module b20s(CK,G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G6762,G6805,G6806,G6807,G6761,G6760,G6808,G6809,G6759,G6758,G6797,G6798,G6799,G6800,G6801,G6802,G6803,G6804,G6763,G6796,G647,G644);
input CK,G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32;
output G6762,G6805,G6806,G6807,G6761,G6760,G6808,G6809,G6759,G6758,G6797,G6798,G6799,G6800,G6801,G6802,G6803,G6804,G6763,G6796,G647,G644;

  wire G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,
       G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,G40,
       G41,G42,G43,G44,G45,G46,G47,G48,G49,G50,G51,G52,G53,G54,G55,G56,G57,G58,G59,G60,
       G61,G62,G63,G64,G65,G66,G67,G68,G69,G70,G71,G72,G73,G74,G75,G76,G77,G78,G79,G80,
       G81,G82,G83,G84,G85,G86,G87,G88,G89,G90,G91,G92,G93,G94,G95,G96,G97,G98,G99,G100,
       G101,G102,G103,G104,G105,G106,G107,G108,G109,G110,G111,G112,G113,G114,G115,G116,G117,G118,G119,G120,
       G121,G122,G123,G124,G125,G126,G127,G128,G129,G130,G131,G132,G133,G134,G135,G136,G137,G138,G139,G140,
       G141,G142,G143,G144,G145,G146,G147,G148,G149,G150,G151,G152,G153,G154,G155,G156,G157,G158,G159,G160,
       G161,G162,G163,G164,G165,G166,G167,G168,G169,G170,G171,G172,G173,G174,G175,G176,G177,G178,G179,G180,
       G181,G182,G183,G184,G185,G186,G187,G188,G189,G190,G191,G192,G193,G194,G195,G196,G197,G198,G199,G200,
       G201,G202,G203,G204,G205,G206,G207,G208,G209,G210,G211,G212,G213,G214,G215,G216,G217,G218,G219,G220,
       G221,G222,G223,G224,G225,G226,G227,G228,G229,G230,G231,G232,G233,G234,G235,G236,G237,G238,G239,G240,
       G241,G242,G243,G244,G245,G246,G247,G248,G249,G250,G251,G252,G253,G254,G255,G256,G257,G258,G259,G260,
       G261,G262,G263,G264,G265,G266,G267,G268,G269,G270,G271,G272,G273,G274,G275,G276,G277,G278,G279,G280,
       G281,G282,G283,G284,G285,G286,G287,G288,G289,G290,G291,G292,G293,G294,G295,G296,G297,G298,G299,G300,
       G301,G302,G303,G304,G305,G306,G307,G308,G309,G310,G311,G312,G313,G314,G315,G316,G317,G318,G319,G320,
       G321,G322,G323,G324,G325,G326,G327,G328,G329,G330,G331,G332,G333,G334,G335,G336,G337,G338,G339,G340,
       G341,G342,G343,G344,G345,G346,G347,G348,G349,G350,G351,G352,G353,G354,G355,G356,G357,G358,G359,G360,
       G361,G362,G363,G364,G365,G366,G367,G368,G369,G370,G371,G372,G373,G374,G375,G376,G377,G378,G379,G380,
       G381,G382,G383,G384,G385,G386,G387,G388,G389,G390,G391,G392,G393,G394,G395,G396,G397,G398,G399,G400,
       G401,G402,G403,G404,G405,G406,G407,G408,G409,G410,G411,G412,G413,G414,G415,G416,G417,G418,G419,G420,
       G421,G422,G423,G424,G425,G426,G427,G428,G429,G430,G431,G432,G433,G434,G435,G436,G437,G438,G439,G440,
       G441,G442,G443,G444,G445,G446,G447,G448,G449,G450,G451,G452,G453,G454,G455,G456,G457,G458,G459,G460,
       G461,G462,G463,G464,G465,G466,G467,G468,G469,G470,G471,G472,G473,G474,G475,G476,G477,G478,G479,G480,
       G481,G482,G483,G484,G485,G486,G487,G488,G489,G490,G491,G492,G493,G494,G495,G496,G497,G498,G499,G500,
       G501,G502,G503,G504,G505,G506,G507,G508,G509,G510,G511,G512,G513,G514,G515,G516,G517,G518,G519,G520,
       G521,G522,G523,G524,G525,G526,G527,G528,G529,G530,G531,G532,G533,G534,G535,G536,G537,G538,G539,G540,
       G541,G542,G543,G544,G545,G546,G547,G548,G549,G550,G551,G552,G553,G554,G555,G556,G557,G558,G559,G560,
       G561,G562,G563,G564,G565,G566,G567,G568,G569,G570,G571,G572,G573,G574,G575,G576,G577,G578,G579,G580,
       G581,G582,G583,G584,G585,G586,G587,G588,G589,G590,G591,G592,G593,G594,G595,G596,G597,G598,G599,G600,
       G601,G602,G603,G604,G605,G606,G607,G608,G609,G610,G611,G612,G613,G614,G615,G616,G617,G618,G619,G620,
       G621,G622,G623,G624,G625,G626,G627,G628,G629,G630,G631,G632,G633,G634,G635,G636,G637,G638,G639,G640,
       G641,G642,G643,G644,G645,G646,G647,G648,G649,G650,G651,G652,G653,G654,G655,G656,G657,G658,G659,G660,
       G661,G662,G663,G664,G665,G666,G667,G668,G669,G670,G671,G672,G673,G674,G675,G676,G677,G678,G679,G680,
       G681,G682,G683,G684,G685,G686,G687,G688,G689,G690,G691,G692,G693,G694,G695,G696,G697,G698,G699,G700,
       G701,G702,G703,G704,G705,G706,G707,G708,G709,G710,G711,G712,G713,G714,G715,G716,G717,G718,G719,G720,
       G721,G722,G723,G724,G725,G726,G727,G728,G729,G730,G731,G732,G733,G734,G735,G736,G737,G738,G739,G740,
       G741,G742,G743,G744,G745,G746,G747,G748,G749,G750,G751,G752,G753,G754,G755,G756,G757,G758,G759,G760,
       G761,G762,G763,G764,G765,G766,G767,G768,G769,G770,G771,G772,G773,G774,G775,G776,G777,G778,G779,G780,
       G781,G782,G783,G784,G785,G786,G787,G788,G789,G790,G791,G792,G793,G794,G795,G796,G797,G798,G799,G800,
       G801,G802,G803,G804,G805,G806,G807,G808,G809,G810,G811,G812,G813,G814,G815,G816,G817,G818,G819,G820,
       G821,G822,G823,G824,G825,G826,G827,G828,G829,G830,G831,G832,G833,G834,G835,G836,G837,G838,G839,G840,
       G841,G842,G843,G844,G845,G846,G847,G848,G849,G850,G851,G852,G853,G854,G855,G856,G857,G858,G859,G860,
       G861,G862,G863,G864,G865,G866,G867,G868,G869,G870,G871,G872,G873,G874,G875,G876,G877,G878,G879,G880,
       G881,G882,G883,G884,G885,G886,G887,G888,G889,G890,G891,G892,G893,G894,G895,G896,G897,G898,G899,G900,
       G901,G902,G903,G904,G905,G906,G907,G908,G909,G910,G911,G912,G913,G914,G915,G916,G917,G918,G919,G920,
       G921,G922,G923,G924,G925,G926,G927,G928,G929,G930,G931,G932,G933,G934,G935,G936,G937,G938,G939,G940,
       G941,G942,G943,G944,G945,G946,G947,G948,G949,G950,G951,G952,G953,G954,G955,G956,G957,G958,G959,G960,
       G961,G962,G963,G964,G965,G966,G967,G968,G969,G970,G971,G972,G973,G974,G975,G976,G977,G978,G979,G980,
       G981,G982,G983,G984,G985,G986,G987,G988,G989,G990,G991,G992,G993,G994,G995,G996,G997,G998,G999,G1000,
       G1001,G1002,G1003,G1004,G1005,G1006,G1007,G1008,G1009,G1010,G1011,G1012,G1013,G1014,G1015,G1016,G1017,G1018,G1019,G1020,
       G1021,G1022,G1023,G1024,G1025,G1026,G1027,G1028,G1029,G1030,G1031,G1032,G1033,G1034,G1035,G1036,G1037,G1038,G1039,G1040,
       G1041,G1042,G1043,G1044,G1045,G1046,G1047,G1048,G1049,G1050,G1051,G1052,G1053,G1054,G1055,G1056,G1057,G1058,G1059,G1060,
       G1061,G1062,G1063,G1064,G1065,G1066,G1067,G1068,G1069,G1070,G1071,G1072,G1073,G1074,G1075,G1076,G1077,G1078,G1079,G1080,
       G1081,G1082,G1083,G1084,G1085,G1086,G1087,G1088,G1089,G1090,G1091,G1092,G1093,G1094,G1095,G1096,G1097,G1098,G1099,G1100,
       G1101,G1102,G1103,G1104,G1105,G1106,G1107,G1108,G1109,G1110,G1111,G1112,G1113,G1114,G1115,G1116,G1117,G1118,G1119,G1120,
       G1121,G1122,G1123,G1124,G1125,G1126,G1127,G1128,G1129,G1130,G1131,G1132,G1133,G1134,G1135,G1136,G1137,G1138,G1139,G1140,
       G1141,G1142,G1143,G1144,G1145,G1146,G1147,G1148,G1149,G1150,G1151,G1152,G1153,G1154,G1155,G1156,G1157,G1158,G1159,G1160,
       G1161,G1162,G1163,G1164,G1165,G1166,G1167,G1168,G1169,G1170,G1171,G1172,G1173,G1174,G1175,G1176,G1177,G1178,G1179,G1180,
       G1181,G1182,G1183,G1184,G1185,G1186,G1187,G1188,G1189,G1190,G1191,G1192,G1193,G1194,G1195,G1196,G1197,G1198,G1199,G1200,
       G1201,G1202,G1203,G1204,G1205,G1206,G1207,G1208,G1209,G1210,G1211,G1212,G1213,G1214,G1215,G1216,G1217,G1218,G1219,G1220,
       G1221,G1222,G1223,G1224,G1225,G1226,G1227,G1228,G1229,G1230,G1231,G1232,G1233,G1234,G1235,G1236,G1237,G1238,G1239,G1240,
       G1241,G1242,G1243,G1244,G1245,G1246,G1247,G1248,G1249,G1250,G1251,G1252,G1253,G1254,G1255,G1256,G1257,G1258,G1259,G1260,
       G1261,G1262,G1263,G1264,G1265,G1266,G1267,G1268,G1269,G1270,G1271,G1272,G1273,G1274,G1275,G1276,G1277,G1278,G1279,G1280,
       G1281,G1282,G1283,G1284,G1285,G1286,G1287,G1288,G1289,G1290,G1291,G1292,G1293,G1294,G1295,G1296,G1297,G1298,G1299,G1300,
       G1301,G1302,G1303,G1304,G1305,G1306,G1307,G1308,G1309,G1310,G1311,G1312,G1313,G1314,G1315,G1316,G1317,G1318,G1319,G1320,
       G1321,G1322,G1323,G1324,G1325,G1326,G1327,G1328,G1329,G1330,G1331,G1332,G1333,G1334,G1335,G1336,G1337,G1338,G1339,G1340,
       G1341,G1342,G1343,G1344,G1345,G1346,G1347,G1348,G1349,G1350,G1351,G1352,G1353,G1354,G1355,G1356,G1357,G1358,G1359,G1360,
       G1361,G1362,G1363,G1364,G1365,G1366,G1367,G1368,G1369,G1370,G1371,G1372,G1373,G1374,G1375,G1376,G1377,G1378,G1379,G1380,
       G1381,G1382,G1383,G1384,G1385,G1386,G1387,G1388,G1389,G1390,G1391,G1392,G1393,G1394,G1395,G1396,G1397,G1398,G1399,G1400,
       G1401,G1402,G1403,G1404,G1405,G1406,G1407,G1408,G1409,G1410,G1411,G1412,G1413,G1414,G1415,G1416,G1417,G1418,G1419,G1420,
       G1421,G1422,G1423,G1424,G1425,G1426,G1427,G1428,G1429,G1430,G1431,G1432,G1433,G1434,G1435,G1436,G1437,G1438,G1439,G1440,
       G1441,G1442,G1443,G1444,G1445,G1446,G1447,G1448,G1449,G1450,G1451,G1452,G1453,G1454,G1455,G1456,G1457,G1458,G1459,G1460,
       G1461,G1462,G1463,G1464,G1465,G1466,G1467,G1468,G1469,G1470,G1471,G1472,G1473,G1474,G1475,G1476,G1477,G1478,G1479,G1480,
       G1481,G1482,G1483,G1484,G1485,G1486,G1487,G1488,G1489,G1490,G1491,G1492,G1493,G1494,G1495,G1496,G1497,G1498,G1499,G1500,
       G1501,G1502,G1503,G1504,G1505,G1506,G1507,G1508,G1509,G1510,G1511,G1512,G1513,G1514,G1515,G1516,G1517,G1518,G1519,G1520,
       G1521,G1522,G1523,G1524,G1525,G1526,G1527,G1528,G1529,G1530,G1531,G1532,G1533,G1534,G1535,G1536,G1537,G1538,G1539,G1540,
       G1541,G1542,G1543,G1544,G1545,G1546,G1547,G1548,G1549,G1550,G1551,G1552,G1553,G1554,G1555,G1556,G1557,G1558,G1559,G1560,
       G1561,G1562,G1563,G1564,G1565,G1566,G1567,G1568,G1569,G1570,G1571,G1572,G1573,G1574,G1575,G1576,G1577,G1578,G1579,G1580,
       G1581,G1582,G1583,G1584,G1585,G1586,G1587,G1588,G1589,G1590,G1591,G1592,G1593,G1594,G1595,G1596,G1597,G1598,G1599,G1600,
       G1601,G1602,G1603,G1604,G1605,G1606,G1607,G1608,G1609,G1610,G1611,G1612,G1613,G1614,G1615,G1616,G1617,G1618,G1619,G1620,
       G1621,G1622,G1623,G1624,G1625,G1626,G1627,G1628,G1629,G1630,G1631,G1632,G1633,G1634,G1635,G1636,G1637,G1638,G1639,G1640,
       G1641,G1642,G1643,G1644,G1645,G1646,G1647,G1648,G1649,G1650,G1651,G1652,G1653,G1654,G1655,G1656,G1657,G1658,G1659,G1660,
       G1661,G1662,G1663,G1664,G1665,G1666,G1667,G1668,G1669,G1670,G1671,G1672,G1673,G1674,G1675,G1676,G1677,G1678,G1679,G1680,
       G1681,G1682,G1683,G1684,G1685,G1686,G1687,G1688,G1689,G1690,G1691,G1692,G1693,G1694,G1695,G1696,G1697,G1698,G1699,G1700,
       G1701,G1702,G1703,G1704,G1705,G1706,G1707,G1708,G1709,G1710,G1711,G1712,G1713,G1714,G1715,G1716,G1717,G1718,G1719,G1720,
       G1721,G1722,G1723,G1724,G1725,G1726,G1727,G1728,G1729,G1730,G1731,G1732,G1733,G1734,G1735,G1736,G1737,G1738,G1739,G1740,
       G1741,G1742,G1743,G1744,G1745,G1746,G1747,G1748,G1749,G1750,G1751,G1752,G1753,G1754,G1755,G1756,G1757,G1758,G1759,G1760,
       G1761,G1762,G1763,G1764,G1765,G1766,G1767,G1768,G1769,G1770,G1771,G1772,G1773,G1774,G1775,G1776,G1777,G1778,G1779,G1780,
       G1781,G1782,G1783,G1784,G1785,G1786,G1787,G1788,G1789,G1790,G1791,G1792,G1793,G1794,G1795,G1796,G1797,G1798,G1799,G1800,
       G1801,G1802,G1803,G1804,G1805,G1806,G1807,G1808,G1809,G1810,G1811,G1812,G1813,G1814,G1815,G1816,G1817,G1818,G1819,G1820,
       G1821,G1822,G1823,G1824,G1825,G1826,G1827,G1828,G1829,G1830,G1831,G1832,G1833,G1834,G1835,G1836,G1837,G1838,G1839,G1840,
       G1841,G1842,G1843,G1844,G1845,G1846,G1847,G1848,G1849,G1850,G1851,G1852,G1853,G1854,G1855,G1856,G1857,G1858,G1859,G1860,
       G1861,G1862,G1863,G1864,G1865,G1866,G1867,G1868,G1869,G1870,G1871,G1872,G1873,G1874,G1875,G1876,G1877,G1878,G1879,G1880,
       G1881,G1882,G1883,G1884,G1885,G1886,G1887,G1888,G1889,G1890,G1891,G1892,G1893,G1894,G1895,G1896,G1897,G1898,G1899,G1900,
       G1901,G1902,G1903,G1904,G1905,G1906,G1907,G1908,G1909,G1910,G1911,G1912,G1913,G1914,G1915,G1916,G1917,G1918,G1919,G1920,
       G1921,G1922,G1923,G1924,G1925,G1926,G1927,G1928,G1929,G1930,G1931,G1932,G1933,G1934,G1935,G1936,G1937,G1938,G1939,G1940,
       G1941,G1942,G1943,G1944,G1945,G1946,G1947,G1948,G1949,G1950,G1951,G1952,G1953,G1954,G1955,G1956,G1957,G1958,G1959,G1960,
       G1961,G1962,G1963,G1964,G1965,G1966,G1967,G1968,G1969,G1970,G1971,G1972,G1973,G1974,G1975,G1976,G1977,G1978,G1979,G1980,
       G1981,G1982,G1983,G1984,G1985,G1986,G1987,G1988,G1989,G1990,G1991,G1992,G1993,G1994,G1995,G1996,G1997,G1998,G1999,G2000,
       G2001,G2002,G2003,G2004,G2005,G2006,G2007,G2008,G2009,G2010,G2011,G2012,G2013,G2014,G2015,G2016,G2017,G2018,G2019,G2020,
       G2021,G2022,G2023,G2024,G2025,G2026,G2027,G2028,G2029,G2030,G2031,G2032,G2033,G2034,G2035,G2036,G2037,G2038,G2039,G2040,
       G2041,G2042,G2043,G2044,G2045,G2046,G2047,G2048,G2049,G2050,G2051,G2052,G2053,G2054,G2055,G2056,G2057,G2058,G2059,G2060,
       G2061,G2062,G2063,G2064,G2065,G2066,G2067,G2068,G2069,G2070,G2071,G2072,G2073,G2074,G2075,G2076,G2077,G2078,G2079,G2080,
       G2081,G2082,G2083,G2084,G2085,G2086,G2087,G2088,G2089,G2090,G2091,G2092,G2093,G2094,G2095,G2096,G2097,G2098,G2099,G2100,
       G2101,G2102,G2103,G2104,G2105,G2106,G2107,G2108,G2109,G2110,G2111,G2112,G2113,G2114,G2115,G2116,G2117,G2118,G2119,G2120,
       G2121,G2122,G2123,G2124,G2125,G2126,G2127,G2128,G2129,G2130,G2131,G2132,G2133,G2134,G2135,G2136,G2137,G2138,G2139,G2140,
       G2141,G2142,G2143,G2144,G2145,G2146,G2147,G2148,G2149,G2150,G2151,G2152,G2153,G2154,G2155,G2156,G2157,G2158,G2159,G2160,
       G2161,G2162,G2163,G2164,G2165,G2166,G2167,G2168,G2169,G2170,G2171,G2172,G2173,G2174,G2175,G2176,G2177,G2178,G2179,G2180,
       G2181,G2182,G2183,G2184,G2185,G2186,G2187,G2188,G2189,G2190,G2191,G2192,G2193,G2194,G2195,G2196,G2197,G2198,G2199,G2200,
       G2201,G2202,G2203,G2204,G2205,G2206,G2207,G2208,G2209,G2210,G2211,G2212,G2213,G2214,G2215,G2216,G2217,G2218,G2219,G2220,
       G2221,G2222,G2223,G2224,G2225,G2226,G2227,G2228,G2229,G2230,G2231,G2232,G2233,G2234,G2235,G2236,G2237,G2238,G2239,G2240,
       G2241,G2242,G2243,G2244,G2245,G2246,G2247,G2248,G2249,G2250,G2251,G2252,G2253,G2254,G2255,G2256,G2257,G2258,G2259,G2260,
       G2261,G2262,G2263,G2264,G2265,G2266,G2267,G2268,G2269,G2270,G2271,G2272,G2273,G2274,G2275,G2276,G2277,G2278,G2279,G2280,
       G2281,G2282,G2283,G2284,G2285,G2286,G2287,G2288,G2289,G2290,G2291,G2292,G2293,G2294,G2295,G2296,G2297,G2298,G2299,G2300,
       G2301,G2302,G2303,G2304,G2305,G2306,G2307,G2308,G2309,G2310,G2311,G2312,G2313,G2314,G2315,G2316,G2317,G2318,G2319,G2320,
       G2321,G2322,G2323,G2324,G2325,G2326,G2327,G2328,G2329,G2330,G2331,G2332,G2333,G2334,G2335,G2336,G2337,G2338,G2339,G2340,
       G2341,G2342,G2343,G2344,G2345,G2346,G2347,G2348,G2349,G2350,G2351,G2352,G2353,G2354,G2355,G2356,G2357,G2358,G2359,G2360,
       G2361,G2362,G2363,G2364,G2365,G2366,G2367,G2368,G2369,G2370,G2371,G2372,G2373,G2374,G2375,G2376,G2377,G2378,G2379,G2380,
       G2381,G2382,G2383,G2384,G2385,G2386,G2387,G2388,G2389,G2390,G2391,G2392,G2393,G2394,G2395,G2396,G2397,G2398,G2399,G2400,
       G2401,G2402,G2403,G2404,G2405,G2406,G2407,G2408,G2409,G2410,G2411,G2412,G2413,G2414,G2415,G2416,G2417,G2418,G2419,G2420,
       G2421,G2422,G2423,G2424,G2425,G2426,G2427,G2428,G2429,G2430,G2431,G2432,G2433,G2434,G2435,G2436,G2437,G2438,G2439,G2440,
       G2441,G2442,G2443,G2444,G2445,G2446,G2447,G2448,G2449,G2450,G2451,G2452,G2453,G2454,G2455,G2456,G2457,G2458,G2459,G2460,
       G2461,G2462,G2463,G2464,G2465,G2466,G2467,G2468,G2469,G2470,G2471,G2472,G2473,G2474,G2475,G2476,G2477,G2478,G2479,G2480,
       G2481,G2482,G2483,G2484,G2485,G2486,G2487,G2488,G2489,G2490,G2491,G2492,G2493,G2494,G2495,G2496,G2497,G2498,G2499,G2500,
       G2501,G2502,G2503,G2504,G2505,G2506,G2507,G2508,G2509,G2510,G2511,G2512,G2513,G2514,G2515,G2516,G2517,G2518,G2519,G2520,
       G2521,G2522,G2523,G2524,G2525,G2526,G2527,G2528,G2529,G2530,G2531,G2532,G2533,G2534,G2535,G2536,G2537,G2538,G2539,G2540,
       G2541,G2542,G2543,G2544,G2545,G2546,G2547,G2548,G2549,G2550,G2551,G2552,G2553,G2554,G2555,G2556,G2557,G2558,G2559,G2560,
       G2561,G2562,G2563,G2564,G2565,G2566,G2567,G2568,G2569,G2570,G2571,G2572,G2573,G2574,G2575,G2576,G2577,G2578,G2579,G2580,
       G2581,G2582,G2583,G2584,G2585,G2586,G2587,G2588,G2589,G2590,G2591,G2592,G2593,G2594,G2595,G2596,G2597,G2598,G2599,G2600,
       G2601,G2602,G2603,G2604,G2605,G2606,G2607,G2608,G2609,G2610,G2611,G2612,G2613,G2614,G2615,G2616,G2617,G2618,G2619,G2620,
       G2621,G2622,G2623,G2624,G2625,G2626,G2627,G2628,G2629,G2630,G2631,G2632,G2633,G2634,G2635,G2636,G2637,G2638,G2639,G2640,
       G2641,G2642,G2643,G2644,G2645,G2646,G2647,G2648,G2649,G2650,G2651,G2652,G2653,G2654,G2655,G2656,G2657,G2658,G2659,G2660,
       G2661,G2662,G2663,G2664,G2665,G2666,G2667,G2668,G2669,G2670,G2671,G2672,G2673,G2674,G2675,G2676,G2677,G2678,G2679,G2680,
       G2681,G2682,G2683,G2684,G2685,G2686,G2687,G2688,G2689,G2690,G2691,G2692,G2693,G2694,G2695,G2696,G2697,G2698,G2699,G2700,
       G2701,G2702,G2703,G2704,G2705,G2706,G2707,G2708,G2709,G2710,G2711,G2712,G2713,G2714,G2715,G2716,G2717,G2718,G2719,G2720,
       G2721,G2722,G2723,G2724,G2725,G2726,G2727,G2728,G2729,G2730,G2731,G2732,G2733,G2734,G2735,G2736,G2737,G2738,G2739,G2740,
       G2741,G2742,G2743,G2744,G2745,G2746,G2747,G2748,G2749,G2750,G2751,G2752,G2753,G2754,G2755,G2756,G2757,G2758,G2759,G2760,
       G2761,G2762,G2763,G2764,G2765,G2766,G2767,G2768,G2769,G2770,G2771,G2772,G2773,G2774,G2775,G2776,G2777,G2778,G2779,G2780,
       G2781,G2782,G2783,G2784,G2785,G2786,G2787,G2788,G2789,G2790,G2791,G2792,G2793,G2794,G2795,G2796,G2797,G2798,G2799,G2800,
       G2801,G2802,G2803,G2804,G2805,G2806,G2807,G2808,G2809,G2810,G2811,G2812,G2813,G2814,G2815,G2816,G2817,G2818,G2819,G2820,
       G2821,G2822,G2823,G2824,G2825,G2826,G2827,G2828,G2829,G2830,G2831,G2832,G2833,G2834,G2835,G2836,G2837,G2838,G2839,G2840,
       G2841,G2842,G2843,G2844,G2845,G2846,G2847,G2848,G2849,G2850,G2851,G2852,G2853,G2854,G2855,G2856,G2857,G2858,G2859,G2860,
       G2861,G2862,G2863,G2864,G2865,G2866,G2867,G2868,G2869,G2870,G2871,G2872,G2873,G2874,G2875,G2876,G2877,G2878,G2879,G2880,
       G2881,G2882,G2883,G2884,G2885,G2886,G2887,G2888,G2889,G2890,G2891,G2892,G2893,G2894,G2895,G2896,G2897,G2898,G2899,G2900,
       G2901,G2902,G2903,G2904,G2905,G2906,G2907,G2908,G2909,G2910,G2911,G2912,G2913,G2914,G2915,G2916,G2917,G2918,G2919,G2920,
       G2921,G2922,G2923,G2924,G2925,G2926,G2927,G2928,G2929,G2930,G2931,G2932,G2933,G2934,G2935,G2936,G2937,G2938,G2939,G2940,
       G2941,G2942,G2943,G2944,G2945,G2946,G2947,G2948,G2949,G2950,G2951,G2952,G2953,G2954,G2955,G2956,G2957,G2958,G2959,G2960,
       G2961,G2962,G2963,G2964,G2965,G2966,G2967,G2968,G2969,G2970,G2971,G2972,G2973,G2974,G2975,G2976,G2977,G2978,G2979,G2980,
       G2981,G2982,G2983,G2984,G2985,G2986,G2987,G2988,G2989,G2990,G2991,G2992,G2993,G2994,G2995,G2996,G2997,G2998,G2999,G3000,
       G3001,G3002,G3003,G3004,G3005,G3006,G3007,G3008,G3009,G3010,G3011,G3012,G3013,G3014,G3015,G3016,G3017,G3018,G3019,G3020,
       G3021,G3022,G3023,G3024,G3025,G3026,G3027,G3028,G3029,G3030,G3031,G3032,G3033,G3034,G3035,G3036,G3037,G3038,G3039,G3040,
       G3041,G3042,G3043,G3044,G3045,G3046,G3047,G3048,G3049,G3050,G3051,G3052,G3053,G3054,G3055,G3056,G3057,G3058,G3059,G3060,
       G3061,G3062,G3063,G3064,G3065,G3066,G3067,G3068,G3069,G3070,G3071,G3072,G3073,G3074,G3075,G3076,G3077,G3078,G3079,G3080,
       G3081,G3082,G3083,G3084,G3085,G3086,G3087,G3088,G3089,G3090,G3091,G3092,G3093,G3094,G3095,G3096,G3097,G3098,G3099,G3100,
       G3101,G3102,G3103,G3104,G3105,G3106,G3107,G3108,G3109,G3110,G3111,G3112,G3113,G3114,G3115,G3116,G3117,G3118,G3119,G3120,
       G3121,G3122,G3123,G3124,G3125,G3126,G3127,G3128,G3129,G3130,G3131,G3132,G3133,G3134,G3135,G3136,G3137,G3138,G3139,G3140,
       G3141,G3142,G3143,G3144,G3145,G3146,G3147,G3148,G3149,G3150,G3151,G3152,G3153,G3154,G3155,G3156,G3157,G3158,G3159,G3160,
       G3161,G3162,G3163,G3164,G3165,G3166,G3167,G3168,G3169,G3170,G3171,G3172,G3173,G3174,G3175,G3176,G3177,G3178,G3179,G3180,
       G3181,G3182,G3183,G3184,G3185,G3186,G3187,G3188,G3189,G3190,G3191,G3192,G3193,G3194,G3195,G3196,G3197,G3198,G3199,G3200,
       G3201,G3202,G3203,G3204,G3205,G3206,G3207,G3208,G3209,G3210,G3211,G3212,G3213,G3214,G3215,G3216,G3217,G3218,G3219,G3220,
       G3221,G3222,G3223,G3224,G3225,G3226,G3227,G3228,G3229,G3230,G3231,G3232,G3233,G3234,G3235,G3236,G3237,G3238,G3239,G3240,
       G3241,G3242,G3243,G3244,G3245,G3246,G3247,G3248,G3249,G3250,G3251,G3252,G3253,G3254,G3255,G3256,G3257,G3258,G3259,G3260,
       G3261,G3262,G3263,G3264,G3265,G3266,G3267,G3268,G3269,G3270,G3271,G3272,G3273,G3274,G3275,G3276,G3277,G3278,G3279,G3280,
       G3281,G3282,G3283,G3284,G3285,G3286,G3287,G3288,G3289,G3290,G3291,G3292,G3293,G3294,G3295,G3296,G3297,G3298,G3299,G3300,
       G3301,G3302,G3303,G3304,G3305,G3306,G3307,G3308,G3309,G3310,G3311,G3312,G3313,G3314,G3315,G3316,G3317,G3318,G3319,G3320,
       G3321,G3322,G3323,G3324,G3325,G3326,G3327,G3328,G3329,G3330,G3331,G3332,G3333,G3334,G3335,G3336,G3337,G3338,G3339,G3340,
       G3341,G3342,G3343,G3344,G3345,G3346,G3347,G3348,G3349,G3350,G3351,G3352,G3353,G3354,G3355,G3356,G3357,G3358,G3359,G3360,
       G3361,G3362,G3363,G3364,G3365,G3366,G3367,G3368,G3369,G3370,G3371,G3372,G3373,G3374,G3375,G3376,G3377,G3378,G3379,G3380,
       G3381,G3382,G3383,G3384,G3385,G3386,G3387,G3388,G3389,G3390,G3391,G3392,G3393,G3394,G3395,G3396,G3397,G3398,G3399,G3400,
       G3401,G3402,G3403,G3404,G3405,G3406,G3407,G3408,G3409,G3410,G3411,G3412,G3413,G3414,G3415,G3416,G3417,G3418,G3419,G3420,
       G3421,G3422,G3423,G3424,G3425,G3426,G3427,G3428,G3429,G3430,G3431,G3432,G3433,G3434,G3435,G3436,G3437,G3438,G3439,G3440,
       G3441,G3442,G3443,G3444,G3445,G3446,G3447,G3448,G3449,G3450,G3451,G3452,G3453,G3454,G3455,G3456,G3457,G3458,G3459,G3460,
       G3461,G3462,G3463,G3464,G3465,G3466,G3467,G3468,G3469,G3470,G3471,G3472,G3473,G3474,G3475,G3476,G3477,G3478,G3479,G3480,
       G3481,G3482,G3483,G3484,G3485,G3486,G3487,G3488,G3489,G3490,G3491,G3492,G3493,G3494,G3495,G3496,G3497,G3498,G3499,G3500,
       G3501,G3502,G3503,G3504,G3505,G3506,G3507,G3508,G3509,G3510,G3511,G3512,G3513,G3514,G3515,G3516,G3517,G3518,G3519,G3520,
       G3521,G3522,G3523,G3524,G3525,G3526,G3527,G3528,G3529,G3530,G3531,G3532,G3533,G3534,G3535,G3536,G3537,G3538,G3539,G3540,
       G3541,G3542,G3543,G3544,G3545,G3546,G3547,G3548,G3549,G3550,G3551,G3552,G3553,G3554,G3555,G3556,G3557,G3558,G3559,G3560,
       G3561,G3562,G3563,G3564,G3565,G3566,G3567,G3568,G3569,G3570,G3571,G3572,G3573,G3574,G3575,G3576,G3577,G3578,G3579,G3580,
       G3581,G3582,G3583,G3584,G3585,G3586,G3587,G3588,G3589,G3590,G3591,G3592,G3593,G3594,G3595,G3596,G3597,G3598,G3599,G3600,
       G3601,G3602,G3603,G3604,G3605,G3606,G3607,G3608,G3609,G3610,G3611,G3612,G3613,G3614,G3615,G3616,G3617,G3618,G3619,G3620,
       G3621,G3622,G3623,G3624,G3625,G3626,G3627,G3628,G3629,G3630,G3631,G3632,G3633,G3634,G3635,G3636,G3637,G3638,G3639,G3640,
       G3641,G3642,G3643,G3644,G3645,G3646,G3647,G3648,G3649,G3650,G3651,G3652,G3653,G3654,G3655,G3656,G3657,G3658,G3659,G3660,
       G3661,G3662,G3663,G3664,G3665,G3666,G3667,G3668,G3669,G3670,G3671,G3672,G3673,G3674,G3675,G3676,G3677,G3678,G3679,G3680,
       G3681,G3682,G3683,G3684,G3685,G3686,G3687,G3688,G3689,G3690,G3691,G3692,G3693,G3694,G3695,G3696,G3697,G3698,G3699,G3700,
       G3701,G3702,G3703,G3704,G3705,G3706,G3707,G3708,G3709,G3710,G3711,G3712,G3713,G3714,G3715,G3716,G3717,G3718,G3719,G3720,
       G3721,G3722,G3723,G3724,G3725,G3726,G3727,G3728,G3729,G3730,G3731,G3732,G3733,G3734,G3735,G3736,G3737,G3738,G3739,G3740,
       G3741,G3742,G3743,G3744,G3745,G3746,G3747,G3748,G3749,G3750,G3751,G3752,G3753,G3754,G3755,G3756,G3757,G3758,G3759,G3760,
       G3761,G3762,G3763,G3764,G3765,G3766,G3767,G3768,G3769,G3770,G3771,G3772,G3773,G3774,G3775,G3776,G3777,G3778,G3779,G3780,
       G3781,G3782,G3783,G3784,G3785,G3786,G3787,G3788,G3789,G3790,G3791,G3792,G3793,G3794,G3795,G3796,G3797,G3798,G3799,G3800,
       G3801,G3802,G3803,G3804,G3805,G3806,G3807,G3808,G3809,G3810,G3811,G3812,G3813,G3814,G3815,G3816,G3817,G3818,G3819,G3820,
       G3821,G3822,G3823,G3824,G3825,G3826,G3827,G3828,G3829,G3830,G3831,G3832,G3833,G3834,G3835,G3836,G3837,G3838,G3839,G3840,
       G3841,G3842,G3843,G3844,G3845,G3846,G3847,G3848,G3849,G3850,G3851,G3852,G3853,G3854,G3855,G3856,G3857,G3858,G3859,G3860,
       G3861,G3862,G3863,G3864,G3865,G3866,G3867,G3868,G3869,G3870,G3871,G3872,G3873,G3874,G3875,G3876,G3877,G3878,G3879,G3880,
       G3881,G3882,G3883,G3884,G3885,G3886,G3887,G3888,G3889,G3890,G3891,G3892,G3893,G3894,G3895,G3896,G3897,G3898,G3899,G3900,
       G3901,G3902,G3903,G3904,G3905,G3906,G3907,G3908,G3909,G3910,G3911,G3912,G3913,G3914,G3915,G3916,G3917,G3918,G3919,G3920,
       G3921,G3922,G3923,G3924,G3925,G3926,G3927,G3928,G3929,G3930,G3931,G3932,G3933,G3934,G3935,G3936,G3937,G3938,G3939,G3940,
       G3941,G3942,G3943,G3944,G3945,G3946,G3947,G3948,G3949,G3950,G3951,G3952,G3953,G3954,G3955,G3956,G3957,G3958,G3959,G3960,
       G3961,G3962,G3963,G3964,G3965,G3966,G3967,G3968,G3969,G3970,G3971,G3972,G3973,G3974,G3975,G3976,G3977,G3978,G3979,G3980,
       G3981,G3982,G3983,G3984,G3985,G3986,G3987,G3988,G3989,G3990,G3991,G3992,G3993,G3994,G3995,G3996,G3997,G3998,G3999,G4000,
       G4001,G4002,G4003,G4004,G4005,G4006,G4007,G4008,G4009,G4010,G4011,G4012,G4013,G4014,G4015,G4016,G4017,G4018,G4019,G4020,
       G4021,G4022,G4023,G4024,G4025,G4026,G4027,G4028,G4029,G4030,G4031,G4032,G4033,G4034,G4035,G4036,G4037,G4038,G4039,G4040,
       G4041,G4042,G4043,G4044,G4045,G4046,G4047,G4048,G4049,G4050,G4051,G4052,G4053,G4054,G4055,G4056,G4057,G4058,G4059,G4060,
       G4061,G4062,G4063,G4064,G4065,G4066,G4067,G4068,G4069,G4070,G4071,G4072,G4073,G4074,G4075,G4076,G4077,G4078,G4079,G4080,
       G4081,G4082,G4083,G4084,G4085,G4086,G4087,G4088,G4089,G4090,G4091,G4092,G4093,G4094,G4095,G4096,G4097,G4098,G4099,G4100,
       G4101,G4102,G4103,G4104,G4105,G4106,G4107,G4108,G4109,G4110,G4111,G4112,G4113,G4114,G4115,G4116,G4117,G4118,G4119,G4120,
       G4121,G4122,G4123,G4124,G4125,G4126,G4127,G4128,G4129,G4130,G4131,G4132,G4133,G4134,G4135,G4136,G4137,G4138,G4139,G4140,
       G4141,G4142,G4143,G4144,G4145,G4146,G4147,G4148,G4149,G4150,G4151,G4152,G4153,G4154,G4155,G4156,G4157,G4158,G4159,G4160,
       G4161,G4162,G4163,G4164,G4165,G4166,G4167,G4168,G4169,G4170,G4171,G4172,G4173,G4174,G4175,G4176,G4177,G4178,G4179,G4180,
       G4181,G4182,G4183,G4184,G4185,G4186,G4187,G4188,G4189,G4190,G4191,G4192,G4193,G4194,G4195,G4196,G4197,G4198,G4199,G4200,
       G4201,G4202,G4203,G4204,G4205,G4206,G4207,G4208,G4209,G4210,G4211,G4212,G4213,G4214,G4215,G4216,G4217,G4218,G4219,G4220,
       G4221,G4222,G4223,G4224,G4225,G4226,G4227,G4228,G4229,G4230,G4231,G4232,G4233,G4234,G4235,G4236,G4237,G4238,G4239,G4240,
       G4241,G4242,G4243,G4244,G4245,G4246,G4247,G4248,G4249,G4250,G4251,G4252,G4253,G4254,G4255,G4256,G4257,G4258,G4259,G4260,
       G4261,G4262,G4263,G4264,G4265,G4266,G4267,G4268,G4269,G4270,G4271,G4272,G4273,G4274,G4275,G4276,G4277,G4278,G4279,G4280,
       G4281,G4282,G4283,G4284,G4285,G4286,G4287,G4288,G4289,G4290,G4291,G4292,G4293,G4294,G4295,G4296,G4297,G4298,G4299,G4300,
       G4301,G4302,G4303,G4304,G4305,G4306,G4307,G4308,G4309,G4310,G4311,G4312,G4313,G4314,G4315,G4316,G4317,G4318,G4319,G4320,
       G4321,G4322,G4323,G4324,G4325,G4326,G4327,G4328,G4329,G4330,G4331,G4332,G4333,G4334,G4335,G4336,G4337,G4338,G4339,G4340,
       G4341,G4342,G4343,G4344,G4345,G4346,G4347,G4348,G4349,G4350,G4351,G4352,G4353,G4354,G4355,G4356,G4357,G4358,G4359,G4360,
       G4361,G4362,G4363,G4364,G4365,G4366,G4367,G4368,G4369,G4370,G4371,G4372,G4373,G4374,G4375,G4376,G4377,G4378,G4379,G4380,
       G4381,G4382,G4383,G4384,G4385,G4386,G4387,G4388,G4389,G4390,G4391,G4392,G4393,G4394,G4395,G4396,G4397,G4398,G4399,G4400,
       G4401,G4402,G4403,G4404,G4405,G4406,G4407,G4408,G4409,G4410,G4411,G4412,G4413,G4414,G4415,G4416,G4417,G4418,G4419,G4420,
       G4421,G4422,G4423,G4424,G4425,G4426,G4427,G4428,G4429,G4430,G4431,G4432,G4433,G4434,G4435,G4436,G4437,G4438,G4439,G4440,
       G4441,G4442,G4443,G4444,G4445,G4446,G4447,G4448,G4449,G4450,G4451,G4452,G4453,G4454,G4455,G4456,G4457,G4458,G4459,G4460,
       G4461,G4462,G4463,G4464,G4465,G4466,G4467,G4468,G4469,G4470,G4471,G4472,G4473,G4474,G4475,G4476,G4477,G4478,G4479,G4480,
       G4481,G4482,G4483,G4484,G4485,G4486,G4487,G4488,G4489,G4490,G4491,G4492,G4493,G4494,G4495,G4496,G4497,G4498,G4499,G4500,
       G4501,G4502,G4503,G4504,G4505,G4506,G4507,G4508,G4509,G4510,G4511,G4512,G4513,G4514,G4515,G4516,G4517,G4518,G4519,G4520,
       G4521,G4522,G4523,G4524,G4525,G4526,G4527,G4528,G4529,G4530,G4531,G4532,G4533,G4534,G4535,G4536,G4537,G4538,G4539,G4540,
       G4541,G4542,G4543,G4544,G4545,G4546,G4547,G4548,G4549,G4550,G4551,G4552,G4553,G4554,G4555,G4556,G4557,G4558,G4559,G4560,
       G4561,G4562,G4563,G4564,G4565,G4566,G4567,G4568,G4569,G4570,G4571,G4572,G4573,G4574,G4575,G4576,G4577,G4578,G4579,G4580,
       G4581,G4582,G4583,G4584,G4585,G4586,G4587,G4588,G4589,G4590,G4591,G4592,G4593,G4594,G4595,G4596,G4597,G4598,G4599,G4600,
       G4601,G4602,G4603,G4604,G4605,G4606,G4607,G4608,G4609,G4610,G4611,G4612,G4613,G4614,G4615,G4616,G4617,G4618,G4619,G4620,
       G4621,G4622,G4623,G4624,G4625,G4626,G4627,G4628,G4629,G4630,G4631,G4632,G4633,G4634,G4635,G4636,G4637,G4638,G4639,G4640,
       G4641,G4642,G4643,G4644,G4645,G4646,G4647,G4648,G4649,G4650,G4651,G4652,G4653,G4654,G4655,G4656,G4657,G4658,G4659,G4660,
       G4661,G4662,G4663,G4664,G4665,G4666,G4667,G4668,G4669,G4670,G4671,G4672,G4673,G4674,G4675,G4676,G4677,G4678,G4679,G4680,
       G4681,G4682,G4683,G4684,G4685,G4686,G4687,G4688,G4689,G4690,G4691,G4692,G4693,G4694,G4695,G4696,G4697,G4698,G4699,G4700,
       G4701,G4702,G4703,G4704,G4705,G4706,G4707,G4708,G4709,G4710,G4711,G4712,G4713,G4714,G4715,G4716,G4717,G4718,G4719,G4720,
       G4721,G4722,G4723,G4724,G4725,G4726,G4727,G4728,G4729,G4730,G4731,G4732,G4733,G4734,G4735,G4736,G4737,G4738,G4739,G4740,
       G4741,G4742,G4743,G4744,G4745,G4746,G4747,G4748,G4749,G4750,G4751,G4752,G4753,G4754,G4755,G4756,G4757,G4758,G4759,G4760,
       G4761,G4762,G4763,G4764,G4765,G4766,G4767,G4768,G4769,G4770,G4771,G4772,G4773,G4774,G4775,G4776,G4777,G4778,G4779,G4780,
       G4781,G4782,G4783,G4784,G4785,G4786,G4787,G4788,G4789,G4790,G4791,G4792,G4793,G4794,G4795,G4796,G4797,G4798,G4799,G4800,
       G4801,G4802,G4803,G4804,G4805,G4806,G4807,G4808,G4809,G4810,G4811,G4812,G4813,G4814,G4815,G4816,G4817,G4818,G4819,G4820,
       G4821,G4822,G4823,G4824,G4825,G4826,G4827,G4828,G4829,G4830,G4831,G4832,G4833,G4834,G4835,G4836,G4837,G4838,G4839,G4840,
       G4841,G4842,G4843,G4844,G4845,G4846,G4847,G4848,G4849,G4850,G4851,G4852,G4853,G4854,G4855,G4856,G4857,G4858,G4859,G4860,
       G4861,G4862,G4863,G4864,G4865,G4866,G4867,G4868,G4869,G4870,G4871,G4872,G4873,G4874,G4875,G4876,G4877,G4878,G4879,G4880,
       G4881,G4882,G4883,G4884,G4885,G4886,G4887,G4888,G4889,G4890,G4891,G4892,G4893,G4894,G4895,G4896,G4897,G4898,G4899,G4900,
       G4901,G4902,G4903,G4904,G4905,G4906,G4907,G4908,G4909,G4910,G4911,G4912,G4913,G4914,G4915,G4916,G4917,G4918,G4919,G4920,
       G4921,G4922,G4923,G4924,G4925,G4926,G4927,G4928,G4929,G4930,G4931,G4932,G4933,G4934,G4935,G4936,G4937,G4938,G4939,G4940,
       G4941,G4942,G4943,G4944,G4945,G4946,G4947,G4948,G4949,G4950,G4951,G4952,G4953,G4954,G4955,G4956,G4957,G4958,G4959,G4960,
       G4961,G4962,G4963,G4964,G4965,G4966,G4967,G4968,G4969,G4970,G4971,G4972,G4973,G4974,G4975,G4976,G4977,G4978,G4979,G4980,
       G4981,G4982,G4983,G4984,G4985,G4986,G4987,G4988,G4989,G4990,G4991,G4992,G4993,G4994,G4995,G4996,G4997,G4998,G4999,G5000,
       G5001,G5002,G5003,G5004,G5005,G5006,G5007,G5008,G5009,G5010,G5011,G5012,G5013,G5014,G5015,G5016,G5017,G5018,G5019,G5020,
       G5021,G5022,G5023,G5024,G5025,G5026,G5027,G5028,G5029,G5030,G5031,G5032,G5033,G5034,G5035,G5036,G5037,G5038,G5039,G5040,
       G5041,G5042,G5043,G5044,G5045,G5046,G5047,G5048,G5049,G5050,G5051,G5052,G5053,G5054,G5055,G5056,G5057,G5058,G5059,G5060,
       G5061,G5062,G5063,G5064,G5065,G5066,G5067,G5068,G5069,G5070,G5071,G5072,G5073,G5074,G5075,G5076,G5077,G5078,G5079,G5080,
       G5081,G5082,G5083,G5084,G5085,G5086,G5087,G5088,G5089,G5090,G5091,G5092,G5093,G5094,G5095,G5096,G5097,G5098,G5099,G5100,
       G5101,G5102,G5103,G5104,G5105,G5106,G5107,G5108,G5109,G5110,G5111,G5112,G5113,G5114,G5115,G5116,G5117,G5118,G5119,G5120,
       G5121,G5122,G5123,G5124,G5125,G5126,G5127,G5128,G5129,G5130,G5131,G5132,G5133,G5134,G5135,G5136,G5137,G5138,G5139,G5140,
       G5141,G5142,G5143,G5144,G5145,G5146,G5147,G5148,G5149,G5150,G5151,G5152,G5153,G5154,G5155,G5156,G5157,G5158,G5159,G5160,
       G5161,G5162,G5163,G5164,G5165,G5166,G5167,G5168,G5169,G5170,G5171,G5172,G5173,G5174,G5175,G5176,G5177,G5178,G5179,G5180,
       G5181,G5182,G5183,G5184,G5185,G5186,G5187,G5188,G5189,G5190,G5191,G5192,G5193,G5194,G5195,G5196,G5197,G5198,G5199,G5200,
       G5201,G5202,G5203,G5204,G5205,G5206,G5207,G5208,G5209,G5210,G5211,G5212,G5213,G5214,G5215,G5216,G5217,G5218,G5219,G5220,
       G5221,G5222,G5223,G5224,G5225,G5226,G5227,G5228,G5229,G5230,G5231,G5232,G5233,G5234,G5235,G5236,G5237,G5238,G5239,G5240,
       G5241,G5242,G5243,G5244,G5245,G5246,G5247,G5248,G5249,G5250,G5251,G5252,G5253,G5254,G5255,G5256,G5257,G5258,G5259,G5260,
       G5261,G5262,G5263,G5264,G5265,G5266,G5267,G5268,G5269,G5270,G5271,G5272,G5273,G5274,G5275,G5276,G5277,G5278,G5279,G5280,
       G5281,G5282,G5283,G5284,G5285,G5286,G5287,G5288,G5289,G5290,G5291,G5292,G5293,G5294,G5295,G5296,G5297,G5298,G5299,G5300,
       G5301,G5302,G5303,G5304,G5305,G5306,G5307,G5308,G5309,G5310,G5311,G5312,G5313,G5314,G5315,G5316,G5317,G5318,G5319,G5320,
       G5321,G5322,G5323,G5324,G5325,G5326,G5327,G5328,G5329,G5330,G5331,G5332,G5333,G5334,G5335,G5336,G5337,G5338,G5339,G5340,
       G5341,G5342,G5343,G5344,G5345,G5346,G5347,G5348,G5349,G5350,G5351,G5352,G5353,G5354,G5355,G5356,G5357,G5358,G5359,G5360,
       G5361,G5362,G5363,G5364,G5365,G5366,G5367,G5368,G5369,G5370,G5371,G5372,G5373,G5374,G5375,G5376,G5377,G5378,G5379,G5380,
       G5381,G5382,G5383,G5384,G5385,G5386,G5387,G5388,G5389,G5390,G5391,G5392,G5393,G5394,G5395,G5396,G5397,G5398,G5399,G5400,
       G5401,G5402,G5403,G5404,G5405,G5406,G5407,G5408,G5409,G5410,G5411,G5412,G5413,G5414,G5415,G5416,G5417,G5418,G5419,G5420,
       G5421,G5422,G5423,G5424,G5425,G5426,G5427,G5428,G5429,G5430,G5431,G5432,G5433,G5434,G5435,G5436,G5437,G5438,G5439,G5440,
       G5441,G5442,G5443,G5444,G5445,G5446,G5447,G5448,G5449,G5450,G5451,G5452,G5453,G5454,G5455,G5456,G5457,G5458,G5459,G5460,
       G5461,G5462,G5463,G5464,G5465,G5466,G5467,G5468,G5469,G5470,G5471,G5472,G5473,G5474,G5475,G5476,G5477,G5478,G5479,G5480,
       G5481,G5482,G5483,G5484,G5485,G5486,G5487,G5488,G5489,G5490,G5491,G5492,G5493,G5494,G5495,G5496,G5497,G5498,G5499,G5500,
       G5501,G5502,G5503,G5504,G5505,G5506,G5507,G5508,G5509,G5510,G5511,G5512,G5513,G5514,G5515,G5516,G5517,G5518,G5519,G5520,
       G5521,G5522,G5523,G5524,G5525,G5526,G5527,G5528,G5529,G5530,G5531,G5532,G5533,G5534,G5535,G5536,G5537,G5538,G5539,G5540,
       G5541,G5542,G5543,G5544,G5545,G5546,G5547,G5548,G5549,G5550,G5551,G5552,G5553,G5554,G5555,G5556,G5557,G5558,G5559,G5560,
       G5561,G5562,G5563,G5564,G5565,G5566,G5567,G5568,G5569,G5570,G5571,G5572,G5573,G5574,G5575,G5576,G5577,G5578,G5579,G5580,
       G5581,G5582,G5583,G5584,G5585,G5586,G5587,G5588,G5589,G5590,G5591,G5592,G5593,G5594,G5595,G5596,G5597,G5598,G5599,G5600,
       G5601,G5602,G5603,G5604,G5605,G5606,G5607,G5608,G5609,G5610,G5611,G5612,G5613,G5614,G5615,G5616,G5617,G5618,G5619,G5620,
       G5621,G5622,G5623,G5624,G5625,G5626,G5627,G5628,G5629,G5630,G5631,G5632,G5633,G5634,G5635,G5636,G5637,G5638,G5639,G5640,
       G5641,G5642,G5643,G5644,G5645,G5646,G5647,G5648,G5649,G5650,G5651,G5652,G5653,G5654,G5655,G5656,G5657,G5658,G5659,G5660,
       G5661,G5662,G5663,G5664,G5665,G5666,G5667,G5668,G5669,G5670,G5671,G5672,G5673,G5674,G5675,G5676,G5677,G5678,G5679,G5680,
       G5681,G5682,G5683,G5684,G5685,G5686,G5687,G5688,G5689,G5690,G5691,G5692,G5693,G5694,G5695,G5696,G5697,G5698,G5699,G5700,
       G5701,G5702,G5703,G5704,G5705,G5706,G5707,G5708,G5709,G5710,G5711,G5712,G5713,G5714,G5715,G5716,G5717,G5718,G5719,G5720,
       G5721,G5722,G5723,G5724,G5725,G5726,G5727,G5728,G5729,G5730,G5731,G5732,G5733,G5734,G5735,G5736,G5737,G5738,G5739,G5740,
       G5741,G5742,G5743,G5744,G5745,G5746,G5747,G5748,G5749,G5750,G5751,G5752,G5753,G5754,G5755,G5756,G5757,G5758,G5759,G5760,
       G5761,G5762,G5763,G5764,G5765,G5766,G5767,G5768,G5769,G5770,G5771,G5772,G5773,G5774,G5775,G5776,G5777,G5778,G5779,G5780,
       G5781,G5782,G5783,G5784,G5785,G5786,G5787,G5788,G5789,G5790,G5791,G5792,G5793,G5794,G5795,G5796,G5797,G5798,G5799,G5800,
       G5801,G5802,G5803,G5804,G5805,G5806,G5807,G5808,G5809,G5810,G5811,G5812,G5813,G5814,G5815,G5816,G5817,G5818,G5819,G5820,
       G5821,G5822,G5823,G5824,G5825,G5826,G5827,G5828,G5829,G5830,G5831,G5832,G5833,G5834,G5835,G5836,G5837,G5838,G5839,G5840,
       G5841,G5842,G5843,G5844,G5845,G5846,G5847,G5848,G5849,G5850,G5851,G5852,G5853,G5854,G5855,G5856,G5857,G5858,G5859,G5860,
       G5861,G5862,G5863,G5864,G5865,G5866,G5867,G5868,G5869,G5870,G5871,G5872,G5873,G5874,G5875,G5876,G5877,G5878,G5879,G5880,
       G5881,G5882,G5883,G5884,G5885,G5886,G5887,G5888,G5889,G5890,G5891,G5892,G5893,G5894,G5895,G5896,G5897,G5898,G5899,G5900,
       G5901,G5902,G5903,G5904,G5905,G5906,G5907,G5908,G5909,G5910,G5911,G5912,G5913,G5914,G5915,G5916,G5917,G5918,G5919,G5920,
       G5921,G5922,G5923,G5924,G5925,G5926,G5927,G5928,G5929,G5930,G5931,G5932,G5933,G5934,G5935,G5936,G5937,G5938,G5939,G5940,
       G5941,G5942,G5943,G5944,G5945,G5946,G5947,G5948,G5949,G5950,G5951,G5952,G5953,G5954,G5955,G5956,G5957,G5958,G5959,G5960,
       G5961,G5962,G5963,G5964,G5965,G5966,G5967,G5968,G5969,G5970,G5971,G5972,G5973,G5974,G5975,G5976,G5977,G5978,G5979,G5980,
       G5981,G5982,G5983,G5984,G5985,G5986,G5987,G5988,G5989,G5990,G5991,G5992,G5993,G5994,G5995,G5996,G5997,G5998,G5999,G6000,
       G6001,G6002,G6003,G6004,G6005,G6006,G6007,G6008,G6009,G6010,G6011,G6012,G6013,G6014,G6015,G6016,G6017,G6018,G6019,G6020,
       G6021,G6022,G6023,G6024,G6025,G6026,G6027,G6028,G6029,G6030,G6031,G6032,G6033,G6034,G6035,G6036,G6037,G6038,G6039,G6040,
       G6041,G6042,G6043,G6044,G6045,G6046,G6047,G6048,G6049,G6050,G6051,G6052,G6053,G6054,G6055,G6056,G6057,G6058,G6059,G6060,
       G6061,G6062,G6063,G6064,G6065,G6066,G6067,G6068,G6069,G6070,G6071,G6072,G6073,G6074,G6075,G6076,G6077,G6078,G6079,G6080,
       G6081,G6082,G6083,G6084,G6085,G6086,G6087,G6088,G6089,G6090,G6091,G6092,G6093,G6094,G6095,G6096,G6097,G6098,G6099,G6100,
       G6101,G6102,G6103,G6104,G6105,G6106,G6107,G6108,G6109,G6110,G6111,G6112,G6113,G6114,G6115,G6116,G6117,G6118,G6119,G6120,
       G6121,G6122,G6123,G6124,G6125,G6126,G6127,G6128,G6129,G6130,G6131,G6132,G6133,G6134,G6135,G6136,G6137,G6138,G6139,G6140,
       G6141,G6142,G6143,G6144,G6145,G6146,G6147,G6148,G6149,G6150,G6151,G6152,G6153,G6154,G6155,G6156,G6157,G6158,G6159,G6160,
       G6161,G6162,G6163,G6164,G6165,G6166,G6167,G6168,G6169,G6170,G6171,G6172,G6173,G6174,G6175,G6176,G6177,G6178,G6179,G6180,
       G6181,G6182,G6183,G6184,G6185,G6186,G6187,G6188,G6189,G6190,G6191,G6192,G6193,G6194,G6195,G6196,G6197,G6198,G6199,G6200,
       G6201,G6202,G6203,G6204,G6205,G6206,G6207,G6208,G6209,G6210,G6211,G6212,G6213,G6214,G6215,G6216,G6217,G6218,G6219,G6220,
       G6221,G6222,G6223,G6224,G6225,G6226,G6227,G6228,G6229,G6230,G6231,G6232,G6233,G6234,G6235,G6236,G6237,G6238,G6239,G6240,
       G6241,G6242,G6243,G6244,G6245,G6246,G6247,G6248,G6249,G6250,G6251,G6252,G6253,G6254,G6255,G6256,G6257,G6258,G6259,G6260,
       G6261,G6262,G6263,G6264,G6265,G6266,G6267,G6268,G6269,G6270,G6271,G6272,G6273,G6274,G6275,G6276,G6277,G6278,G6279,G6280,
       G6281,G6282,G6283,G6284,G6285,G6286,G6287,G6288,G6289,G6290,G6291,G6292,G6293,G6294,G6295,G6296,G6297,G6298,G6299,G6300,
       G6301,G6302,G6303,G6304,G6305,G6306,G6307,G6308,G6309,G6310,G6311,G6312,G6313,G6314,G6315,G6316,G6317,G6318,G6319,G6320,
       G6321,G6322,G6323,G6324,G6325,G6326,G6327,G6328,G6329,G6330,G6331,G6332,G6333,G6334,G6335,G6336,G6337,G6338,G6339,G6340,
       G6341,G6342,G6343,G6344,G6345,G6346,G6347,G6348,G6349,G6350,G6351,G6352,G6353,G6354,G6355,G6356,G6357,G6358,G6359,G6360,
       G6361,G6362,G6363,G6364,G6365,G6366,G6367,G6368,G6369,G6370,G6371,G6372,G6373,G6374,G6375,G6376,G6377,G6378,G6379,G6380,
       G6381,G6382,G6383,G6384,G6385,G6386,G6387,G6388,G6389,G6390,G6391,G6392,G6393,G6394,G6395,G6396,G6397,G6398,G6399,G6400,
       G6401,G6402,G6403,G6404,G6405,G6406,G6407,G6408,G6409,G6410,G6411,G6412,G6413,G6414,G6415,G6416,G6417,G6418,G6419,G6420,
       G6421,G6422,G6423,G6424,G6425,G6426,G6427,G6428,G6429,G6430,G6431,G6432,G6433,G6434,G6435,G6436,G6437,G6438,G6439,G6440,
       G6441,G6442,G6443,G6444,G6445,G6446,G6447,G6448,G6449,G6450,G6451,G6452,G6453,G6454,G6455,G6456,G6457,G6458,G6459,G6460,
       G6461,G6462,G6463,G6464,G6465,G6466,G6467,G6468,G6469,G6470,G6471,G6472,G6473,G6474,G6475,G6476,G6477,G6478,G6479,G6480,
       G6481,G6482,G6483,G6484,G6485,G6486,G6487,G6488,G6489,G6490,G6491,G6492,G6493,G6494,G6495,G6496,G6497,G6498,G6499,G6500,
       G6501,G6502,G6503,G6504,G6505,G6506,G6507,G6508,G6509,G6510,G6511,G6512,G6513,G6514,G6515,G6516,G6517,G6518,G6519,G6520,
       G6521,G6522,G6523,G6524,G6525,G6526,G6527,G6528,G6529,G6530,G6531,G6532,G6533,G6534,G6535,G6536,G6537,G6538,G6539,G6540,
       G6541,G6542,G6543,G6544,G6545,G6546,G6547,G6548,G6549,G6550,G6551,G6552,G6553,G6554,G6555,G6556,G6557,G6558,G6559,G6560,
       G6561,G6562,G6563,G6564,G6565,G6566,G6567,G6568,G6569,G6570,G6571,G6572,G6573,G6574,G6575,G6576,G6577,G6578,G6579,G6580,
       G6581,G6582,G6583,G6584,G6585,G6586,G6587,G6588,G6589,G6590,G6591,G6592,G6593,G6594,G6595,G6596,G6597,G6598,G6599,G6600,
       G6601,G6602,G6603,G6604,G6605,G6606,G6607,G6608,G6609,G6610,G6611,G6612,G6613,G6614,G6615,G6616,G6617,G6618,G6619,G6620,
       G6621,G6622,G6623,G6624,G6625,G6626,G6627,G6628,G6629,G6630,G6631,G6632,G6633,G6634,G6635,G6636,G6637,G6638,G6639,G6640,
       G6641,G6642,G6643,G6644,G6645,G6646,G6647,G6648,G6649,G6650,G6651,G6652,G6653,G6654,G6655,G6656,G6657,G6658,G6659,G6660,
       G6661,G6662,G6663,G6664,G6665,G6666,G6667,G6668,G6669,G6670,G6671,G6672,G6673,G6674,G6675,G6676,G6677,G6678,G6679,G6680,
       G6681,G6682,G6683,G6684,G6685,G6686,G6687,G6688,G6689,G6690,G6691,G6692,G6693,G6694,G6695,G6696,G6697,G6698,G6699,G6700,
       G6701,G6702,G6703,G6704,G6705,G6706,G6707,G6708,G6709,G6710,G6711,G6712,G6713,G6714,G6715,G6716,G6717,G6718,G6719,G6720,
       G6721,G6722,G6723,G6724,G6725,G6726,G6727,G6728,G6729,G6730,G6731,G6732,G6733,G6734,G6735,G6736,G6737,G6738,G6739,G6740,
       G6741,G6742,G6743,G6744,G6745,G6746,G6747,G6748,G6749,G6750,G6751,G6752,G6753,G6754,G6755,G6756,G6757,G6758,G6759,G6760,
       G6761,G6762,G6763,G6764,G6765,G6766,G6767,G6768,G6769,G6770,G6771,G6772,G6773,G6774,G6775,G6776,G6777,G6778,G6779,G6780,
       G6781,G6782,G6783,G6784,G6785,G6786,G6787,G6788,G6789,G6790,G6791,G6792,G6793,G6794,G6795,G6796,G6797,G6798,G6799,G6800,
       G6801,G6802,G6803,G6804,G6805,G6806,G6807,G6808,G6809,G6810,G6811,G6812,G6813,G6814,G6815,G6816,G6817,G6818,G6819,G6820,
       G6821,G6822,G6823,G6824,G6825,G6826,G6827,G6828,G6829,G6830,G6831,G6832,G6833,G6834,G6835,G6836,G6837,G6838,G6839,G6840,
       G6841,G6842,G6843,G6844,G6845,G6846,G6847,G6848,G6849,G6850,G6851,G6852,G6853,G6854,G6855,G6856,G6857,G6858,G6859,G6860,
       G6861,G6862,G6863,G6864,G6865,G6866,G6867,G6868,G6869,G6870,G6871,G6872,G6873,G6874,G6875,G6876,G6877,G6878,G6879,G6880,
       G6881,G6882,G6883,G6884,G6885,G6886,G6887,G6888,G6889,G6890,G6891,G6892,G6893,G6894,G6895,G6896,G6897,G6898,G6899,G6900,
       G6901,G6902,G6903,G6904,G6905,G6906,G6907,G6908,G6909,G6910,G6911,G6912,G6913,G6914,G6915,G6916,G6917,G6918,G6919,G6920,
       G6921,G6922,G6923,G6924,G6925,G6926,G6927,G6928,G6929,G6930,G6931,G6932,G6933,G6934,G6935,G6936,G6937,G6938,G6939,G6940,
       G6941,G6942,G6943,G6944,G6945,G6946,G6947,G6948,G6949,G6950,G6951,G6952,G6953,G6954,G6955,G6956,G6957,G6958,G6959,G6960,
       G6961,G6962,G6963,G6964,G6965,G6966,G6967,G6968,G6969,G6970,G6971,G6972,G6973,G6974,G6975,G6976,G6977,G6978,G6979,G6980,
       G6981,G6982,G6983,G6984,G6985,G6986,G6987,G6988,G6989,G6990,G6991,G6992,G6993,G6994,G6995,G6996,G6997,G6998,G6999,G7000,
       G7001,G7002,G7003,G7004,G7005,G7006,G7007,G7008,G7009,G7010,G7011,G7012,G7013,G7014,G7015,G7016,G7017,G7018,G7019,G7020,
       G7021,G7022,G7023,G7024,G7025,G7026,G7027,G7028,G7029,G7030,G7031,G7032,G7033,G7034,G7035,G7036,G7037,G7038,G7039,G7040,
       G7041,G7042,G7043,G7044,G7045,G7046,G7047,G7048,G7049,G7050,G7051,G7052,G7053,G7054,G7055,G7056,G7057,G7058,G7059,G7060,
       G7061,G7062,G7063,G7064,G7065,G7066,G7067,G7068,G7069,G7070,G7071,G7072,G7073,G7074,G7075,G7076,G7077,G7078,G7079,G7080,
       G7081,G7082,G7083,G7084,G7085,G7086,G7087,G7088,G7089,G7090,G7091,G7092,G7093,G7094,G7095,G7096,G7097,G7098,G7099,G7100,
       G7101,G7102,G7103,G7104,G7105,G7106,G7107,G7108,G7109,G7110,G7111,G7112,G7113,G7114,G7115,G7116,G7117,G7118,G7119,G7120,
       G7121,G7122,G7123,G7124,G7125,G7126,G7127,G7128,G7129,G7130,G7131,G7132,G7133,G7134,G7135,G7136,G7137,G7138,G7139,G7140,
       G7141,G7142,G7143,G7144,G7145,G7146,G7147,G7148,G7149,G7150,G7151,G7152,G7153,G7154,G7155,G7156,G7157,G7158,G7159,G7160,
       G7161,G7162,G7163,G7164,G7165,G7166,G7167,G7168,G7169,G7170,G7171,G7172,G7173,G7174,G7175,G7176,G7177,G7178,G7179,G7180,
       G7181,G7182,G7183,G7184,G7185,G7186,G7187,G7188,G7189,G7190,G7191,G7192,G7193,G7194,G7195,G7196,G7197,G7198,G7199,G7200,
       G7201,G7202,G7203,G7204,G7205,G7206,G7207,G7208,G7209,G7210,G7211,G7212,G7213,G7214,G7215,G7216,G7217,G7218,G7219,G7220,
       G7221,G7222,G7223,G7224,G7225,G7226,G7227,G7228,G7229,G7230,G7231,G7232,G7233,G7234,G7235,G7236,G7237,G7238,G7239,G7240,
       G7241,G7242,G7243,G7244,G7245,G7246,G7247,G7248,G7249,G7250,G7251,G7252,G7253,G7254,G7255,G7256,G7257,G7258,G7259,G7260,
       G7261,G7262,G7263,G7264,G7265,G7266,G7267,G7268,G7269,G7270,G7271,G7272,G7273,G7274,G7275,G7276,G7277,G7278,G7279,G7280,
       G7281,G7282,G7283,G7284,G7285,G7286,G7287,G7288,G7289,G7290,G7291,G7292,G7293,G7294,G7295,G7296,G7297,G7298,G7299,G7300,
       G7301,G7302,G7303,G7304,G7305,G7306,G7307,G7308,G7309,G7310,G7311,G7312,G7313,G7314,G7315,G7316,G7317,G7318,G7319,G7320,
       G7321,G7322,G7323,G7324,G7325,G7326,G7327,G7328,G7329,G7330,G7331,G7332,G7333,G7334,G7335,G7336,G7337,G7338,G7339,G7340,
       G7341,G7342,G7343,G7344,G7345,G7346,G7347,G7348,G7349,G7350,G7351,G7352,G7353,G7354,G7355,G7356,G7357,G7358,G7359,G7360,
       G7361,G7362,G7363,G7364,G7365,G7366,G7367,G7368,G7369,G7370,G7371,G7372,G7373,G7374,G7375,G7376,G7377,G7378,G7379,G7380,
       G7381,G7382,G7383,G7384,G7385,G7386,G7387,G7388,G7389,G7390,G7391,G7392,G7393,G7394,G7395,G7396,G7397,G7398,G7399,G7400,
       G7401,G7402,G7403,G7404,G7405,G7406,G7407,G7408,G7409,G7410,G7411,G7412,G7413,G7414,G7415,G7416,G7417,G7418,G7419,G7420,
       G7421,G7422,G7423,G7424,G7425,G7426,G7427,G7428,G7429,G7430,G7431,G7432,G7433,G7434,G7435,G7436,G7437,G7438,G7439,G7440,
       G7441,G7442,G7443,G7444,G7445,G7446,G7447,G7448,G7449,G7450,G7451,G7452,G7453,G7454,G7455,G7456,G7457,G7458,G7459,G7460,
       G7461,G7462,G7463,G7464,G7465,G7466,G7467,G7468,G7469,G7470,G7471,G7472,G7473,G7474,G7475,G7476,G7477,G7478,G7479,G7480,
       G7481,G7482,G7483,G7484,G7485,G7486,G7487,G7488,G7489,G7490,G7491,G7492,G7493,G7494,G7495,G7496,G7497,G7498,G7499,G7500,
       G7501,G7502,G7503,G7504,G7505,G7506,G7507,G7508,G7509,G7510,G7511,G7512,G7513,G7514,G7515,G7516,G7517,G7518,G7519,G7520,
       G7521,G7522,G7523,G7524,G7525,G7526,G7527,G7528,G7529,G7530,G7531,G7532,G7533,G7534,G7535,G7536,G7537,G7538,G7539,G7540,
       G7541,G7542,G7543,G7544,G7545,G7546,G7547,G7548,G7549,G7550,G7551,G7552,G7553,G7554,G7555,G7556,G7557,G7558,G7559,G7560,
       G7561,G7562,G7563,G7564,G7565,G7566,G7567,G7568,G7569,G7570,G7571,G7572,G7573,G7574,G7575,G7576,G7577,G7578,G7579,G7580,
       G7581,G7582,G7583,G7584,G7585,G7586,G7587,G7588,G7589,G7590,G7591,G7592,G7593,G7594,G7595,G7596,G7597,G7598,G7599,G7600,
       G7601,G7602,G7603,G7604,G7605,G7606,G7607,G7608,G7609,G7610,G7611,G7612,G7613,G7614,G7615,G7616,G7617,G7618,G7619,G7620,
       G7621,G7622,G7623,G7624,G7625,G7626,G7627,G7628,G7629,G7630,G7631,G7632,G7633,G7634,G7635,G7636,G7637,G7638,G7639,G7640,
       G7641,G7642,G7643,G7644,G7645,G7646,G7647,G7648,G7649,G7650,G7651,G7652,G7653,G7654,G7655,G7656,G7657,G7658,G7659,G7660,
       G7661,G7662,G7663,G7664,G7665,G7666,G7667,G7668,G7669,G7670,G7671,G7672,G7673,G7674,G7675,G7676,G7677,G7678,G7679,G7680,
       G7681,G7682,G7683,G7684,G7685,G7686,G7687,G7688,G7689,G7690,G7691,G7692,G7693,G7694,G7695,G7696,G7697,G7698,G7699,G7700,
       G7701,G7702,G7703,G7704,G7705,G7706,G7707,G7708,G7709,G7710,G7711,G7712,G7713,G7714,G7715,G7716,G7717,G7718,G7719,G7720,
       G7721,G7722,G7723,G7724,G7725,G7726,G7727,G7728,G7729,G7730,G7731,G7732,G7733,G7734,G7735,G7736,G7737,G7738,G7739,G7740,
       G7741,G7742,G7743,G7744,G7745,G7746,G7747,G7748,G7749,G7750,G7751,G7752,G7753,G7754,G7755,G7756,G7757,G7758,G7759,G7760,
       G7761,G7762,G7763,G7764,G7765,G7766,G7767,G7768,G7769,G7770,G7771,G7772,G7773,G7774,G7775,G7776,G7777,G7778,G7779,G7780,
       G7781,G7782,G7783,G7784,G7785,G7786,G7787,G7788,G7789,G7790,G7791,G7792,G7793,G7794,G7795,G7796,G7797,G7798,G7799,G7800,
       G7801,G7802,G7803,G7804,G7805,G7806,G7807,G7808,G7809,G7810,G7811,G7812,G7813,G7814,G7815,G7816,G7817,G7818,G7819,G7820,
       G7821,G7822,G7823,G7824,G7825,G7826,G7827,G7828,G7829,G7830,G7831,G7832,G7833,G7834,G7835,G7836,G7837,G7838,G7839,G7840,
       G7841,G7842,G7843,G7844,G7845,G7846,G7847,G7848,G7849,G7850,G7851,G7852,G7853,G7854,G7855,G7856,G7857,G7858,G7859,G7860,
       G7861,G7862,G7863,G7864,G7865,G7866,G7867,G7868,G7869,G7870,G7871,G7872,G7873,G7874,G7875,G7876,G7877,G7878,G7879,G7880,
       G7881,G7882,G7883,G7884,G7885,G7886,G7887,G7888,G7889,G7890,G7891,G7892,G7893,G7894,G7895,G7896,G7897,G7898,G7899,G7900,
       G7901,G7902,G7903,G7904,G7905,G7906,G7907,G7908,G7909,G7910,G7911,G7912,G7913,G7914,G7915,G7916,G7917,G7918,G7919,G7920,
       G7921,G7922,G7923,G7924,G7925,G7926,G7927,G7928,G7929,G7930,G7931,G7932,G7933,G7934,G7935,G7936,G7937,G7938,G7939,G7940,
       G7941,G7942,G7943,G7944,G7945,G7946,G7947,G7948,G7949,G7950,G7951,G7952,G7953,G7954,G7955,G7956,G7957,G7958,G7959,G7960,
       G7961,G7962,G7963,G7964,G7965,G7966,G7967,G7968,G7969,G7970,G7971,G7972,G7973,G7974,G7975,G7976,G7977,G7978,G7979,G7980,
       G7981,G7982,G7983,G7984,G7985,G7986,G7987,G7988,G7989,G7990,G7991,G7992,G7993,G7994,G7995,G7996,G7997,G7998,G7999,G8000,
       G8001,G8002,G8003,G8004,G8005,G8006,G8007,G8008,G8009,G8010,G8011,G8012,G8013,G8014,G8015,G8016,G8017,G8018,G8019,G8020,
       G8021,G8022,G8023,G8024,G8025,G8026,G8027,G8028,G8029,G8030,G8031,G8032,G8033,G8034,G8035,G8036,G8037,G8038,G8039,G8040,
       G8041,G8042,G8043,G8044,G8045,G8046,G8047,G8048,G8049,G8050,G8051,G8052,G8053,G8054,G8055,G8056,G8057,G8058,G8059,G8060,
       G8061,G8062,G8063,G8064,G8065,G8066,G8067,G8068,G8069,G8070,G8071,G8072,G8073,G8074,G8075,G8076,G8077,G8078,G8079,G8080,
       G8081,G8082,G8083,G8084,G8085,G8086,G8087,G8088,G8089,G8090,G8091,G8092,G8093,G8094,G8095,G8096,G8097,G8098,G8099,G8100,
       G8101,G8102,G8103,G8104,G8105,G8106,G8107,G8108,G8109,G8110,G8111,G8112,G8113,G8114,G8115,G8116,G8117,G8118,G8119,G8120,
       G8121,G8122,G8123,G8124,G8125,G8126,G8127,G8128,G8129,G8130,G8131,G8132,G8133,G8134,G8135,G8136,G8137,G8138,G8139,G8140,
       G8141,G8142,G8143,G8144,G8145,G8146,G8147,G8148,G8149,G8150,G8151,G8152,G8153,G8154,G8155,G8156,G8157,G8158,G8159,G8160,
       G8161,G8162,G8163,G8164,G8165,G8166,G8167,G8168,G8169,G8170,G8171,G8172,G8173,G8174,G8175,G8176,G8177,G8178,G8179,G8180,
       G8181,G8182,G8183,G8184,G8185,G8186,G8187,G8188,G8189,G8190,G8191,G8192,G8193,G8194,G8195,G8196,G8197,G8198,G8199,G8200,
       G8201,G8202,G8203,G8204,G8205,G8206,G8207,G8208,G8209,G8210,G8211,G8212,G8213,G8214,G8215,G8216,G8217,G8218,G8219,G8220,
       G8221,G8222,G8223,G8224,G8225,G8226,G8227,G8228,G8229,G8230,G8231,G8232,G8233,G8234,G8235,G8236,G8237,G8238,G8239,G8240,
       G8241,G8242,G8243,G8244,G8245,G8246,G8247,G8248,G8249,G8250,G8251,G8252,G8253,G8254,G8255,G8256,G8257,G8258,G8259,G8260,
       G8261,G8262,G8263,G8264,G8265,G8266,G8267,G8268,G8269,G8270,G8271,G8272,G8273,G8274,G8275,G8276,G8277,G8278,G8279,G8280,
       G8281,G8282,G8283,G8284,G8285,G8286,G8287,G8288,G8289,G8290,G8291,G8292,G8293,G8294,G8295,G8296,G8297,G8298,G8299,G8300,
       G8301,G8302,G8303,G8304,G8305,G8306,G8307,G8308,G8309,G8310,G8311,G8312,G8313,G8314,G8315,G8316,G8317,G8318,G8319,G8320,
       G8321,G8322,G8323,G8324,G8325,G8326,G8327,G8328,G8329,G8330,G8331,G8332,G8333,G8334,G8335,G8336,G8337,G8338,G8339,G8340,
       G8341,G8342,G8343,G8344,G8345,G8346,G8347,G8348,G8349,G8350,G8351,G8352,G8353,G8354,G8355,G8356,G8357,G8358,G8359,G8360,
       G8361,G8362,G8363,G8364,G8365,G8366,G8367,G8368,G8369,G8370,G8371,G8372,G8373,G8374,G8375,G8376,G8377,G8378,G8379,G8380,
       G8381,G8382,G8383,G8384,G8385,G8386,G8387,G8388,G8389,G8390,G8391,G8392,G8393,G8394,G8395,G8396,G8397,G8398,G8399,G8400,
       G8401,G8402,G8403,G8404,G8405,G8406,G8407,G8408,G8409,G8410,G8411,G8412,G8413,G8414,G8415,G8416,G8417,G8418,G8419,G8420,
       G8421,G8422,G8423,G8424,G8425,G8426,G8427,G8428,G8429,G8430,G8431,G8432,G8433,G8434,G8435,G8436,G8437,G8438,G8439,G8440,
       G8441,G8442,G8443,G8444,G8445,G8446,G8447,G8448,G8449,G8450,G8451,G8452,G8453,G8454,G8455,G8456,G8457,G8458,G8459,G8460,
       G8461,G8462,G8463,G8464,G8465,G8466,G8467,G8468,G8469,G8470,G8471,G8472,G8473,G8474,G8475,G8476,G8477,G8478,G8479,G8480,
       G8481,G8482,G8483,G8484,G8485,G8486,G8487,G8488,G8489,G8490,G8491,G8492,G8493,G8494,G8495,G8496,G8497,G8498,G8499,G8500,
       G8501,G8502,G8503,G8504,G8505,G8506,G8507,G8508,G8509,G8510,G8511,G8512,G8513,G8514,G8515,G8516,G8517,G8518,G8519,G8520,
       G8521,G8522,G8523,G8524,G8525,G8526,G8527,G8528,G8529,G8530,G8531,G8532,G8533,G8534,G8535,G8536,G8537,G8538,G8539,G8540,
       G8541,G8542,G8543,G8544,G8545,G8546,G8547,G8548,G8549,G8550,G8551,G8552,G8553,G8554,G8555,G8556,G8557,G8558,G8559,G8560,
       G8561,G8562,G8563,G8564,G8565,G8566,G8567,G8568,G8569,G8570,G8571,G8572,G8573,G8574,G8575,G8576,G8577,G8578,G8579,G8580,
       G8581,G8582,G8583,G8584,G8585,G8586,G8587,G8588,G8589,G8590,G8591,G8592,G8593,G8594,G8595,G8596,G8597,G8598,G8599,G8600,
       G8601,G8602,G8603,G8604,G8605,G8606,G8607,G8608,G8609,G8610,G8611,G8612,G8613,G8614,G8615,G8616,G8617,G8618,G8619,G8620,
       G8621,G8622,G8623,G8624,G8625,G8626,G8627,G8628,G8629,G8630,G8631,G8632,G8633,G8634,G8635,G8636,G8637,G8638,G8639,G8640,
       G8641,G8642,G8643,G8644,G8645,G8646,G8647,G8648,G8649,G8650,G8651,G8652,G8653,G8654,G8655,G8656,G8657,G8658,G8659,G8660,
       G8661,G8662,G8663,G8664,G8665,G8666,G8667,G8668,G8669,G8670,G8671,G8672,G8673,G8674,G8675,G8676,G8677,G8678,G8679,G8680,
       G8681,G8682,G8683,G8684,G8685,G8686,G8687,G8688,G8689,G8690,G8691,G8692,G8693,G8694,G8695,G8696,G8697,G8698,G8699,G8700,
       G8701,G8702,G8703,G8704,G8705,G8706,G8707,G8708,G8709,G8710,G8711,G8712,G8713,G8714,G8715,G8716,G8717,G8718,G8719,G8720,
       G8721,G8722,G8723,G8724,G8725,G8726,G8727,G8728,G8729,G8730,G8731,G8732,G8733,G8734,G8735,G8736,G8737,G8738,G8739,G8740,
       G8741,G8742,G8743,G8744,G8745,G8746,G8747,G8748,G8749,G8750,G8751,G8752,G8753,G8754,G8755,G8756,G8757,G8758,G8759,G8760,
       G8761,G8762,G8763,G8764,G8765,G8766,G8767,G8768,G8769,G8770,G8771,G8772,G8773,G8774,G8775,G8776,G8777,G8778,G8779,G8780,
       G8781,G8782,G8783,G8784,G8785,G8786,G8787,G8788,G8789,G8790,G8791,G8792,G8793,G8794,G8795,G8796,G8797,G8798,G8799,G8800,
       G8801,G8802,G8803,G8804,G8805,G8806,G8807,G8808,G8809,G8810,G8811,G8812,G8813,G8814,G8815,G8816,G8817,G8818,G8819,G8820,
       G8821,G8822,G8823,G8824,G8825,G8826,G8827,G8828,G8829,G8830,G8831,G8832,G8833,G8834,G8835,G8836,G8837,G8838,G8839,G8840,
       G8841,G8842,G8843,G8844,G8845,G8846,G8847,G8848,G8849,G8850,G8851,G8852,G8853,G8854,G8855,G8856,G8857,G8858,G8859,G8860,
       G8861,G8862,G8863,G8864,G8865,G8866,G8867,G8868,G8869,G8870,G8871,G8872,G8873,G8874,G8875,G8876,G8877,G8878,G8879,G8880,
       G8881,G8882,G8883,G8884,G8885,G8886,G8887,G8888,G8889,G8890,G8891,G8892,G8893,G8894,G8895,G8896,G8897,G8898,G8899,G8900,
       G8901,G8902,G8903,G8904,G8905,G8906,G8907,G8908,G8909,G8910,G8911,G8912,G8913,G8914,G8915,G8916,G8917,G8918,G8919,G8920,
       G8921,G8922,G8923,G8924,G8925,G8926,G8927,G8928,G8929,G8930,G8931,G8932,G8933,G8934,G8935,G8936,G8937,G8938,G8939,G8940,
       G8941,G8942,G8943,G8944,G8945,G8946,G8947,G8948,G8949,G8950,G8951,G8952,G8953,G8954,G8955,G8956,G8957,G8958,G8959,G8960,
       G8961,G8962,G8963,G8964,G8965,G8966,G8967,G8968,G8969,G8970,G8971,G8972,G8973,G8974,G8975,G8976,G8977,G8978,G8979,G8980,
       G8981,G8982,G8983,G8984,G8985,G8986,G8987,G8988,G8989,G8990,G8991,G8992,G8993,G8994,G8995,G8996,G8997,G8998,G8999,G9000,
       G9001,G9002,G9003,G9004,G9005,G9006,G9007,G9008,G9009,G9010,G9011,G9012,G9013,G9014,G9015,G9016,G9017,G9018,G9019,G9020,
       G9021,G9022,G9023,G9024,G9025,G9026,G9027,G9028,G9029,G9030,G9031,G9032,G9033,G9034,G9035,G9036,G9037,G9038,G9039,G9040,
       G9041,G9042,G9043,G9044,G9045,G9046,G9047,G9048,G9049,G9050,G9051,G9052,G9053,G9054,G9055,G9056,G9057,G9058,G9059,G9060,
       G9061,G9062,G9063,G9064,G9065,G9066,G9067,G9068,G9069,G9070,G9071,G9072,G9073,G9074,G9075,G9076,G9077,G9078,G9079,G9080,
       G9081,G9082,G9083,G9084,G9085,G9086,G9087,G9088,G9089,G9090,G9091,G9092,G9093,G9094,G9095,G9096,G9097,G9098,G9099,G9100,
       G9101,G9102,G9103,G9104,G9105,G9106,G9107,G9108,G9109,G9110,G9111,G9112,G9113,G9114,G9115,G9116,G9117,G9118,G9119,G9120,
       G9121,G9122,G9123,G9124,G9125,G9126,G9127,G9128,G9129,G9130,G9131,G9132,G9133,G9134,G9135,G9136,G9137,G9138,G9139,G9140,
       G9141,G9142,G9143,G9144,G9145,G9146,G9147,G9148,G9149,G9150,G9151,G9152,G9153,G9154,G9155,G9156,G9157,G9158,G9159,G9160,
       G9161,G9162,G9163,G9164,G9165,G9166,G9167,G9168,G9169,G9170,G9171,G9172,G9173,G9174,G9175,G9176,G9177,G9178,G9179,G9180,
       G9181,G9182,G9183,G9184,G9185,G9186,G9187,G9188,G9189,G9190,G9191,G9192,G9193,G9194,G9195,G9196,G9197,G9198,G9199,G9200,
       G9201,G9202,G9203,G9204,G9205,G9206,G9207,G9208,G9209,G9210,G9211,G9212,G9213,G9214,G9215,G9216,G9217,G9218,G9219,G9220,
       G9221,G9222,G9223,G9224,G9225,G9226,G9227,G9228,G9229,G9230,G9231,G9232,G9233,G9234,G9235,G9236,G9237,G9238,G9239,G9240,
       G9241,G9242,G9243,G9244,G9245,G9246,G9247,G9248,G9249,G9250,G9251,G9252,G9253,G9254,G9255,G9256,G9257,G9258,G9259,G9260,
       G9261,G9262,G9263,G9264,G9265,G9266,G9267,G9268,G9269,G9270,G9271,G9272,G9273,G9274,G9275,G9276,G9277,G9278,G9279,G9280,
       G9281,G9282,G9283,G9284,G9285,G9286,G9287,G9288,G9289,G9290,G9291,G9292,G9293,G9294,G9295,G9296,G9297,G9298,G9299,G9300,
       G9301,G9302,G9303,G9304,G9305,G9306,G9307,G9308,G9309,G9310,G9311,G9312,G9313,G9314,G9315,G9316,G9317,G9318,G9319,G9320,
       G9321,G9322,G9323,G9324,G9325,G9326,G9327,G9328,G9329,G9330,G9331,G9332,G9333,G9334,G9335,G9336,G9337,G9338,G9339,G9340,
       G9341,G9342,G9343,G9344,G9345,G9346,G9347,G9348,G9349,G9350,G9351,G9352,G9353,G9354,G9355,G9356,G9357,G9358,G9359,G9360,
       G9361,G9362,G9363,G9364,G9365,G9366,G9367,G9368,G9369,G9370,G9371,G9372,G9373,G9374,G9375,G9376,G9377,G9378,G9379,G9380,
       G9381,G9382,G9383,G9384,G9385,G9386,G9387,G9388,G9389,G9390,G9391,G9392,G9393,G9394,G9395,G9396,G9397,G9398,G9399,G9400,
       G9401,G9402,G9403,G9404,G9405,G9406,G9407,G9408,G9409,G9410,G9411,G9412,G9413,G9414,G9415,G9416,G9417,G9418,G9419,G9420,
       G9421,G9422,G9423,G9424,G9425,G9426,G9427,G9428,G9429,G9430,G9431,G9432,G9433,G9434,G9435,G9436,G9437,G9438,G9439,G9440,
       G9441,G9442,G9443,G9444,G9445,G9446,G9447,G9448,G9449,G9450,G9451,G9452,G9453,G9454,G9455,G9456,G9457,G9458,G9459,G9460,
       G9461,G9462,G9463,G9464,G9465,G9466,G9467,G9468,G9469,G9470,G9471,G9472,G9473,G9474,G9475,G9476,G9477,G9478,G9479,G9480,
       G9481,G9482,G9483,G9484,G9485,G9486,G9487,G9488,G9489,G9490,G9491,G9492,G9493,G9494,G9495,G9496,G9497,G9498,G9499,G9500,
       G9501,G9502,G9503,G9504,G9505,G9506,G9507,G9508,G9509,G9510,G9511,G9512,G9513,G9514,G9515,G9516,G9517,G9518,G9519,G9520,
       G9521,G9522,G9523,G9524,G9525,G9526,G9527,G9528,G9529,G9530,G9531,G9532,G9533,G9534,G9535,G9536,G9537,G9538,G9539,G9540,
       G9541,G9542,G9543,G9544,G9545,G9546,G9547,G9548,G9549,G9550,G9551,G9552,G9553,G9554,G9555,G9556,G9557,G9558,G9559,G9560,
       G9561,G9562,G9563,G9564,G9565,G9566,G9567,G9568,G9569,G9570,G9571,G9572,G9573,G9574,G9575,G9576,G9577,G9578,G9579,G9580,
       G9581,G9582,G9583,G9584,G9585,G9586,G9587,G9588,G9589,G9590,G9591,G9592,G9593,G9594,G9595,G9596,G9597,G9598,G9599,G9600,
       G9601,G9602,G9603,G9604,G9605,G9606,G9607,G9608,G9609,G9610,G9611,G9612,G9613,G9614,G9615,G9616,G9617,G9618,G9619,G9620,
       G9621,G9622,G9623,G9624,G9625,G9626,G9627,G9628,G9629,G9630,G9631,G9632,G9633,G9634,G9635,G9636,G9637,G9638,G9639,G9640,
       G9641,G9642,G9643,G9644,G9645,G9646,G9647,G9648,G9649,G9650,G9651,G9652,G9653,G9654,G9655,G9656,G9657,G9658,G9659,G9660,
       G9661,G9662,G9663,G9664,G9665,G9666,G9667,G9668,G9669,G9670,G9671,G9672,G9673,G9674,G9675,G9676,G9677,G9678,G9679,G9680,
       G9681,G9682,G9683,G9684,G9685,G9686,G9687,G9688,G9689,G9690,G9691,G9692,G9693,G9694,G9695,G9696,G9697,G9698,G9699,G9700,
       G9701,G9702,G9703,G9704,G9705,G9706,G9707,G9708,G9709,G9710,G9711,G9712,G9713,G9714,G9715,G9716,G9717,G9718,G9719,G9720,
       G9721,G9722,G9723,G9724,G9725,G9726,G9727,G9728,G9729,G9730,G9731,G9732,G9733,G9734,G9735,G9736,G9737,G9738,G9739,G9740,
       G9741,G9742,G9743,G9744,G9745,G9746,G9747,G9748,G9749,G9750,G9751,G9752,G9753,G9754,G9755,G9756,G9757,G9758,G9759,G9760,
       G9761,G9762,G9763,G9764,G9765,G9766,G9767,G9768,G9769,G9770,G9771,G9772,G9773,G9774,G9775,G9776,G9777,G9778,G9779,G9780,
       G9781,G9782,G9783,G9784,G9785,G9786,G9787,G9788,G9789,G9790,G9791,G9792,G9793,G9794,G9795,G9796,G9797,G9798,G9799,G9800,
       G9801,G9802,G9803,G9804,G9805,G9806,G9807,G9808,G9809,G9810,G9811,G9812,G9813,G9814,G9815,G9816,G9817,G9818,G9819,G9820,
       G9821,G9822,G9823,G9824,G9825,G9826,G9827,G9828,G9829,G9830,G9831,G9832,G9833,G9834,G9835,G9836,G9837,G9838,G9839,G9840,
       G9841,G9842,G9843,G9844,G9845,G9846,G9847,G9848,G9849,G9850,G9851,G9852,G9853,G9854,G9855,G9856,G9857,G9858,G9859,G9860,
       G9861,G9862,G9863,G9864,G9865,G9866,G9867,G9868,G9869,G9870,G9871,G9872,G9873,G9874,G9875,G9876,G9877,G9878,G9879,G9880,
       G9881,G9882,G9883,G9884,G9885,G9886,G9887,G9888,G9889,G9890,G9891,G9892,G9893,G9894,G9895,G9896,G9897,G9898,G9899,G9900,
       G9901,G9902,G9903,G9904,G9905,G9906,G9907,G9908,G9909,G9910,G9911,G9912,G9913,G9914,G9915,G9916,G9917,G9918,G9919,G9920,
       G9921,G9922,G9923,G9924,G9925,G9926,G9927,G9928,G9929,G9930,G9931,G9932,G9933,G9934,G9935,G9936,G9937,G9938,G9939,G9940,
       G9941,G9942,G9943,G9944,G9945,G9946,G9947,G9948,G9949,G9950,G9951,G9952,G9953,G9954,G9955,G9956,G9957,G9958,G9959,G9960,
       G9961,G9962,G9963,G9964,G9965,G9966,G9967,G9968,G9969,G9970,G9971,G9972,G9973,G9974,G9975,G9976,G9977,G9978,G9979,G9980,
       G9981,G9982,G9983,G9984,G9985,G9986,G9987,G9988,G9989,G9990,G9991,G9992,G9993,G9994,G9995,G9996,G9997,G9998,G9999,G10000,
       G10001,G10002,G10003,G10004,G10005,G10006,G10007,G10008,G10009,G10010,G10011,G10012,G10013,G10014,G10015,G10016,G10017,G10018,G10019,G10020,
       G10021,G10022,G10023,G10024,G10025,G10026,G10027,G10028,G10029,G10030,G10031,G10032,G10033,G10034,G10035,G10036,G10037,G10038,G10039,G10040,
       G10041,G10042,G10043,G10044,G10045,G10046,G10047,G10048,G10049,G10050,G10051,G10052,G10053,G10054,G10055,G10056,G10057,G10058,G10059,G10060,
       G10061,G10062,G10063,G10064,G10065,G10066,G10067,G10068,G10069,G10070,G10071,G10072,G10073,G10074,G10075,G10076,G10077,G10078,G10079,G10080,
       G10081,G10082,G10083,G10084,G10085,G10086,G10087,G10088,G10089,G10090,G10091,G10092,G10093,G10094,G10095,G10096,G10097,G10098,G10099,G10100,
       G10101,G10102,G10103,G10104,G10105,G10106,G10107,G10108,G10109,G10110,G10111,G10112,G10113,G10114,G10115,G10116,G10117,G10118,G10119,G10120,
       G10121,G10122,G10123,G10124,G10125,G10126,G10127,G10128,G10129,G10130,G10131,G10132,G10133,G10134,G10135,G10136,G10137,G10138,G10139,G10140,
       G10141,G10142,G10143,G10144,G10145,G10146,G10147,G10148,G10149,G10150,G10151,G10152,G10153,G10154,G10155,G10156,G10157,G10158,G10159,G10160,
       G10161,G10162,G10163,G10164,G10165,G10166,G10167,G10168,G10169,G10170,G10171,G10172,G10173,G10174,G10175,G10176,G10177,G10178,G10179,G10180,
       G10181,G10182,G10183,G10184,G10185,G10186,G10187,G10188,G10189,G10190,G10191,G10192,G10193,G10194,G10195,G10196,G10197,G10198,G10199,G10200,
       G10201,G10202,G10203,G10204,G10205,G10206,G10207,G10208,G10209,G10210,G10211,G10212,G10213,G10214,G10215,G10216,G10217,G10218,G10219,G10220,
       G10221,G10222,G10223,G10224,G10225,G10226,G10227,G10228,G10229,G10230,G10231,G10232,G10233,G10234,G10235,G10236,G10237,G10238,G10239,G10240,
       G10241,G10242,G10243,G10244,G10245,G10246,G10247,G10248,G10249,G10250,G10251,G10252,G10253,G10254,G10255,G10256,G10257,G10258,G10259,G10260,
       G10261,G10262,G10263,G10264,G10265,G10266,G10267,G10268,G10269,G10270,G10271,G10272,G10273,G10274,G10275,G10276,G10277,G10278,G10279,G10280,
       G10281,G10282,G10283,G10284,G10285,G10286,G10287,G10288,G10289,G10290,G10291,G10292,G10293,G10294,G10295,G10296,G10297,G10298,G10299,G10300,
       G10301,G10302,G10303,G10304,G10305,G10306,G10307,G10308,G10309,G10310,G10311,G10312,G10313,G10314,G10315,G10316,G10317,G10318,G10319,G10320,
       G10321,G10322,G10323,G10324,G10325,G10326,G10327,G10328,G10329,G10330,G10331,G10332,G10333,G10334,G10335,G10336,G10337,G10338,G10339,G10340,
       G10341,G10342,G10343,G10344,G10345,G10346,G10347,G10348,G10349,G10350,G10351,G10352,G10353,G10354,G10355,G10356,G10357,G10358,G10359,G10360,
       G10361,G10362,G10363,G10364,G10365,G10366,G10367,G10368,G10369,G10370,G10371,G10372,G10373,G10374,G10375,G10376,G10377,G10378,G10379,G10380,
       G10381,G10382,G10383,G10384,G10385,G10386,G10387,G10388,G10389,G10390,G10391,G10392,G10393,G10394,G10395,G10396,G10397,G10398,G10399,G10400,
       G10401,G10402,G10403,G10404,G10405,G10406,G10407,G10408,G10409,G10410,G10411,G10412,G10413,G10414,G10415,G10416,G10417,G10418,G10419,G10420,
       G10421,G10422,G10423,G10424,G10425,G10426,G10427,G10428,G10429,G10430,G10431,G10432,G10433,G10434,G10435,G10436,G10437,G10438,G10439,G10440,
       G10441,G10442,G10443,G10444,G10445,G10446,G10447,G10448,G10449,G10450,G10451,G10452,G10453,G10454,G10455,G10456,G10457,G10458,G10459,G10460,
       G10461,G10462,G10463,G10464,G10465,G10466,G10467,G10468,G10469,G10470,G10471,G10472,G10473,G10474,G10475,G10476,G10477,G10478,G10479,G10480,
       G10481,G10482,G10483,G10484,G10485,G10486,G10487,G10488,G10489,G10490,G10491,G10492,G10493,G10494,G10495,G10496,G10497,G10498,G10499,G10500,
       G10501,G10502,G10503,G10504,G10505,G10506,G10507,G10508,G10509,G10510,G10511,G10512,G10513,G10514,G10515,G10516,G10517,G10518,G10519,G10520,
       G10521,G10522,G10523,G10524,G10525,G10526,G10527,G10528,G10529,G10530,G10531,G10532,G10533,G10534,G10535,G10536,G10537,G10538,G10539,G10540,
       G10541,G10542,G10543,G10544,G10545,G10546,G10547,G10548,G10549,G10550,G10551,G10552,G10553,G10554,G10555,G10556,G10557,G10558,G10559,G10560,
       G10561,G10562,G10563,G10564,G10565,G10566,G10567,G10568,G10569,G10570,G10571,G10572,G10573,G10574,G10575,G10576,G10577,G10578,G10579,G10580,
       G10581,G10582,G10583,G10584,G10585,G10586,G10587,G10588,G10589,G10590,G10591,G10592,G10593,G10594,G10595,G10596,G10597,G10598,G10599,G10600,
       G10601,G10602,G10603,G10604,G10605,G10606,G10607,G10608,G10609,G10610,G10611,G10612,G10613,G10614,G10615,G10616,G10617,G10618,G10619,G10620,
       G10621,G10622,G10623,G10624,G10625,G10626,G10627,G10628,G10629,G10630,G10631,G10632,G10633,G10634,G10635,G10636,G10637,G10638,G10639,G10640,
       G10641,G10642,G10643,G10644,G10645,G10646,G10647,G10648,G10649,G10650,G10651,G10652,G10653,G10654,G10655,G10656,G10657,G10658,G10659,G10660,
       G10661,G10662,G10663,G10664,G10665,G10666,G10667,G10668,G10669,G10670,G10671,G10672,G10673,G10674,G10675,G10676,G10677,G10678,G10679,G10680,
       G10681,G10682,G10683,G10684,G10685,G10686,G10687,G10688,G10689,G10690,G10691,G10692,G10693,G10694,G10695,G10696,G10697,G10698,G10699,G10700,
       G10701,G10702,G10703,G10704,G10705,G10706,G10707,G10708,G10709,G10710,G10711,G10712,G10713,G10714,G10715,G10716,G10717,G10718,G10719,G10720,
       G10721,G10722,G10723,G10724,G10725,G10726,G10727,G10728,G10729,G10730,G10731,G10732,G10733,G10734,G10735,G10736,G10737,G10738,G10739,G10740,
       G10741,G10742,G10743,G10744,G10745,G10746,G10747,G10748,G10749,G10750,G10751,G10752,G10753,G10754,G10755,G10756,G10757,G10758,G10759,G10760,
       G10761,G10762,G10763,G10764,G10765,G10766,G10767,G10768,G10769,G10770,G10771,G10772,G10773,G10774,G10775,G10776,G10777,G10778,G10779,G10780,
       G10781,G10782,G10783,G10784,G10785,G10786,G10787,G10788,G10789,G10790,G10791,G10792,G10793,G10794,G10795,G10796,G10797,G10798,G10799,G10800,
       G10801,G10802,G10803,G10804,G10805,G10806,G10807,G10808,G10809,G10810,G10811,G10812,G10813,G10814,G10815,G10816,G10817,G10818,G10819,G10820,
       G10821,G10822,G10823,G10824,G10825,G10826,G10827,G10828,G10829,G10830,G10831,G10832,G10833,G10834,G10835,G10836,G10837,G10838,G10839,G10840,
       G10841,G10842,G10843,G10844,G10845,G10846,G10847,G10848,G10849,G10850,G10851,G10852,G10853,G10854,G10855,G10856,G10857,G10858,G10859,G10860,
       G10861,G10862,G10863,G10864,G10865,G10866,G10867,G10868,G10869,G10870,G10871,G10872,G10873,G10874,G10875,G10876,G10877,G10878,G10879,G10880,
       G10881,G10882,G10883,G10884,G10885,G10886,G10887,G10888,G10889,G10890,G10891,G10892,G10893,G10894,G10895,G10896,G10897,G10898,G10899,G10900,
       G10901,G10902,G10903,G10904,G10905,G10906,G10907,G10908,G10909,G10910,G10911,G10912,G10913,G10914,G10915,G10916,G10917,G10918,G10919,G10920,
       G10921,G10922,G10923,G10924,G10925,G10926,G10927,G10928,G10929,G10930,G10931,G10932,G10933,G10934,G10935,G10936,G10937,G10938,G10939,G10940,
       G10941,G10942,G10943,G10944,G10945,G10946,G10947,G10948,G10949,G10950,G10951,G10952,G10953,G10954,G10955,G10956,G10957,G10958,G10959,G10960,
       G10961,G10962,G10963,G10964,G10965,G10966,G10967,G10968,G10969,G10970,G10971,G10972,G10973,G10974,G10975,G10976,G10977,G10978,G10979,G10980,
       G10981,G10982,G10983,G10984,G10985,G10986,G10987,G10988,G10989,G10990,G10991,G10992,G10993,G10994,G10995,G10996,G10997,G10998,G10999,G11000,
       G11001,G11002,G11003,G11004,G11005,G11006,G11007,G11008,G11009,G11010,G11011,G11012,G11013,G11014,G11015,G11016,G11017,G11018,G11019,G11020,
       G11021,G11022,G11023,G11024,G11025,G11026,G11027,G11028,G11029,G11030,G11031,G11032,G11033,G11034,G11035,G11036,G11037,G11038,G11039,G11040,
       G11041,G11042,G11043,G11044,G11045,G11046,G11047,G11048,G11049,G11050,G11051,G11052,G11053,G11054,G11055,G11056,G11057,G11058,G11059,G11060,
       G11061,G11062,G11063,G11064,G11065,G11066,G11067,G11068,G11069,G11070,G11071,G11072,G11073,G11074,G11075,G11076,G11077,G11078,G11079,G11080,
       G11081,G11082,G11083,G11084,G11085,G11086,G11087,G11088,G11089,G11090,G11091,G11092,G11093,G11094,G11095,G11096,G11097,G11098,G11099,G11100,
       G11101,G11102,G11103,G11104,G11105,G11106,G11107,G11108,G11109,G11110,G11111,G11112,G11113,G11114,G11115,G11116,G11117,G11118,G11119,G11120,
       G11121,G11122,G11123,G11124,G11125,G11126,G11127,G11128,G11129,G11130,G11131,G11132,G11133,G11134,G11135,G11136,G11137,G11138,G11139,G11140,
       G11141,G11142,G11143,G11144,G11145,G11146,G11147,G11148,G11149,G11150,G11151,G11152,G11153,G11154,G11155,G11156,G11157,G11158,G11159,G11160,
       G11161,G11162,G11163,G11164,G11165,G11166,G11167,G11168,G11169,G11170,G11171,G11172,G11173,G11174,G11175,G11176,G11177,G11178,G11179,G11180,
       G11181,G11182,G11183,G11184,G11185,G11186,G11187,G11188,G11189,G11190,G11191,G11192,G11193,G11194,G11195,G11196,G11197,G11198,G11199,G11200,
       G11201,G11202,G11203,G11204,G11205,G11206,G11207,G11208,G11209,G11210,G11211,G11212,G11213,G11214,G11215,G11216,G11217,G11218,G11219,G11220,
       G11221,G11222,G11223,G11224,G11225,G11226,G11227,G11228,G11229,G11230,G11231,G11232,G11233,G11234,G11235,G11236,G11237,G11238,G11239,G11240,
       G11241,G11242,G11243,G11244,G11245,G11246,G11247,G11248,G11249,G11250,G11251,G11252,G11253,G11254,G11255,G11256,G11257,G11258,G11259,G11260,
       G11261,G11262,G11263,G11264,G11265,G11266,G11267,G11268,G11269,G11270,G11271,G11272,G11273,G11274,G11275,G11276,G11277,G11278,G11279,G11280,
       G11281,G11282,G11283,G11284,G11285,G11286,G11287,G11288,G11289,G11290,G11291,G11292,G11293,G11294,G11295,G11296,G11297,G11298,G11299,G11300,
       G11301,G11302,G11303,G11304,G11305,G11306,G11307,G11308,G11309,G11310,G11311,G11312,G11313,G11314,G11315,G11316,G11317,G11318,G11319,G11320,
       G11321,G11322,G11323,G11324,G11325,G11326,G11327,G11328,G11329,G11330,G11331,G11332,G11333,G11334,G11335,G11336,G11337,G11338,G11339,G11340,
       G11341,G11342,G11343,G11344,G11345,G11346,G11347,G11348,G11349,G11350,G11351,G11352,G11353,G11354,G11355,G11356,G11357,G11358,G11359,G11360,
       G11361,G11362,G11363,G11364,G11365,G11366,G11367,G11368,G11369,G11370,G11371,G11372,G11373,G11374,G11375,G11376,G11377,G11378,G11379,G11380,
       G11381,G11382,G11383,G11384,G11385,G11386,G11387,G11388,G11389,G11390,G11391,G11392,G11393,G11394,G11395,G11396,G11397,G11398,G11399,G11400,
       G11401,G11402,G11403,G11404,G11405,G11406,G11407,G11408,G11409,G11410,G11411,G11412,G11413,G11414,G11415,G11416,G11417,G11418,G11419,G11420,
       G11421,G11422,G11423,G11424,G11425,G11426,G11427,G11428,G11429,G11430,G11431,G11432,G11433,G11434,G11435,G11436,G11437,G11438,G11439,G11440,
       G11441,G11442,G11443,G11444,G11445,G11446,G11447,G11448,G11449,G11450,G11451,G11452,G11453,G11454,G11455,G11456,G11457,G11458,G11459,G11460,
       G11461,G11462,G11463,G11464,G11465,G11466,G11467,G11468,G11469,G11470,G11471,G11472,G11473,G11474,G11475,G11476,G11477,G11478,G11479,G11480,
       G11481,G11482,G11483,G11484,G11485,G11486,G11487,G11488,G11489,G11490,G11491,G11492,G11493,G11494,G11495,G11496,G11497,G11498,G11499,G11500,
       G11501,G11502,G11503,G11504,G11505,G11506,G11507,G11508,G11509,G11510,G11511,G11512,G11513,G11514,G11515,G11516,G11517,G11518,G11519,G11520,
       G11521,G11522,G11523,G11524,G11525,G11526,G11527,G11528,G11529,G11530,G11531,G11532,G11533,G11534,G11535,G11536,G11537,G11538,G11539,G11540,
       G11541,G11542,G11543,G11544,G11545,G11546,G11547,G11548,G11549,G11550,G11551,G11552,G11553,G11554,G11555,G11556,G11557,G11558,G11559,G11560,
       G11561,G11562,G11563,G11564,G11565,G11566,G11567,G11568,G11569,G11570,G11571,G11572,G11573,G11574,G11575,G11576,G11577,G11578,G11579,G11580,
       G11581,G11582,G11583,G11584,G11585,G11586,G11587,G11588,G11589,G11590,G11591,G11592,G11593,G11594,G11595,G11596,G11597,G11598,G11599,G11600,
       G11601,G11602,G11603,G11604,G11605,G11606,G11607,G11608,G11609,G11610,G11611,G11612,G11613,G11614,G11615,G11616,G11617,G11618,G11619,G11620,
       G11621,G11622,G11623,G11624,G11625,G11626,G11627,G11628,G11629,G11630,G11631,G11632,G11633,G11634,G11635,G11636,G11637,G11638,G11639,G11640,
       G11641,G11642,G11643,G11644,G11645,G11646,G11647,G11648,G11649,G11650,G11651,G11652,G11653,G11654,G11655,G11656,G11657,G11658,G11659,G11660,
       G11661,G11662,G11663,G11664,G11665,G11666,G11667,G11668,G11669,G11670,G11671,G11672,G11673,G11674,G11675,G11676,G11677,G11678,G11679,G11680,
       G11681,G11682,G11683,G11684,G11685,G11686,G11687,G11688,G11689,G11690,G11691,G11692,G11693,G11694,G11695,G11696,G11697,G11698,G11699,G11700,
       G11701,G11702,G11703,G11704,G11705,G11706,G11707,G11708,G11709,G11710,G11711,G11712,G11713,G11714,G11715,G11716,G11717,G11718,G11719,G11720,
       G11721,G11722,G11723,G11724,G11725,G11726,G11727,G11728,G11729,G11730,G11731,G11732,G11733,G11734,G11735,G11736,G11737,G11738,G11739,G11740,
       G11741,G11742,G11743,G11744,G11745,G11746,G11747,G11748,G11749,G11750,G11751,G11752,G11753,G11754,G11755,G11756,G11757,G11758,G11759,G11760,
       G11761,G11762,G11763,G11764,G11765,G11766,G11767,G11768,G11769,G11770,G11771,G11772,G11773,G11774,G11775,G11776,G11777,G11778,G11779,G11780,
       G11781,G11782,G11783,G11784,G11785,G11786,G11787,G11788,G11789,G11790,G11791,G11792,G11793,G11794,G11795,G11796,G11797,G11798,G11799,G11800,
       G11801,G11802,G11803,G11804,G11805,G11806,G11807,G11808,G11809,G11810,G11811,G11812,G11813,G11814,G11815,G11816,G11817,G11818,G11819,G11820,
       G11821,G11822,G11823,G11824,G11825,G11826,G11827,G11828,G11829,G11830,G11831,G11832,G11833,G11834,G11835,G11836,G11837,G11838,G11839,G11840,
       G11841,G11842,G11843,G11844,G11845,G11846,G11847,G11848,G11849,G11850,G11851,G11852,G11853,G11854,G11855,G11856,G11857,G11858,G11859,G11860,
       G11861,G11862,G11863,G11864,G11865,G11866,G11867,G11868,G11869,G11870,G11871,G11872,G11873,G11874,G11875,G11876,G11877,G11878,G11879,G11880,
       G11881,G11882,G11883,G11884,G11885,G11886,G11887,G11888,G11889,G11890,G11891,G11892,G11893,G11894,G11895,G11896,G11897,G11898,G11899,G11900,
       G11901,G11902,G11903,G11904,G11905,G11906,G11907,G11908,G11909,G11910,G11911,G11912,G11913,G11914,G11915,G11916,G11917,G11918,G11919,G11920,
       G11921,G11922,G11923,G11924,G11925,G11926,G11927,G11928,G11929,G11930,G11931,G11932,G11933,G11934,G11935,G11936,G11937,G11938,G11939,G11940,
       G11941,G11942,G11943,G11944,G11945,G11946,G11947,G11948,G11949,G11950,G11951,G11952,G11953,G11954,G11955,G11956,G11957,G11958,G11959,G11960,
       G11961,G11962,G11963,G11964,G11965,G11966,G11967,G11968,G11969,G11970,G11971,G11972,G11973,G11974,G11975,G11976,G11977,G11978,G11979,G11980,
       G11981,G11982,G11983,G11984,G11985,G11986,G11987,G11988,G11989,G11990,G11991,G11992,G11993,G11994,G11995,G11996,G11997,G11998,G11999,G12000,
       G12001,G12002,G12003,G12004,G12005,G12006,G12007,G12008,G12009,G12010,G12011,G12012,G12013,G12014,G12015,G12016,G12017,G12018,G12019,G12020,
       G12021,G12022,G12023,G12024,G12025,G12026,G12027,G12028,G12029,G12030,G12031,G12032,G12033,G12034,G12035,G12036,G12037,G12038,G12039,G12040,
       G12041,G12042,G12043,G12044,G12045,G12046,G12047,G12048,G12049,G12050,G12051,G12052,G12053,G12054,G12055,G12056,G12057,G12058,G12059,G12060,
       G12061,G12062,G12063,G12064,G12065,G12066,G12067,G12068,G12069,G12070,G12071,G12072,G12073,G12074,G12075,G12076,G12077,G12078,G12079,G12080,
       G12081,G12082,G12083,G12084,G12085,G12086,G12087,G12088,G12089,G12090,G12091,G12092,G12093,G12094,G12095,G12096,G12097,G12098,G12099,G12100,
       G12101,G12102,G12103,G12104,G12105,G12106,G12107,G12108,G12109,G12110,G12111,G12112,G12113,G12114,G12115,G12116,G12117,G12118,G12119,G12120,
       G12121,G12122,G12123,G12124,G12125,G12126,G12127,G12128,G12129,G12130,G12131,G12132,G12133,G12134,G12135,G12136,G12137,G12138,G12139,G12140,
       G12141,G12142,G12143,G12144,G12145,G12146,G12147,G12148,G12149,G12150,G12151,G12152,G12153,G12154,G12155,G12156,G12157,G12158,G12159,G12160,
       G12161,G12162,G12163,G12164,G12165,G12166,G12167,G12168,G12169,G12170,G12171,G12172,G12173,G12174,G12175,G12176,G12177,G12178,G12179,G12180,
       G12181,G12182,G12183,G12184,G12185,G12186,G12187,G12188,G12189,G12190,G12191,G12192,G12193,G12194,G12195,G12196,G12197,G12198,G12199,G12200,
       G12201,G12202,G12203,G12204,G12205,G12206,G12207,G12208,G12209,G12210,G12211,G12212,G12213,G12214,G12215,G12216,G12217,G12218,G12219,G12220,
       G12221,G12222,G12223,G12224,G12225,G12226,G12227,G12228,G12229,G12230,G12231,G12232,G12233,G12234,G12235,G12236,G12237,G12238,G12239,G12240,
       G12241,G12242,G12243,G12244,G12245,G12246,G12247,G12248,G12249,G12250,G12251,G12252,G12253,G12254,G12255,G12256,G12257,G12258,G12259,G12260,
       G12261,G12262,G12263,G12264,G12265,G12266,G12267,G12268,G12269,G12270,G12271,G12272,G12273,G12274,G12275,G12276,G12277,G12278,G12279,G12280,
       G12281,G12282,G12283,G12284,G12285,G12286,G12287,G12288,G12289,G12290,G12291,G12292,G12293,G12294,G12295,G12296,G12297,G12298,G12299,G12300,
       G12301,G12302,G12303,G12304,G12305,G12306,G12307,G12308,G12309,G12310,G12311,G12312,G12313,G12314,G12315,G12316,G12317,G12318,G12319,G12320,
       G12321,G12322,G12323,G12324,G12325,G12326,G12327,G12328,G12329,G12330,G12331,G12332,G12333,G12334,G12335,G12336,G12337,G12338,G12339,G12340,
       G12341,G12342,G12343,G12344,G12345,G12346,G12347,G12348,G12349,G12350,G12351,G12352,G12353,G12354,G12355,G12356,G12357,G12358,G12359,G12360,
       G12361,G12362,G12363,G12364,G12365,G12366,G12367,G12368,G12369,G12370,G12371,G12372,G12373,G12374,G12375,G12376,G12377,G12378,G12379,G12380,
       G12381,G12382,G12383,G12384,G12385,G12386,G12387,G12388,G12389,G12390,G12391,G12392,G12393,G12394,G12395,G12396,G12397,G12398,G12399,G12400,
       G12401,G12402,G12403,G12404,G12405,G12406,G12407,G12408,G12409,G12410,G12411,G12412,G12413,G12414,G12415,G12416,G12417,G12418,G12419,G12420,
       G12421,G12422,G12423,G12424,G12425,G12426,G12427,G12428,G12429,G12430,G12431,G12432,G12433,G12434,G12435,G12436,G12437,G12438,G12439,G12440,
       G12441,G12442,G12443,G12444,G12445,G12446,G12447,G12448,G12449,G12450,G12451,G12452,G12453,G12454,G12455,G12456,G12457,G12458,G12459,G12460,
       G12461,G12462,G12463,G12464,G12465,G12466,G12467,G12468,G12469,G12470,G12471,G12472,G12473,G12474,G12475,G12476,G12477,G12478,G12479,G12480,
       G12481,G12482,G12483,G12484,G12485,G12486,G12487,G12488,G12489,G12490,G12491,G12492,G12493,G12494,G12495,G12496,G12497,G12498,G12499,G12500,
       G12501,G12502,G12503,G12504,G12505,G12506,G12507,G12508,G12509,G12510,G12511,G12512,G12513,G12514,G12515,G12516,G12517,G12518,G12519,G12520,
       G12521,G12522,G12523,G12524,G12525,G12526,G12527,G12528,G12529,G12530,G12531,G12532,G12533,G12534,G12535,G12536,G12537,G12538,G12539,G12540,
       G12541,G12542,G12543,G12544,G12545,G12546,G12547,G12548,G12549,G12550,G12551,G12552,G12553,G12554,G12555,G12556,G12557,G12558,G12559,G12560,
       G12561,G12562,G12563,G12564,G12565,G12566,G12567,G12568,G12569,G12570,G12571,G12572,G12573,G12574,G12575,G12576,G12577,G12578,G12579,G12580,
       G12581,G12582,G12583,G12584,G12585,G12586,G12587,G12588,G12589,G12590,G12591,G12592,G12593,G12594,G12595,G12596,G12597,G12598,G12599,G12600,
       G12601,G12602,G12603,G12604,G12605,G12606,G12607,G12608,G12609,G12610,G12611,G12612,G12613,G12614,G12615,G12616,G12617,G12618,G12619,G12620,
       G12621,G12622,G12623,G12624,G12625,G12626,G12627,G12628,G12629,G12630,G12631,G12632,G12633,G12634,G12635,G12636,G12637,G12638,G12639,G12640,
       G12641,G12642,G12643,G12644,G12645,G12646,G12647,G12648,G12649,G12650,G12651,G12652,G12653,G12654,G12655,G12656,G12657,G12658,G12659,G12660,
       G12661,G12662,G12663,G12664,G12665,G12666,G12667,G12668,G12669,G12670,G12671,G12672,G12673,G12674,G12675,G12676,G12677,G12678,G12679,G12680,
       G12681,G12682,G12683,G12684,G12685,G12686,G12687,G12688,G12689,G12690,G12691,G12692,G12693,G12694,G12695,G12696,G12697,G12698,G12699,G12700,
       G12701,G12702,G12703,G12704,G12705,G12706,G12707,G12708,G12709,G12710,G12711,G12712,G12713,G12714,G12715,G12716,G12717,G12718,G12719,G12720,
       G12721,G12722,G12723,G12724,G12725,G12726,G12727,G12728,G12729,G12730,G12731,G12732,G12733,G12734,G12735,G12736,G12737,G12738,G12739,G12740,
       G12741,G12742,G12743,G12744,G12745,G12746,G12747,G12748,G12749,G12750,G12751,G12752,G12753,G12754,G12755,G12756,G12757,G12758,G12759,G12760,
       G12761,G12762,G12763,G12764,G12765,G12766,G12767,G12768,G12769,G12770,G12771,G12772,G12773,G12774,G12775,G12776,G12777,G12778,G12779,G12780,
       G12781,G12782,G12783,G12784,G12785,G12786,G12787,G12788,G12789,G12790,G12791,G12792,G12793,G12794,G12795,G12796,G12797,G12798,G12799,G12800,
       G12801,G12802,G12803,G12804,G12805,G12806,G12807,G12808,G12809,G12810,G12811,G12812,G12813,G12814,G12815,G12816,G12817,G12818,G12819,G12820,
       G12821,G12822,G12823,G12824,G12825,G12826,G12827,G12828,G12829,G12830,G12831,G12832,G12833,G12834,G12835,G12836,G12837,G12838,G12839,G12840,
       G12841,G12842,G12843,G12844,G12845,G12846,G12847,G12848,G12849,G12850,G12851,G12852,G12853,G12854,G12855,G12856,G12857,G12858,G12859,G12860,
       G12861,G12862,G12863,G12864,G12865,G12866,G12867,G12868,G12869,G12870,G12871,G12872,G12873,G12874,G12875,G12876,G12877,G12878,G12879,G12880,
       G12881,G12882,G12883,G12884,G12885,G12886,G12887,G12888,G12889,G12890,G12891,G12892,G12893,G12894,G12895,G12896,G12897,G12898,G12899,G12900,
       G12901,G12902,G12903,G12904,G12905,G12906,G12907,G12908,G12909,G12910,G12911,G12912,G12913,G12914,G12915,G12916,G12917,G12918,G12919,G12920,
       G12921,G12922,G12923,G12924,G12925,G12926,G12927,G12928,G12929,G12930,G12931,G12932,G12933,G12934,G12935,G12936,G12937,G12938,G12939,G12940,
       G12941,G12942,G12943,G12944,G12945,G12946,G12947,G12948,G12949,G12950,G12951,G12952,G12953,G12954,G12955,G12956,G12957,G12958,G12959,G12960,
       G12961,G12962,G12963,G12964,G12965,G12966,G12967,G12968,G12969,G12970,G12971,G12972,G12973,G12974,G12975,G12976,G12977,G12978,G12979,G12980,
       G12981,G12982,G12983,G12984,G12985,G12986,G12987,G12988,G12989,G12990,G12991,G12992,G12993,G12994,G12995,G12996,G12997,G12998,G12999,G13000,
       G13001,G13002,G13003,G13004,G13005,G13006,G13007,G13008,G13009,G13010,G13011,G13012,G13013,G13014,G13015,G13016,G13017,G13018,G13019,G13020,
       G13021,G13022,G13023,G13024,G13025,G13026,G13027,G13028,G13029,G13030,G13031,G13032,G13033,G13034,G13035,G13036,G13037,G13038,G13039,G13040,
       G13041,G13042,G13043,G13044,G13045,G13046,G13047,G13048,G13049,G13050,G13051,G13052,G13053,G13054,G13055,G13056,G13057,G13058,G13059,G13060,
       G13061,G13062,G13063,G13064,G13065,G13066,G13067,G13068,G13069,G13070,G13071,G13072,G13073,G13074,G13075,G13076,G13077,G13078,G13079,G13080,
       G13081,G13082,G13083,G13084,G13085,G13086,G13087,G13088,G13089,G13090,G13091,G13092,G13093,G13094,G13095,G13096,G13097,G13098,G13099,G13100,
       G13101,G13102,G13103,G13104,G13105,G13106,G13107,G13108,G13109,G13110,G13111,G13112,G13113,G13114,G13115,G13116,G13117,G13118,G13119,G13120,
       G13121,G13122,G13123,G13124,G13125,G13126,G13127,G13128,G13129,G13130,G13131,G13132,G13133,G13134,G13135,G13136,G13137,G13138,G13139,G13140,
       G13141,G13142,G13143,G13144,G13145,G13146,G13147,G13148,G13149,G13150,G13151,G13152,G13153,G13154,G13155,G13156,G13157,G13158,G13159,G13160,
       G13161,G13162,G13163,G13164,G13165,G13166,G13167,G13168,G13169,G13170,G13171,G13172,G13173,G13174,G13175,G13176,G13177,G13178,G13179,G13180,
       G13181,G13182,G13183,G13184,G13185,G13186,G13187,G13188,G13189,G13190,G13191,G13192,G13193,G13194,G13195,G13196,G13197,G13198,G13199,G13200,
       G13201,G13202,G13203,G13204,G13205,G13206,G13207,G13208,G13209,G13210,G13211,G13212,G13213,G13214,G13215,G13216,G13217,G13218,G13219,G13220,
       G13221,G13222,G13223,G13224,G13225,G13226,G13227,G13228,G13229,G13230,G13231,G13232,G13233,G13234,G13235,G13236,G13237,G13238,G13239,G13240,
       G13241,G13242,G13243,G13244,G13245,G13246,G13247,G13248,G13249,G13250,G13251,G13252,G13253,G13254,G13255,G13256,G13257,G13258,G13259,G13260,
       G13261,G13262,G13263,G13264,G13265,G13266,G13267,G13268,G13269,G13270,G13271,G13272,G13273,G13274,G13275,G13276,G13277,G13278,G13279,G13280,
       G13281,G13282,G13283,G13284,G13285,G13286,G13287,G13288,G13289,G13290,G13291,G13292,G13293,G13294,G13295,G13296,G13297,G13298,G13299,G13300,
       G13301,G13302,G13303,G13304,G13305,G13306,G13307,G13308,G13309,G13310,G13311,G13312,G13313,G13314,G13315,G13316,G13317,G13318,G13319,G13320,
       G13321,G13322,G13323,G13324,G13325,G13326,G13327,G13328,G13329,G13330,G13331,G13332,G13333,G13334,G13335,G13336,G13337,G13338,G13339,G13340,
       G13341,G13342,G13343,G13344,G13345,G13346,G13347,G13348,G13349,G13350,G13351,G13352,G13353,G13354,G13355,G13356,G13357,G13358,G13359,G13360,
       G13361,G13362,G13363,G13364,G13365,G13366,G13367,G13368,G13369,G13370,G13371,G13372,G13373,G13374,G13375,G13376,G13377,G13378,G13379,G13380,
       G13381,G13382,G13383,G13384,G13385,G13386,G13387,G13388,G13389,G13390,G13391,G13392,G13393,G13394,G13395,G13396,G13397,G13398,G13399,G13400,
       G13401,G13402,G13403,G13404,G13405,G13406,G13407,G13408,G13409,G13410,G13411,G13412,G13413,G13414,G13415,G13416,G13417,G13418,G13419,G13420,
       G13421,G13422,G13423,G13424,G13425,G13426,G13427,G13428,G13429,G13430,G13431,G13432,G13433,G13434,G13435,G13436,G13437,G13438,G13439,G13440,
       G13441,G13442,G13443,G13444,G13445,G13446,G13447,G13448,G13449,G13450,G13451,G13452,G13453,G13454,G13455,G13456,G13457,G13458,G13459,G13460,
       G13461,G13462,G13463,G13464,G13465,G13466,G13467,G13468,G13469,G13470,G13471,G13472,G13473,G13474,G13475,G13476,G13477,G13478,G13479,G13480,
       G13481,G13482,G13483,G13484,G13485,G13486,G13487,G13488,G13489,G13490,G13491,G13492,G13493,G13494,G13495,G13496,G13497,G13498,G13499,G13500,
       G13501,G13502,G13503,G13504,G13505,G13506,G13507,G13508,G13509,G13510,G13511,G13512,G13513,G13514,G13515,G13516,G13517,G13518,G13519,G13520,
       G13521,G13522,G13523,G13524,G13525,G13526,G13527,G13528,G13529,G13530,G13531,G13532,G13533,G13534,G13535,G13536,G13537,G13538,G13539,G13540,
       G13541,G13542,G13543,G13544,G13545,G13546,G13547,G13548,G13549,G13550,G13551,G13552,G13553,G13554,G13555,G13556,G13557,G13558,G13559,G13560,
       G13561,G13562,G13563,G13564,G13565,G13566,G13567,G13568,G13569,G13570,G13571,G13572,G13573,G13574,G13575,G13576,G13577,G13578,G13579,G13580,
       G13581,G13582,G13583,G13584,G13585,G13586,G13587,G13588,G13589,G13590,G13591,G13592,G13593,G13594,G13595,G13596,G13597,G13598,G13599,G13600,
       G13601,G13602,G13603,G13604,G13605,G13606,G13607,G13608,G13609,G13610,G13611,G13612,G13613,G13614,G13615,G13616,G13617,G13618,G13619,G13620,
       G13621,G13622,G13623,G13624,G13625,G13626,G13627,G13628,G13629,G13630,G13631,G13632,G13633,G13634,G13635,G13636,G13637,G13638,G13639,G13640,
       G13641,G13642,G13643,G13644,G13645,G13646,G13647,G13648,G13649,G13650,G13651,G13652,G13653,G13654,G13655,G13656,G13657,G13658,G13659,G13660,
       G13661,G13662,G13663,G13664,G13665,G13666,G13667,G13668,G13669,G13670,G13671,G13672,G13673,G13674,G13675,G13676,G13677,G13678,G13679,G13680,
       G13681,G13682,G13683,G13684,G13685,G13686,G13687,G13688,G13689,G13690,G13691,G13692,G13693,G13694,G13695,G13696,G13697,G13698,G13699,G13700,
       G13701,G13702,G13703,G13704,G13705,G13706,G13707,G13708,G13709,G13710,G13711,G13712,G13713,G13714,G13715,G13716,G13717,G13718,G13719,G13720,
       G13721,G13722,G13723,G13724,G13725,G13726,G13727,G13728,G13729,G13730,G13731,G13732,G13733,G13734,G13735,G13736,G13737,G13738,G13739,G13740,
       G13741,G13742,G13743,G13744,G13745,G13746,G13747,G13748,G13749,G13750,G13751,G13752,G13753,G13754,G13755,G13756,G13757,G13758,G13759,G13760,
       G13761,G13762,G13763,G13764,G13765,G13766,G13767,G13768,G13769,G13770,G13771,G13772,G13773,G13774,G13775,G13776,G13777,G13778,G13779,G13780,
       G13781,G13782,G13783,G13784,G13785,G13786,G13787,G13788,G13789,G13790,G13791,G13792,G13793,G13794,G13795,G13796,G13797,G13798,G13799,G13800,
       G13801,G13802,G13803,G13804,G13805,G13806,G13807,G13808,G13809,G13810,G13811,G13812,G13813,G13814,G13815,G13816,G13817,G13818,G13819,G13820,
       G13821,G13822,G13823,G13824,G13825,G13826,G13827,G13828,G13829,G13830,G13831,G13832,G13833,G13834,G13835,G13836,G13837,G13838,G13839,G13840,
       G13841,G13842,G13843,G13844,G13845,G13846,G13847,G13848,G13849,G13850,G13851,G13852,G13853,G13854,G13855,G13856,G13857,G13858,G13859,G13860,
       G13861,G13862,G13863,G13864,G13865,G13866,G13867,G13868,G13869,G13870,G13871,G13872,G13873,G13874,G13875,G13876,G13877,G13878,G13879,G13880,
       G13881,G13882,G13883,G13884,G13885,G13886,G13887,G13888,G13889,G13890,G13891,G13892,G13893,G13894,G13895,G13896,G13897,G13898,G13899,G13900,
       G13901,G13902,G13903,G13904,G13905,G13906,G13907,G13908,G13909,G13910,G13911,G13912,G13913,G13914,G13915,G13916,G13917,G13918,G13919,G13920,
       G13921,G13922,G13923,G13924,G13925,G13926,G13927,G13928,G13929,G13930,G13931,G13932,G13933,G13934,G13935,G13936,G13937,G13938,G13939,G13940,
       G13941,G13942,G13943,G13944,G13945,G13946,G13947,G13948,G13949,G13950,G13951,G13952,G13953,G13954,G13955,G13956,G13957,G13958,G13959,G13960,
       G13961,G13962,G13963,G13964,G13965,G13966,G13967,G13968,G13969,G13970,G13971,G13972,G13973,G13974,G13975,G13976,G13977,G13978,G13979,G13980,
       G13981,G13982,G13983,G13984,G13985,G13986,G13987,G13988,G13989,G13990,G13991,G13992,G13993,G13994,G13995,G13996,G13997,G13998,G13999,G14000,
       G14001,G14002,G14003,G14004,G14005,G14006,G14007,G14008,G14009,G14010,G14011,G14012,G14013,G14014,G14015,G14016,G14017,G14018,G14019,G14020,
       G14021,G14022,G14023,G14024,G14025,G14026,G14027,G14028,G14029,G14030,G14031,G14032,G14033,G14034,G14035,G14036,G14037,G14038,G14039,G14040,
       G14041,G14042,G14043,G14044,G14045,G14046,G14047,G14048,G14049,G14050,G14051,G14052,G14053,G14054,G14055,G14056,G14057,G14058,G14059,G14060,
       G14061,G14062,G14063,G14064,G14065,G14066,G14067,G14068,G14069,G14070,G14071,G14072,G14073,G14074,G14075,G14076,G14077,G14078,G14079,G14080,
       G14081,G14082,G14083,G14084,G14085,G14086,G14087,G14088,G14089,G14090,G14091,G14092,G14093,G14094,G14095,G14096,G14097,G14098,G14099,G14100,
       G14101,G14102,G14103,G14104,G14105,G14106,G14107,G14108,G14109,G14110,G14111,G14112,G14113,G14114,G14115,G14116,G14117,G14118,G14119,G14120,
       G14121,G14122,G14123,G14124,G14125,G14126,G14127,G14128,G14129,G14130,G14131,G14132,G14133,G14134,G14135,G14136,G14137,G14138,G14139,G14140,
       G14141,G14142,G14143,G14144,G14145,G14146,G14147,G14148,G14149,G14150,G14151,G14152,G14153,G14154,G14155,G14156,G14157,G14158,G14159,G14160,
       G14161,G14162,G14163,G14164,G14165,G14166,G14167,G14168,G14169,G14170,G14171,G14172,G14173,G14174,G14175,G14176,G14177,G14178,G14179,G14180,
       G14181,G14182,G14183,G14184,G14185,G14186,G14187,G14188,G14189,G14190,G14191,G14192,G14193,G14194,G14195,G14196,G14197,G14198,G14199,G14200,
       G14201,G14202,G14203,G14204,G14205,G14206,G14207,G14208,G14209,G14210,G14211,G14212,G14213,G14214,G14215,G14216,G14217,G14218,G14219,G14220,
       G14221,G14222,G14223,G14224,G14225,G14226,G14227,G14228,G14229,G14230,G14231,G14232,G14233,G14234,G14235,G14236,G14237,G14238,G14239,G14240,
       G14241,G14242,G14243,G14244,G14245,G14246,G14247,G14248,G14249,G14250,G14251,G14252,G14253,G14254,G14255,G14256,G14257,G14258,G14259,G14260,
       G14261,G14262,G14263,G14264,G14265,G14266,G14267,G14268,G14269,G14270,G14271,G14272,G14273,G14274,G14275,G14276,G14277,G14278,G14279,G14280,
       G14281,G14282,G14283,G14284,G14285,G14286,G14287,G14288,G14289,G14290,G14291,G14292,G14293,G14294,G14295,G14296,G14297,G14298,G14299,G14300,
       G14301,G14302,G14303,G14304,G14305,G14306,G14307,G14308,G14309,G14310,G14311,G14312,G14313,G14314,G14315,G14316,G14317,G14318,G14319,G14320,
       G14321,G14322,G14323,G14324,G14325,G14326,G14327,G14328,G14329,G14330,G14331,G14332,G14333,G14334,G14335,G14336,G14337,G14338,G14339,G14340,
       G14341,G14342,G14343,G14344,G14345,G14346,G14347,G14348,G14349,G14350,G14351,G14352,G14353,G14354,G14355,G14356,G14357,G14358,G14359,G14360,
       G14361,G14362,G14363,G14364,G14365,G14366,G14367,G14368,G14369,G14370,G14371,G14372,G14373,G14374,G14375,G14376,G14377,G14378,G14379,G14380,
       G14381,G14382,G14383,G14384,G14385,G14386,G14387,G14388,G14389,G14390,G14391,G14392,G14393,G14394,G14395,G14396,G14397,G14398,G14399,G14400,
       G14401,G14402,G14403,G14404,G14405,G14406,G14407,G14408,G14409,G14410,G14411,G14412,G14413,G14414,G14415,G14416,G14417,G14418,G14419,G14420,
       G14421,G14422,G14423,G14424,G14425,G14426,G14427,G14428,G14429,G14430,G14431,G14432,G14433,G14434,G14435,G14436,G14437,G14438,G14439,G14440,
       G14441,G14442,G14443,G14444,G14445,G14446,G14447,G14448,G14449,G14450,G14451,G14452,G14453,G14454,G14455,G14456,G14457,G14458,G14459,G14460,
       G14461,G14462,G14463,G14464,G14465,G14466,G14467,G14468,G14469,G14470,G14471,G14472,G14473,G14474,G14475,G14476,G14477,G14478,G14479,G14480,
       G14481,G14482,G14483,G14484,G14485,G14486,G14487,G14488,G14489,G14490,G14491,G14492,G14493,G14494,G14495,G14496,G14497,G14498,G14499,G14500,
       G14501,G14502,G14503,G14504,G14505,G14506,G14507,G14508,G14509,G14510,G14511,G14512,G14513,G14514,G14515,G14516,G14517,G14518,G14519,G14520,
       G14521,G14522,G14523,G14524,G14525,G14526,G14527,G14528,G14529,G14530,G14531,G14532,G14533,G14534,G14535,G14536,G14537,G14538,G14539,G14540,
       G14541,G14542,G14543,G14544,G14545,G14546,G14547,G14548,G14549,G14550,G14551,G14552,G14553,G14554,G14555,G14556,G14557,G14558,G14559,G14560,
       G14561,G14562,G14563,G14564,G14565,G14566,G14567,G14568,G14569,G14570,G14571,G14572,G14573,G14574,G14575,G14576,G14577,G14578,G14579,G14580,
       G14581,G14582,G14583,G14584,G14585,G14586,G14587,G14588,G14589,G14590,G14591,G14592,G14593,G14594,G14595,G14596,G14597,G14598,G14599,G14600,
       G14601,G14602,G14603,G14604,G14605,G14606,G14607,G14608,G14609,G14610,G14611,G14612,G14613,G14614,G14615,G14616,G14617,G14618,G14619,G14620,
       G14621,G14622,G14623,G14624,G14625,G14626,G14627,G14628,G14629,G14630,G14631,G14632,G14633,G14634,G14635,G14636,G14637,G14638,G14639,G14640,
       G14641,G14642,G14643,G14644,G14645,G14646,G14647,G14648,G14649,G14650,G14651,G14652,G14653,G14654,G14655,G14656,G14657,G14658,G14659,G14660,
       G14661,G14662,G14663,G14664,G14665,G14666,G14667,G14668,G14669,G14670,G14671,G14672,G14673,G14674,G14675,G14676,G14677,G14678,G14679,G14680,
       G14681,G14682,G14683,G14684,G14685,G14686,G14687,G14688,G14689,G14690,G14691,G14692,G14693,G14694,G14695,G14696,G14697,G14698,G14699,G14700,
       G14701,G14702,G14703,G14704,G14705,G14706,G14707,G14708,G14709,G14710,G14711,G14712,G14713,G14714,G14715,G14716,G14717,G14718,G14719,G14720,
       G14721,G14722,G14723,G14724,G14725,G14726,G14727,G14728,G14729,G14730,G14731,G14732,G14733,G14734,G14735,G14736,G14737,G14738,G14739,G14740,
       G14741,G14742,G14743,G14744,G14745,G14746,G14747,G14748,G14749,G14750,G14751,G14752,G14753,G14754,G14755,G14756,G14757,G14758,G14759,G14760,
       G14761,G14762,G14763,G14764,G14765,G14766,G14767,G14768,G14769,G14770,G14771,G14772,G14773,G14774,G14775,G14776,G14777,G14778,G14779,G14780,
       G14781,G14782,G14783,G14784,G14785,G14786,G14787,G14788,G14789,G14790,G14791,G14792,G14793,G14794,G14795,G14796,G14797,G14798,G14799,G14800,
       G14801,G14802,G14803,G14804,G14805,G14806,G14807,G14808,G14809,G14810,G14811,G14812,G14813,G14814,G14815,G14816,G14817,G14818,G14819,G14820,
       G14821,G14822,G14823,G14824,G14825,G14826,G14827,G14828,G14829,G14830,G14831,G14832,G14833,G14834,G14835,G14836,G14837,G14838,G14839,G14840,
       G14841,G14842,G14843,G14844,G14845,G14846,G14847,G14848,G14849,G14850,G14851,G14852,G14853,G14854,G14855,G14856,G14857,G14858,G14859,G14860,
       G14861,G14862,G14863,G14864,G14865,G14866,G14867,G14868,G14869,G14870,G14871,G14872,G14873,G14874,G14875,G14876,G14877,G14878,G14879,G14880,
       G14881,G14882,G14883,G14884,G14885,G14886,G14887,G14888,G14889,G14890,G14891,G14892,G14893,G14894,G14895,G14896,G14897,G14898,G14899,G14900,
       G14901,G14902,G14903,G14904,G14905,G14906,G14907,G14908,G14909,G14910,G14911,G14912,G14913,G14914,G14915,G14916,G14917,G14918,G14919,G14920,
       G14921,G14922,G14923,G14924,G14925,G14926,G14927,G14928,G14929,G14930,G14931,G14932,G14933,G14934,G14935,G14936,G14937,G14938,G14939,G14940,
       G14941,G14942,G14943,G14944,G14945,G14946,G14947,G14948,G14949,G14950,G14951,G14952,G14953,G14954,G14955,G14956,G14957,G14958,G14959,G14960,
       G14961,G14962,G14963,G14964,G14965,G14966,G14967,G14968,G14969,G14970,G14971,G14972,G14973,G14974,G14975,G14976,G14977,G14978,G14979,G14980,
       G14981,G14982,G14983,G14984,G14985,G14986,G14987,G14988,G14989,G14990,G14991,G14992,G14993,G14994,G14995,G14996,G14997,G14998,G14999,G15000,
       G15001,G15002,G15003,G15004,G15005,G15006,G15007,G15008,G15009,G15010,G15011,G15012,G15013,G15014,G15015,G15016,G15017,G15018,G15019,G15020,
       G15021,G15022,G15023,G15024,G15025,G15026,G15027,G15028,G15029,G15030,G15031,G15032,G15033,G15034,G15035,G15036,G15037,G15038,G15039,G15040,
       G15041,G15042,G15043,G15044,G15045,G15046,G15047,G15048,G15049,G15050,G15051,G15052,G15053,G15054,G15055,G15056,G15057,G15058,G15059,G15060,
       G15061,G15062,G15063,G15064,G15065,G15066,G15067,G15068,G15069,G15070,G15071,G15072,G15073,G15074,G15075,G15076,G15077,G15078,G15079,G15080,
       G15081,G15082,G15083,G15084,G15085,G15086,G15087,G15088,G15089,G15090,G15091,G15092,G15093,G15094,G15095,G15096,G15097,G15098,G15099,G15100,
       G15101,G15102,G15103,G15104,G15105,G15106,G15107,G15108,G15109,G15110,G15111,G15112,G15113,G15114,G15115,G15116,G15117,G15118,G15119,G15120,
       G15121,G15122,G15123,G15124,G15125,G15126,G15127,G15128,G15129,G15130,G15131,G15132,G15133,G15134,G15135,G15136,G15137,G15138,G15139,G15140,
       G15141,G15142,G15143,G15144,G15145,G15146,G15147,G15148,G15149,G15150,G15151,G15152,G15153,G15154,G15155,G15156,G15157,G15158,G15159,G15160,
       G15161,G15162,G15163,G15164,G15165,G15166,G15167,G15168,G15169,G15170,G15171,G15172,G15173,G15174,G15175,G15176,G15177,G15178,G15179,G15180,
       G15181,G15182,G15183,G15184,G15185,G15186,G15187,G15188,G15189,G15190,G15191,G15192,G15193,G15194,G15195,G15196,G15197,G15198,G15199,G15200,
       G15201,G15202,G15203,G15204,G15205,G15206,G15207,G15208,G15209,G15210,G15211,G15212,G15213,G15214,G15215,G15216,G15217,G15218,G15219,G15220,
       G15221,G15222,G15223,G15224,G15225,G15226,G15227,G15228,G15229,G15230,G15231,G15232,G15233,G15234,G15235,G15236,G15237,G15238,G15239,G15240,
       G15241,G15242,G15243,G15244,G15245,G15246,G15247,G15248,G15249,G15250,G15251,G15252,G15253,G15254,G15255,G15256,G15257,G15258,G15259,G15260,
       G15261,G15262,G15263,G15264,G15265,G15266,G15267,G15268,G15269,G15270,G15271,G15272,G15273,G15274,G15275,G15276,G15277,G15278,G15279,G15280,
       G15281,G15282,G15283,G15284,G15285,G15286,G15287,G15288,G15289,G15290,G15291,G15292,G15293,G15294,G15295,G15296,G15297,G15298,G15299,G15300,
       G15301,G15302,G15303,G15304,G15305,G15306,G15307,G15308,G15309,G15310,G15311,G15312,G15313,G15314,G15315,G15316,G15317,G15318,G15319,G15320,
       G15321,G15322,G15323,G15324,G15325,G15326,G15327,G15328,G15329,G15330,G15331,G15332,G15333,G15334,G15335,G15336,G15337,G15338,G15339,G15340,
       G15341,G15342,G15343,G15344,G15345,G15346,G15347,G15348,G15349,G15350,G15351,G15352,G15353,G15354,G15355,G15356,G15357,G15358,G15359,G15360,
       G15361,G15362,G15363,G15364,G15365,G15366,G15367,G15368,G15369,G15370,G15371,G15372,G15373,G15374,G15375,G15376,G15377,G15378,G15379,G15380,
       G15381,G15382,G15383,G15384,G15385,G15386,G15387,G15388,G15389,G15390,G15391,G15392,G15393,G15394,G15395,G15396,G15397,G15398,G15399,G15400,
       G15401,G15402,G15403,G15404,G15405,G15406,G15407,G15408,G15409,G15410,G15411,G15412,G15413,G15414,G15415,G15416,G15417,G15418,G15419,G15420,
       G15421,G15422,G15423,G15424,G15425,G15426,G15427,G15428,G15429,G15430,G15431,G15432,G15433,G15434,G15435,G15436,G15437,G15438,G15439,G15440,
       G15441,G15442,G15443,G15444,G15445,G15446,G15447,G15448,G15449,G15450,G15451,G15452,G15453,G15454,G15455,G15456,G15457,G15458,G15459,G15460,
       G15461,G15462,G15463,G15464,G15465,G15466,G15467,G15468,G15469,G15470,G15471,G15472,G15473,G15474,G15475,G15476,G15477,G15478,G15479,G15480,
       G15481,G15482,G15483,G15484,G15485,G15486,G15487,G15488,G15489,G15490,G15491,G15492,G15493,G15494,G15495,G15496,G15497,G15498,G15499,G15500,
       G15501,G15502,G15503,G15504,G15505,G15506,G15507,G15508,G15509,G15510,G15511,G15512,G15513,G15514,G15515,G15516,G15517,G15518,G15519,G15520,
       G15521,G15522,G15523,G15524,G15525,G15526,G15527,G15528,G15529,G15530,G15531,G15532,G15533,G15534,G15535,G15536,G15537,G15538,G15539,G15540,
       G15541,G15542,G15543,G15544,G15545,G15546,G15547,G15548,G15549,G15550,G15551,G15552,G15553,G15554,G15555,G15556,G15557,G15558,G15559,G15560,
       G15561,G15562,G15563,G15564,G15565,G15566,G15567,G15568,G15569,G15570,G15571,G15572,G15573,G15574,G15575,G15576,G15577,G15578,G15579,G15580,
       G15581,G15582,G15583,G15584,G15585,G15586,G15587,G15588,G15589,G15590,G15591,G15592,G15593,G15594,G15595,G15596,G15597,G15598,G15599,G15600,
       G15601,G15602,G15603,G15604,G15605,G15606,G15607,G15608,G15609,G15610,G15611,G15612,G15613,G15614,G15615,G15616,G15617,G15618,G15619,G15620,
       G15621,G15622,G15623,G15624,G15625,G15626,G15627,G15628,G15629,G15630,G15631,G15632,G15633,G15634,G15635,G15636,G15637,G15638,G15639,G15640,
       G15641,G15642,G15643,G15644,G15645,G15646,G15647,G15648,G15649,G15650,G15651,G15652,G15653,G15654,G15655,G15656,G15657,G15658,G15659,G15660,
       G15661,G15662,G15663,G15664,G15665,G15666,G15667,G15668,G15669,G15670,G15671,G15672,G15673,G15674,G15675,G15676,G15677,G15678,G15679,G15680,
       G15681,G15682,G15683,G15684,G15685,G15686,G15687,G15688,G15689,G15690,G15691,G15692,G15693,G15694,G15695,G15696,G15697,G15698,G15699,G15700,
       G15701,G15702,G15703,G15704,G15705,G15706,G15707,G15708,G15709,G15710,G15711,G15712,G15713,G15714,G15715,G15716,G15717,G15718,G15719,G15720,
       G15721,G15722,G15723,G15724,G15725,G15726,G15727,G15728,G15729,G15730,G15731,G15732,G15733,G15734,G15735,G15736,G15737,G15738,G15739,G15740,
       G15741,G15742,G15743,G15744,G15745,G15746,G15747,G15748,G15749,G15750,G15751,G15752,G15753,G15754,G15755,G15756,G15757,G15758,G15759,G15760,
       G15761,G15762,G15763,G15764,G15765,G15766,G15767,G15768,G15769,G15770,G15771,G15772,G15773,G15774,G15775,G15776,G15777,G15778,G15779,G15780,
       G15781,G15782,G15783,G15784,G15785,G15786,G15787,G15788,G15789,G15790,G15791,G15792,G15793,G15794,G15795,G15796,G15797,G15798,G15799,G15800,
       G15801,G15802,G15803,G15804,G15805,G15806,G15807,G15808,G15809,G15810,G15811,G15812,G15813,G15814,G15815,G15816,G15817,G15818,G15819,G15820,
       G15821,G15822,G15823,G15824,G15825,G15826,G15827,G15828,G15829,G15830,G15831,G15832,G15833,G15834,G15835,G15836,G15837,G15838,G15839,G15840,
       G15841,G15842,G15843,G15844,G15845,G15846,G15847,G15848,G15849,G15850,G15851,G15852,G15853,G15854,G15855,G15856,G15857,G15858,G15859,G15860,
       G15861,G15862,G15863,G15864,G15865,G15866,G15867,G15868,G15869,G15870,G15871,G15872,G15873,G15874,G15875,G15876,G15877,G15878,G15879,G15880,
       G15881,G15882,G15883,G15884,G15885,G15886,G15887,G15888,G15889,G15890,G15891,G15892,G15893,G15894,G15895,G15896,G15897,G15898,G15899,G15900,
       G15901,G15902,G15903,G15904,G15905,G15906,G15907,G15908,G15909,G15910,G15911,G15912,G15913,G15914,G15915,G15916,G15917,G15918,G15919,G15920,
       G15921,G15922,G15923,G15924,G15925,G15926,G15927,G15928,G15929,G15930,G15931,G15932,G15933,G15934,G15935,G15936,G15937,G15938,G15939,G15940,
       G15941,G15942,G15943,G15944,G15945,G15946,G15947,G15948,G15949,G15950,G15951,G15952,G15953,G15954,G15955,G15956,G15957,G15958,G15959,G15960,
       G15961,G15962,G15963,G15964,G15965,G15966,G15967,G15968,G15969,G15970,G15971,G15972,G15973,G15974,G15975,G15976,G15977,G15978,G15979,G15980,
       G15981,G15982,G15983,G15984,G15985,G15986,G15987,G15988,G15989,G15990,G15991,G15992,G15993,G15994,G15995,G15996,G15997,G15998,G15999,G16000,
       G16001,G16002,G16003,G16004,G16005,G16006,G16007,G16008,G16009,G16010,G16011,G16012,G16013,G16014,G16015,G16016,G16017,G16018,G16019,G16020,
       G16021,G16022,G16023,G16024,G16025,G16026,G16027,G16028,G16029,G16030,G16031,G16032,G16033,G16034,G16035,G16036,G16037,G16038,G16039,G16040,
       G16041,G16042,G16043,G16044,G16045,G16046,G16047,G16048,G16049,G16050,G16051,G16052,G16053,G16054,G16055,G16056,G16057,G16058,G16059,G16060,
       G16061,G16062,G16063,G16064,G16065,G16066,G16067,G16068,G16069,G16070,G16071,G16072,G16073,G16074,G16075,G16076,G16077,G16078,G16079,G16080,
       G16081,G16082,G16083,G16084,G16085,G16086,G16087,G16088,G16089,G16090,G16091,G16092,G16093,G16094,G16095,G16096,G16097,G16098,G16099,G16100,
       G16101,G16102,G16103,G16104,G16105,G16106,G16107,G16108,G16109,G16110,G16111,G16112,G16113,G16114,G16115,G16116,G16117,G16118,G16119,G16120,
       G16121,G16122,G16123,G16124,G16125,G16126,G16127,G16128,G16129,G16130,G16131,G16132,G16133,G16134,G16135,G16136,G16137,G16138,G16139,G16140,
       G16141,G16142,G16143,G16144,G16145,G16146,G16147,G16148,G16149,G16150,G16151,G16152,G16153,G16154,G16155,G16156,G16157,G16158,G16159,G16160,
       G16161,G16162,G16163,G16164,G16165,G16166,G16167,G16168,G16169,G16170,G16171,G16172,G16173,G16174,G16175,G16176,G16177,G16178,G16179,G16180,
       G16181,G16182,G16183,G16184,G16185,G16186,G16187,G16188,G16189,G16190,G16191,G16192,G16193,G16194,G16195,G16196,G16197,G16198,G16199,G16200,
       G16201,G16202,G16203,G16204,G16205,G16206,G16207,G16208,G16209,G16210,G16211,G16212,G16213,G16214,G16215,G16216,G16217,G16218,G16219,G16220,
       G16221,G16222,G16223,G16224,G16225,G16226,G16227,G16228,G16229,G16230,G16231,G16232,G16233,G16234,G16235,G16236,G16237,G16238,G16239,G16240,
       G16241,G16242,G16243,G16244,G16245,G16246,G16247,G16248,G16249,G16250,G16251,G16252,G16253,G16254,G16255,G16256,G16257,G16258,G16259,G16260,
       G16261,G16262,G16263,G16264,G16265,G16266,G16267,G16268,G16269,G16270,G16271,G16272,G16273,G16274,G16275,G16276,G16277,G16278,G16279,G16280,
       G16281,G16282,G16283,G16284,G16285,G16286,G16287,G16288,G16289,G16290,G16291,G16292,G16293,G16294,G16295,G16296,G16297,G16298,G16299,G16300,
       G16301,G16302,G16303,G16304,G16305,G16306,G16307,G16308,G16309,G16310,G16311,G16312,G16313,G16314,G16315,G16316,G16317,G16318,G16319,G16320,
       G16321,G16322,G16323,G16324,G16325,G16326,G16327,G16328,G16329,G16330,G16331,G16332,G16333,G16334,G16335,G16336,G16337,G16338,G16339,G16340,
       G16341,G16342,G16343,G16344,G16345,G16346,G16347,G16348,G16349,G16350,G16351,G16352,G16353,G16354,G16355,G16356,G16357,G16358,G16359,G16360,
       G16361,G16362,G16363,G16364,G16365,G16366,G16367,G16368,G16369,G16370,G16371,G16372,G16373,G16374,G16375,G16376,G16377,G16378,G16379,G16380,
       G16381,G16382,G16383,G16384,G16385,G16386,G16387,G16388,G16389,G16390,G16391,G16392,G16393,G16394,G16395,G16396,G16397,G16398,G16399,G16400,
       G16401,G16402,G16403,G16404,G16405,G16406,G16407,G16408,G16409,G16410,G16411,G16412,G16413,G16414,G16415,G16416,G16417,G16418,G16419,G16420,
       G16421,G16422,G16423,G16424,G16425,G16426,G16427,G16428,G16429,G16430,G16431,G16432,G16433,G16434,G16435,G16436,G16437,G16438,G16439,G16440,
       G16441,G16442,G16443,G16444,G16445,G16446,G16447,G16448,G16449,G16450,G16451,G16452,G16453,G16454,G16455,G16456,G16457,G16458,G16459,G16460,
       G16461,G16462,G16463,G16464,G16465,G16466,G16467,G16468,G16469,G16470,G16471,G16472,G16473,G16474,G16475,G16476,G16477,G16478,G16479,G16480,
       G16481,G16482,G16483,G16484,G16485,G16486,G16487,G16488,G16489,G16490,G16491,G16492,G16493,G16494,G16495,G16496,G16497,G16498,G16499,G16500,
       G16501,G16502,G16503,G16504,G16505,G16506,G16507,G16508,G16509,G16510,G16511,G16512,G16513,G16514,G16515,G16516,G16517,G16518,G16519,G16520,
       G16521,G16522,G16523,G16524,G16525,G16526,G16527,G16528,G16529,G16530,G16531,G16532,G16533,G16534,G16535,G16536,G16537,G16538,G16539,G16540,
       G16541,G16542,G16543,G16544,G16545,G16546,G16547,G16548,G16549,G16550,G16551,G16552,G16553,G16554,G16555,G16556,G16557,G16558,G16559,G16560,
       G16561,G16562,G16563,G16564,G16565,G16566,G16567,G16568,G16569,G16570,G16571,G16572,G16573,G16574,G16575,G16576,G16577,G16578,G16579,G16580,
       G16581,G16582,G16583,G16584,G16585,G16586,G16587,G16588,G16589,G16590,G16591,G16592,G16593,G16594,G16595,G16596,G16597,G16598,G16599,G16600,
       G16601,G16602,G16603,G16604,G16605,G16606,G16607,G16608,G16609,G16610,G16611,G16612,G16613,G16614,G16615,G16616,G16617,G16618,G16619,G16620,
       G16621,G16622,G16623,G16624,G16625,G16626,G16627,G16628,G16629,G16630,G16631,G16632,G16633,G16634,G16635,G16636,G16637,G16638,G16639,G16640,
       G16641,G16642,G16643,G16644,G16645,G16646,G16647,G16648,G16649,G16650,G16651,G16652,G16653,G16654,G16655,G16656,G16657,G16658,G16659,G16660,
       G16661,G16662,G16663,G16664,G16665,G16666,G16667,G16668,G16669,G16670,G16671,G16672,G16673,G16674,G16675,G16676,G16677,G16678,G16679,G16680,
       G16681,G16682,G16683,G16684,G16685,G16686,G16687,G16688,G16689,G16690,G16691,G16692,G16693,G16694,G16695,G16696,G16697,G16698,G16699,G16700,
       G16701,G16702,G16703,G16704,G16705,G16706,G16707,G16708,G16709,G16710,G16711,G16712,G16713,G16714,G16715,G16716,G16717,G16718,G16719,G16720,
       G16721,G16722,G16723,G16724,G16725,G16726,G16727,G16728,G16729,G16730,G16731,G16732,G16733,G16734,G16735,G16736,G16737,G16738,G16739,G16740,
       G16741,G16742,G16743,G16744,G16745,G16746,G16747,G16748,G16749,G16750,G16751,G16752,G16753,G16754,G16755,G16756,G16757,G16758,G16759,G16760,
       G16761,G16762,G16763,G16764,G16765,G16766,G16767,G16768,G16769,G16770,G16771,G16772,G16773,G16774,G16775,G16776,G16777,G16778,G16779,G16780,
       G16781,G16782,G16783,G16784,G16785,G16786,G16787,G16788,G16789,G16790,G16791,G16792,G16793,G16794,G16795,G16796,G16797,G16798,G16799,G16800,
       G16801,G16802,G16803,G16804,G16805,G16806,G16807,G16808,G16809,G16810,G16811,G16812,G16813,G16814,G16815,G16816,G16817,G16818,G16819,G16820,
       G16821,G16822,G16823,G16824,G16825,G16826,G16827,G16828,G16829,G16830,G16831,G16832,G16833,G16834,G16835,G16836,G16837,G16838,G16839,G16840,
       G16841,G16842,G16843,G16844,G16845,G16846,G16847,G16848,G16849,G16850,G16851,G16852,G16853,G16854,G16855,G16856,G16857,G16858,G16859,G16860,
       G16861,G16862,G16863,G16864,G16865,G16866,G16867,G16868,G16869,G16870,G16871,G16872,G16873,G16874,G16875,G16876,G16877,G16878,G16879,G16880,
       G16881,G16882,G16883,G16884,G16885,G16886,G16887,G16888,G16889,G16890,G16891,G16892,G16893,G16894,G16895,G16896,G16897,G16898,G16899,G16900,
       G16901,G16902,G16903,G16904,G16905,G16906,G16907,G16908,G16909,G16910,G16911,G16912,G16913,G16914,G16915,G16916,G16917,G16918,G16919,G16920,
       G16921,G16922,G16923,G16924,G16925,G16926,G16927,G16928,G16929,G16930,G16931,G16932,G16933,G16934,G16935,G16936,G16937,G16938,G16939,G16940,
       G16941,G16942,G16943,G16944,G16945,G16946,G16947,G16948,G16949,G16950,G16951,G16952,G16953,G16954,G16955,G16956,G16957,G16958,G16959,G16960,
       G16961,G16962,G16963,G16964,G16965,G16966,G16967,G16968,G16969,G16970,G16971,G16972,G16973,G16974,G16975,G16976,G16977,G16978,G16979,G16980,
       G16981,G16982,G16983,G16984,G16985,G16986,G16987,G16988,G16989,G16990,G16991,G16992,G16993,G16994,G16995,G16996,G16997,G16998,G16999,G17000,
       G17001,G17002,G17003,G17004,G17005,G17006,G17007,G17008,G17009,G17010,G17011,G17012,G17013,G17014,G17015,G17016,G17017,G17018,G17019,G17020,
       G17021,G17022,G17023,G17024,G17025,G17026,G17027,G17028,G17029,G17030,G17031,G17032,G17033,G17034,G17035,G17036,G17037,G17038,G17039,G17040,
       G17041,G17042,G17043,G17044,G17045,G17046,G17047,G17048,G17049,G17050,G17051,G17052,G17053,G17054,G17055,G17056,G17057,G17058,G17059,G17060,
       G17061,G17062,G17063,G17064,G17065,G17066,G17067,G17068,G17069,G17070,G17071,G17072,G17073,G17074,G17075,G17076,G17077,G17078,G17079,G17080,
       G17081,G17082,G17083,G17084,G17085,G17086,G17087,G17088,G17089,G17090,G17091,G17092,G17093,G17094,G17095,G17096,G17097,G17098,G17099,G17100,
       G17101,G17102,G17103,G17104,G17105,G17106,G17107,G17108,G17109,G17110,G17111,G17112,G17113,G17114,G17115,G17116,G17117,G17118,G17119,G17120,
       G17121,G17122,G17123,G17124,G17125,G17126,G17127,G17128,G17129,G17130,G17131,G17132,G17133,G17134,G17135,G17136,G17137,G17138,G17139,G17140,
       G17141,G17142,G17143,G17144,G17145,G17146,G17147,G17148,G17149,G17150,G17151,G17152,G17153,G17154,G17155,G17156,G17157,G17158,G17159,G17160,
       G17161,G17162,G17163,G17164,G17165,G17166,G17167,G17168,G17169,G17170,G17171,G17172,G17173,G17174,G17175,G17176,G17177,G17178,G17179,G17180,
       G17181,G17182,G17183,G17184,G17185,G17186,G17187,G17188,G17189,G17190,G17191,G17192,G17193,G17194,G17195,G17196,G17197,G17198,G17199,G17200,
       G17201,G17202,G17203,G17204,G17205,G17206,G17207,G17208,G17209,G17210,G17211,G17212,G17213,G17214,G17215,G17216,G17217,G17218,G17219,G17220,
       G17221,G17222,G17223,G17224,G17225,G17226,G17227,G17228,G17229,G17230,G17231,G17232,G17233,G17234,G17235,G17236,G17237,G17238,G17239,G17240,
       G17241,G17242,G17243,G17244,G17245,G17246,G17247,G17248,G17249,G17250,G17251,G17252,G17253,G17254,G17255,G17256,G17257,G17258,G17259,G17260,
       G17261,G17262,G17263,G17264,G17265,G17266,G17267,G17268,G17269,G17270,G17271,G17272,G17273,G17274,G17275,G17276,G17277,G17278,G17279,G17280,
       G17281,G17282,G17283,G17284,G17285,G17286,G17287,G17288,G17289,G17290,G17291,G17292,G17293,G17294,G17295,G17296,G17297,G17298,G17299,G17300,
       G17301,G17302,G17303,G17304,G17305,G17306,G17307,G17308,G17309,G17310,G17311,G17312,G17313,G17314,G17315,G17316,G17317,G17318,G17319,G17320,
       G17321,G17322,G17323,G17324,G17325,G17326,G17327,G17328,G17329,G17330,G17331,G17332,G17333,G17334,G17335,G17336,G17337,G17338,G17339,G17340,
       G17341,G17342,G17343,G17344,G17345,G17346,G17347,G17348,G17349,G17350,G17351,G17352,G17353,G17354,G17355,G17356,G17357,G17358,G17359,G17360,
       G17361,G17362,G17363,G17364,G17365,G17366,G17367,G17368,G17369,G17370,G17371,G17372,G17373,G17374,G17375,G17376,G17377,G17378,G17379,G17380,
       G17381,G17382,G17383,G17384,G17385,G17386,G17387,G17388,G17389,G17390,G17391,G17392,G17393,G17394,G17395,G17396,G17397,G17398,G17399,G17400,
       G17401,G17402,G17403,G17404,G17405,G17406,G17407,G17408,G17409,G17410,G17411,G17412,G17413,G17414,G17415,G17416,G17417,G17418,G17419,G17420,
       G17421,G17422,G17423,G17424,G17425,G17426,G17427,G17428,G17429,G17430,G17431,G17432,G17433,G17434,G17435,G17436,G17437,G17438,G17439,G17440,
       G17441,G17442,G17443,G17444,G17445,G17446,G17447,G17448,G17449,G17450,G17451,G17452,G17453,G17454,G17455,G17456,G17457,G17458,G17459,G17460,
       G17461,G17462,G17463,G17464,G17465,G17466,G17467,G17468,G17469,G17470,G17471,G17472,G17473,G17474,G17475,G17476,G17477,G17478,G17479,G17480,
       G17481,G17482,G17483,G17484,G17485,G17486,G17487,G17488,G17489,G17490,G17491,G17492,G17493,G17494,G17495,G17496,G17497,G17498,G17499,G17500,
       G17501,G17502,G17503,G17504,G17505,G17506,G17507,G17508,G17509,G17510,G17511,G17512,G17513,G17514,G17515,G17516,G17517,G17518,G17519,G17520,
       G17521,G17522,G17523,G17524,G17525,G17526,G17527,G17528,G17529,G17530,G17531,G17532,G17533,G17534,G17535,G17536,G17537,G17538,G17539,G17540,
       G17541,G17542,G17543,G17544,G17545,G17546,G17547,G17548,G17549,G17550,G17551,G17552,G17553,G17554,G17555,G17556,G17557,G17558,G17559,G17560,
       G17561,G17562,G17563,G17564,G17565,G17566,G17567,G17568,G17569,G17570,G17571,G17572,G17573,G17574,G17575,G17576,G17577,G17578,G17579,G17580,
       G17581,G17582,G17583,G17584,G17585,G17586,G17587,G17588,G17589,G17590,G17591,G17592,G17593,G17594,G17595,G17596,G17597,G17598,G17599,G17600,
       G17601,G17602,G17603,G17604,G17605,G17606,G17607,G17608,G17609,G17610,G17611,G17612,G17613,G17614,G17615,G17616,G17617,G17618,G17619,G17620,
       G17621,G17622,G17623,G17624,G17625,G17626,G17627,G17628,G17629,G17630,G17631,G17632,G17633,G17634,G17635,G17636,G17637,G17638,G17639,G17640,
       G17641,G17642,G17643,G17644,G17645,G17646,G17647,G17648,G17649,G17650,G17651,G17652,G17653,G17654,G17655,G17656,G17657,G17658,G17659,G17660,
       G17661,G17662,G17663,G17664,G17665,G17666,G17667,G17668,G17669,G17670,G17671,G17672,G17673,G17674,G17675,G17676,G17677,G17678,G17679,G17680,
       G17681,G17682,G17683,G17684,G17685,G17686,G17687,G17688,G17689,G17690,G17691,G17692,G17693,G17694,G17695,G17696,G17697,G17698,G17699,G17700,
       G17701,G17702,G17703,G17704,G17705,G17706,G17707,G17708,G17709,G17710,G17711,G17712,G17713,G17714,G17715,G17716,G17717,G17718,G17719,G17720,
       G17721,G17722,G17723,G17724,G17725,G17726,G17727,G17728,G17729,G17730,G17731,G17732,G17733,G17734,G17735,G17736,G17737,G17738,G17739,G17740,
       G17741,G17742,G17743,G17744,G17745,G17746,G17747,G17748,G17749,G17750,G17751,G17752,G17753,G17754,G17755,G17756,G17757,G17758,G17759,G17760,
       G17761,G17762,G17763,G17764,G17765,G17766,G17767,G17768,G17769,G17770,G17771,G17772,G17773,G17774,G17775,G17776,G17777,G17778,G17779,G17780,
       G17781,G17782,G17783,G17784,G17785,G17786,G17787,G17788,G17789,G17790,G17791,G17792,G17793,G17794,G17795,G17796,G17797,G17798,G17799,G17800,
       G17801,G17802,G17803,G17804,G17805,G17806,G17807,G17808,G17809,G17810,G17811,G17812,G17813,G17814,G17815,G17816,G17817,G17818,G17819,G17820,
       G17821,G17822,G17823,G17824,G17825,G17826,G17827,G17828,G17829,G17830,G17831,G17832,G17833,G17834,G17835,G17836,G17837,G17838,G17839,G17840,
       G17841,G17842,G17843,G17844,G17845,G17846,G17847,G17848,G17849,G17850,G17851,G17852,G17853,G17854,G17855,G17856,G17857,G17858,G17859,G17860,
       G17861,G17862,G17863,G17864,G17865,G17866,G17867,G17868,G17869,G17870,G17871,G17872,G17873,G17874,G17875,G17876,G17877,G17878,G17879,G17880,
       G17881,G17882,G17883,G17884,G17885,G17886,G17887,G17888,G17889,G17890,G17891,G17892,G17893,G17894,G17895,G17896,G17897,G17898,G17899,G17900,
       G17901,G17902,G17903,G17904,G17905,G17906,G17907,G17908,G17909,G17910,G17911,G17912,G17913,G17914,G17915,G17916,G17917,G17918,G17919,G17920,
       G17921,G17922,G17923,G17924,G17925,G17926,G17927,G17928,G17929,G17930,G17931,G17932,G17933,G17934,G17935,G17936,G17937,G17938,G17939,G17940,
       G17941,G17942,G17943,G17944,G17945,G17946,G17947,G17948,G17949,G17950,G17951,G17952,G17953,G17954,G17955,G17956,G17957,G17958,G17959,G17960,
       G17961,G17962,G17963,G17964,G17965,G17966,G17967,G17968,G17969,G17970,G17971,G17972,G17973,G17974,G17975,G17976,G17977,G17978,G17979,G17980,
       G17981,G17982,G17983,G17984,G17985,G17986,G17987,G17988,G17989,G17990,G17991,G17992,G17993,G17994,G17995,G17996,G17997,G17998,G17999,G18000,
       G18001,G18002,G18003,G18004,G18005,G18006,G18007,G18008,G18009,G18010,G18011,G18012,G18013,G18014,G18015,G18016,G18017,G18018,G18019,G18020,
       G18021,G18022,G18023,G18024,G18025,G18026,G18027,G18028,G18029,G18030,G18031,G18032,G18033,G18034,G18035,G18036,G18037,G18038,G18039,G18040,
       G18041,G18042,G18043,G18044,G18045,G18046,G18047,G18048,G18049,G18050,G18051,G18052,G18053,G18054,G18055,G18056,G18057,G18058,G18059,G18060,
       G18061,G18062,G18063,G18064,G18065,G18066,G18067,G18068,G18069,G18070,G18071,G18072,G18073,G18074,G18075,G18076,G18077,G18078,G18079,G18080,
       G18081,G18082,G18083,G18084,G18085,G18086,G18087,G18088,G18089,G18090,G18091,G18092,G18093,G18094,G18095,G18096,G18097,G18098,G18099,G18100,
       G18101,G18102,G18103,G18104,G18105,G18106,G18107,G18108,G18109,G18110,G18111,G18112,G18113,G18114,G18115,G18116,G18117,G18118,G18119,G18120,
       G18121,G18122,G18123,G18124,G18125,G18126,G18127,G18128,G18129,G18130,G18131,G18132,G18133,G18134,G18135,G18136,G18137,G18138,G18139,G18140,
       G18141,G18142,G18143,G18144,G18145,G18146,G18147,G18148,G18149,G18150,G18151,G18152,G18153,G18154,G18155,G18156,G18157,G18158,G18159,G18160,
       G18161,G18162,G18163,G18164,G18165,G18166,G18167,G18168,G18169,G18170,G18171,G18172,G18173,G18174,G18175,G18176,G18177,G18178,G18179,G18180,
       G18181,G18182,G18183,G18184,G18185,G18186,G18187,G18188,G18189,G18190,G18191,G18192,G18193,G18194,G18195,G18196,G18197,G18198,G18199,G18200,
       G18201,G18202,G18203,G18204,G18205,G18206,G18207,G18208,G18209,G18210,G18211,G18212,G18213,G18214,G18215,G18216,G18217,G18218,G18219,G18220,
       G18221,G18222,G18223,G18224,G18225,G18226,G18227,G18228,G18229,G18230,G18231,G18232,G18233,G18234,G18235,G18236,G18237,G18238,G18239,G18240,
       G18241,G18242,G18243,G18244,G18245,G18246,G18247,G18248,G18249,G18250,G18251,G18252,G18253,G18254,G18255,G18256,G18257,G18258,G18259,G18260,
       G18261,G18262,G18263,G18264,G18265,G18266,G18267,G18268,G18269,G18270,G18271,G18272,G18273,G18274,G18275,G18276,G18277,G18278,G18279,G18280,
       G18281,G18282,G18283,G18284,G18285,G18286,G18287,G18288,G18289,G18290,G18291,G18292,G18293,G18294,G18295,G18296,G18297,G18298,G18299,G18300,
       G18301,G18302,G18303,G18304,G18305,G18306,G18307,G18308,G18309,G18310,G18311,G18312,G18313,G18314,G18315,G18316,G18317,G18318,G18319,G18320,
       G18321,G18322,G18323,G18324,G18325,G18326,G18327,G18328,G18329,G18330,G18331,G18332,G18333,G18334,G18335,G18336,G18337,G18338,G18339,G18340,
       G18341,G18342,G18343,G18344,G18345,G18346,G18347,G18348,G18349,G18350,G18351,G18352,G18353,G18354,G18355,G18356,G18357,G18358,G18359,G18360,
       G18361,G18362,G18363,G18364,G18365,G18366,G18367,G18368,G18369,G18370,G18371,G18372,G18373,G18374,G18375,G18376,G18377,G18378,G18379,G18380,
       G18381,G18382,G18383,G18384,G18385,G18386,G18387,G18388,G18389,G18390,G18391,G18392,G18393,G18394,G18395,G18396,G18397,G18398,G18399,G18400,
       G18401,G18402,G18403,G18404,G18405,G18406,G18407,G18408,G18409,G18410,G18411,G18412,G18413,G18414,G18415,G18416,G18417,G18418,G18419,G18420,
       G18421,G18422,G18423,G18424,G18425,G18426,G18427,G18428,G18429,G18430,G18431,G18432,G18433,G18434,G18435,G18436,G18437,G18438,G18439,G18440,
       G18441,G18442,G18443,G18444,G18445,G18446,G18447,G18448,G18449,G18450,G18451,G18452,G18453,G18454,G18455,G18456,G18457,G18458,G18459,G18460,
       G18461,G18462,G18463,G18464,G18465,G18466,G18467,G18468,G18469,G18470,G18471,G18472,G18473,G18474,G18475,G18476,G18477,G18478,G18479,G18480,
       G18481,G18482,G18483,G18484,G18485,G18486,G18487,G18488,G18489,G18490,G18491,G18492,G18493,G18494,G18495,G18496,G18497,G18498,G18499,G18500,
       G18501,G18502,G18503,G18504,G18505,G18506,G18507,G18508,G18509,G18510,G18511,G18512,G18513,G18514,G18515,G18516,G18517,G18518,G18519,G18520,
       G18521,G18522,G18523,G18524,G18525,G18526,G18527,G18528,G18529,G18530,G18531,G18532,G18533,G18534,G18535,G18536,G18537,G18538,G18539,G18540,
       G18541,G18542,G18543,G18544,G18545,G18546,G18547,G18548,G18549,G18550,G18551,G18552,G18553,G18554,G18555,G18556,G18557,G18558,G18559,G18560,
       G18561,G18562,G18563,G18564,G18565,G18566,G18567,G18568,G18569,G18570,G18571,G18572,G18573,G18574,G18575,G18576,G18577,G18578,G18579,G18580,
       G18581,G18582,G18583,G18584,G18585,G18586,G18587,G18588,G18589,G18590,G18591,G18592,G18593,G18594,G18595,G18596,G18597,G18598,G18599,G18600,
       G18601,G18602,G18603,G18604,G18605,G18606,G18607,G18608,G18609,G18610,G18611,G18612,G18613,G18614,G18615,G18616,G18617,G18618,G18619,G18620,
       G18621,G18622,G18623,G18624,G18625,G18626,G18627,G18628,G18629,G18630,G18631,G18632,G18633,G18634,G18635,G18636,G18637,G18638,G18639,G18640,
       G18641,G18642,G18643,G18644,G18645,G18646,G18647,G18648,G18649,G18650,G18651,G18652,G18653,G18654,G18655,G18656,G18657,G18658,G18659,G18660,
       G18661,G18662,G18663,G18664,G18665,G18666,G18667,G18668,G18669,G18670,G18671,G18672,G18673,G18674,G18675,G18676,G18677,G18678,G18679,G18680,
       G18681,G18682,G18683,G18684,G18685,G18686,G18687,G18688,G18689,G18690,G18691,G18692,G18693,G18694,G18695,G18696,G18697,G18698,G18699,G18700,
       G18701,G18702,G18703,G18704,G18705,G18706,G18707,G18708,G18709,G18710,G18711,G18712,G18713,G18714,G18715,G18716,G18717,G18718,G18719,G18720,
       G18721,G18722,G18723,G18724,G18725,G18726,G18727,G18728,G18729,G18730,G18731,G18732,G18733,G18734,G18735,G18736,G18737,G18738,G18739,G18740,
       G18741,G18742,G18743,G18744,G18745,G18746,G18747,G18748,G18749,G18750,G18751,G18752,G18753,G18754,G18755,G18756,G18757,G18758,G18759,G18760,
       G18761,G18762,G18763,G18764,G18765,G18766,G18767,G18768,G18769,G18770,G18771,G18772,G18773,G18774,G18775,G18776,G18777,G18778,G18779,G18780,
       G18781,G18782,G18783,G18784,G18785,G18786,G18787,G18788,G18789,G18790,G18791,G18792,G18793,G18794,G18795,G18796,G18797,G18798,G18799,G18800,
       G18801,G18802,G18803,G18804,G18805,G18806,G18807,G18808,G18809,G18810,G18811,G18812,G18813,G18814,G18815,G18816,G18817,G18818,G18819,G18820,
       G18821,G18822,G18823,G18824,G18825,G18826,G18827,G18828,G18829,G18830,G18831,G18832,G18833,G18834,G18835,G18836,G18837,G18838,G18839,G18840,
       G18841,G18842,G18843,G18844,G18845,G18846,G18847,G18848,G18849,G18850,G18851,G18852,G18853,G18854,G18855,G18856,G18857,G18858,G18859,G18860,
       G18861,G18862,G18863,G18864,G18865,G18866,G18867,G18868,G18869,G18870,G18871,G18872,G18873,G18874,G18875,G18876,G18877,G18878,G18879,G18880,
       G18881,G18882,G18883,G18884,G18885,G18886,G18887,G18888,G18889,G18890,G18891,G18892,G18893,G18894,G18895,G18896,G18897,G18898,G18899,G18900,
       G18901,G18902,G18903,G18904,G18905,G18906,G18907,G18908,G18909,G18910,G18911,G18912,G18913,G18914,G18915,G18916,G18917,G18918,G18919,G18920,
       G18921,G18922,G18923,G18924,G18925,G18926,G18927,G18928,G18929,G18930,G18931,G18932,G18933,G18934,G18935,G18936,G18937,G18938,G18939,G18940,
       G18941,G18942,G18943,G18944,G18945,G18946,G18947,G18948,G18949,G18950,G18951,G18952,G18953,G18954,G18955,G18956,G18957,G18958,G18959,G18960,
       G18961,G18962,G18963,G18964,G18965,G18966,G18967,G18968,G18969,G18970,G18971,G18972,G18973,G18974,G18975,G18976,G18977,G18978,G18979,G18980,
       G18981,G18982,G18983,G18984,G18985,G18986,G18987,G18988,G18989,G18990,G18991,G18992,G18993,G18994,G18995,G18996,G18997,G18998,G18999,G19000,
       G19001,G19002,G19003,G19004,G19005,G19006,G19007,G19008,G19009,G19010,G19011,G19012,G19013,G19014,G19015,G19016,G19017,G19018,G19019,G19020,
       G19021,G19022,G19023,G19024,G19025,G19026,G19027,G19028,G19029,G19030,G19031,G19032,G19033,G19034,G19035,G19036,G19037,G19038,G19039,G19040,
       G19041,G19042,G19043,G19044,G19045,G19046,G19047,G19048,G19049,G19050,G19051,G19052,G19053,G19054,G19055,G19056,G19057,G19058,G19059,G19060,
       G19061,G19062,G19063,G19064,G19065,G19066,G19067,G19068,G19069,G19070,G19071,G19072,G19073,G19074,G19075,G19076,G19077,G19078,G19079,G19080,
       G19081,G19082,G19083,G19084,G19085,G19086,G19087,G19088,G19089,G19090,G19091,G19092,G19093,G19094,G19095,G19096,G19097,G19098,G19099,G19100,
       G19101,G19102,G19103,G19104,G19105,G19106,G19107,G19108,G19109,G19110,G19111,G19112,G19113,G19114,G19115,G19116,G19117,G19118,G19119,G19120,
       G19121,G19122,G19123,G19124,G19125,G19126,G19127,G19128,G19129,G19130,G19131,G19132,G19133,G19134,G19135,G19136,G19137,G19138,G19139,G19140,
       G19141,G19142,G19143,G19144,G19145,G19146,G19147,G19148,G19149,G19150,G19151,G19152,G19153,G19154,G19155,G19156,G19157,G19158,G19159,G19160,
       G19161,G19162,G19163,G19164,G19165,G19166,G19167,G19168,G19169,G19170,G19171,G19172,G19173,G19174,G19175,G19176,G19177,G19178,G19179,G19180,
       G19181,G19182,G19183,G19184,G19185,G19186,G19187,G19188,G19189,G19190,G19191,G19192,G19193,G19194,G19195,G19196,G19197,G19198,G19199,G19200,
       G19201,G19202,G19203,G19204,G19205,G19206,G19207,G19208,G19209,G19210,G19211,G19212,G19213,G19214,G19215,G19216,G19217,G19218,G19219,G19220,
       G19221,G19222,G19223,G19224,G19225,G19226,G19227,G19228,G19229,G19230,G19231,G19232,G19233,G19234,G19235,G19236,G19237,G19238,G19239,G19240,
       G19241,G19242,G19243,G19244,G19245,G19246,G19247,G19248,G19249,G19250,G19251,G19252,G19253,G19254,G19255,G19256,G19257,G19258,G19259,G19260,
       G19261,G19262,G19263,G19264,G19265,G19266,G19267,G19268,G19269,G19270,G19271,G19272,G19273,G19274,G19275,G19276,G19277,G19278,G19279,G19280,
       G19281,G19282,G19283,G19284,G19285,G19286,G19287,G19288,G19289,G19290,G19291,G19292,G19293,G19294,G19295,G19296,G19297,G19298,G19299,G19300,
       G19301,G19302,G19303,G19304,G19305,G19306,G19307,G19308,G19309,G19310,G19311,G19312,G19313,G19314,G19315,G19316,G19317,G19318,G19319,G19320,
       G19321,G19322,G19323,G19324,G19325,G19326,G19327,G19328,G19329,G19330,G19331,G19332,G19333,G19334,G19335,G19336,G19337,G19338,G19339,G19340,
       G19341,G19342,G19343,G19344,G19345,G19346,G19347,G19348,G19349,G19350,G19351,G19352,G19353,G19354,G19355,G19356,G19357,G19358,G19359,G19360,
       G19361,G19362,G19363,G19364,G19365,G19366,G19367,G19368,G19369,G19370,G19371,G19372,G19373,G19374,G19375,G19376,G19377,G19378,G19379,G19380,
       G19381,G19382,G19383,G19384,G19385,G19386,G19387,G19388,G19389,G19390,G19391,G19392,G19393,G19394,G19395,G19396,G19397,G19398,G19399,G19400,
       G19401,G19402,G19403,G19404,G19405,G19406,G19407,G19408,G19409,G19410,G19411,G19412,G19413,G19414,G19415,G19416,G19417,G19418,G19419,G19420,
       G19421,G19422,G19423,G19424,G19425,G19426,G19427,G19428,G19429,G19430,G19431,G19432,G19433,G19434,G19435,G19436,G19437,G19438,G19439,G19440,
       G19441,G19442,G19443,G19444,G19445,G19446,G19447,G19448,G19449,G19450,G19451,G19452,G19453,G19454,G19455,G19456,G19457,G19458,G19459,G19460,
       G19461,G19462,G19463,G19464,G19465,G19466,G19467,G19468,G19469,G19470,G19471,G19472,G19473,G19474,G19475,G19476,G19477,G19478,G19479,G19480,
       G19481,G19482,G19483,G19484,G19485,G19486,G19487,G19488,G19489,G19490,G19491,G19492,G19493,G19494,G19495,G19496,G19497,G19498,G19499,G19500,
       G19501,G19502,G19503,G19504,G19505,G19506,G19507,G19508,G19509,G19510,G19511,G19512,G19513,G19514,G19515,G19516,G19517,G19518,G19519,G19520,
       G19521,G19522,G19523,G19524,G19525,G19526,G19527,G19528,G19529,G19530,G19531,G19532,G19533,G19534,G19535,G19536,G19537,G19538,G19539,G19540,
       G19541,G19542,G19543,G19544,G19545,G19546,G19547,G19548,G19549,G19550,G19551,G19552,G19553,G19554,G19555,G19556,G19557,G19558,G19559,G19560,
       G19561,G19562,G19563,G19564,G19565,G19566,G19567,G19568,G19569,G19570,G19571,G19572,G19573,G19574,G19575,G19576,G19577,G19578,G19579,G19580,
       G19581,G19582,G19583,G19584,G19585,G19586,G19587,G19588,G19589,G19590,G19591,G19592,G19593,G19594,G19595,G19596,G19597,G19598,G19599,G19600,
       G19601,G19602,G19603,G19604,G19605,G19606,G19607,G19608,G19609,G19610,G19611,G19612,G19613,G19614,G19615,G19616,G19617,G19618,G19619,G19620,
       G19621,G19622,G19623,G19624,G19625,G19626,G19627,G19628,G19629,G19630,G19631,G19632,G19633,G19634,G19635,G19636,G19637,G19638,G19639,G19640,
       G19641,G19642,G19643,G19644,G19645,G19646,G19647,G19648,G19649,G19650,G19651,G19652,G19653,G19654,G19655,G19656,G19657,G19658,G19659,G19660,
       G19661,G19662,G19663,G19664,G19665,G19666,G19667,G19668,G19669,G19670,G19671,G19672,G19673,G19674,G19675,G19676,G19677,G19678,G19679,G19680,
       G19681,G19682,G19683,G19684,G19685,G19686,G19687,G19688,G19689,G19690,G19691,G19692,G19693,G19694,G19695,G19696,G19697,G19698,G19699,G19700,
       G19701,G19702,G19703,G19704,G19705,G19706,G19707,G19708,G19709,G19710,G19711,G19712,G19713,G19714,G19715,G19716,G19717,G19718,G19719,G19720,
       G19721,G19722,G19723,G19724,G19725,G19726,G19727,G19728,G19729,G19730,G19731,G19732,G19733,G19734,G19735,G19736,G19737,G19738,G19739,G19740,
       G19741,G19742,G19743,G19744,G19745,G19746,G19747,G19748,G19749,G19750,G19751,G19752,G19753,G19754,G19755,G19756,G19757,G19758,G19759,G19760,
       G19761,G19762,G19763,G19764,G19765,G19766,G19767,G19768,G19769,G19770,G19771,G19772,G19773,G19774,G19775,G19776,G19777,G19778,G19779,G19780,
       G19781,G19782,G19783,G19784,G19785,G19786,G19787,G19788,G19789,G19790,G19791,G19792,G19793,G19794,G19795,G19796,G19797,G19798,G19799,G19800,
       G19801,G19802,G19803,G19804,G19805,G19806,G19807,G19808,G19809,G19810,G19811,G19812,G19813,G19814,G19815,G19816,G19817,G19818,G19819,G19820,
       G19821,G19822,G19823,G19824,G19825,G19826,G19827,G19828,G19829,G19830,G19831,G19832,G19833,G19834,G19835,G19836,G19837,G19838,G19839,G19840,
       G19841,G19842,G19843,G19844,G19845,G19846,G19847,G19848,G19849,G19850,G19851,G19852,G19853,G19854,G19855,G19856,G19857,G19858,G19859,G19860,
       G19861,G19862,G19863,G19864,G19865,G19866,G19867,G19868,G19869,G19870,G19871,G19872,G19873,G19874,G19875,G19876,G19877,G19878,G19879,G19880,
       G19881,G19882,G19883,G19884,G19885,G19886,G19887,G19888,G19889,G19890,G19891,G19892,G19893,G19894,G19895,G19896,G19897,G19898,G19899,G19900,
       G19901,G19902,G19903,G19904,G19905,G19906,G19907,G19908,G19909,G19910,G19911,G19912,G19913,G19914,G19915,G19916,G19917,G19918,G19919,G19920,
       G19921,G19922,G19923,G19924,G19925,G19926,G19927,G19928,G19929,G19930,G19931,G19932,G19933,G19934,G19935,G19936,G19937,G19938,G19939,G19940,
       G19941,G19942,G19943,G19944,G19945,G19946,G19947,G19948,G19949,G19950,G19951,G19952,G19953,G19954,G19955,G19956,G19957,G19958,G19959,G19960,
       G19961,G19962,G19963,G19964,G19965,G19966,G19967,G19968,G19969,G19970,G19971,G19972,G19973,G19974,G19975,G19976,G19977,G19978,G19979,G19980,
       G19981,G19982,G19983,G19984,G19985,G19986,G19987,G19988,G19989,G19990,G19991,G19992,G19993,G19994,G19995,G19996,G19997,G19998,G19999,G20000,
       G20001,G20002,G20003,G20004,G20005,G20006,G20007,G20008,G20009,G20010,G20011,G20012,G20013,G20014,G20015,G20016,G20017,G20018,G20019,G20020,
       G20021,G20022,G20023,G20024,G20025,G20026,G20027,G20028,G20029,G20030,G20031,G20032,G20033,G20034,G20035,G20036,G20037,G20038,G20039,G20040,
       G20041,G20042,G20043,G20044,G20045,G20046,G20047,G20048,G20049,G20050,G20051,G20052,G20053,G20054,G20055,G20056,G20057,G20058,G20059,G20060,
       G20061,G20062,G20063,G20064,G20065,G20066,G20067,G20068,G20069,G20070,G20071,G20072,G20073,G20074,G20075,G20076,G20077,G20078,G20079,G20080,
       G20081,G20082,G20083,G20084,G20085,G20086,G20087,G20088,G20089,G20090,G20091,G20092,G20093,G20094,G20095,G20096,G20097,G20098,G20099,G20100,
       G20101,G20102,G20103,G20104,G20105,G20106,G20107,G20108,G20109,G20110,G20111,G20112,G20113,G20114,G20115,G20116,G20117,G20118,G20119,G20120,
       G20121,G20122,G20123,G20124,G20125,G20126,G20127,G20128,G20129,G20130,G20131,G20132,G20133,G20134,G20135,G20136,G20137,G20138,G20139,G20140,
       G20141,G20142,G20143,G20144,G20145,G20146,G20147,G20148,G20149,G20150,G20151,G20152,G20153,G20154,G20155,G20156,G20157,G20158,G20159,G20160,
       G20161,G20162,G20163,G20164,G20165,G20166,G20167,G20168,G20169,G20170,G20171,G20172,G20173,G20174,G20175,G20176,G20177,G20178,G20179,G20180,
       G20181,G20182,G20183,G20184,G20185,G20186,G20187,G20188,G20189,G20190,G20191,G20192,G20193,G20194,G20195,G20196,G20197,G20198,G20199,G20200,
       G20201,G20202,G20203,G20204,G20205,G20206,G20207,G20208,G20209,G20210,G20211,G20212,G20213,G20214,G20215,G20216,G20217,G20218,G20219,G20220,
       G20221,G20222,G20223,G20224,G20225,G20226,G20227,G20228,G20229,G20230,G20231,G20232,G20233,G20234,G20235,G20236,G20237,G20238,G20239,G20240,
       G20241,G20242,G20243,G20244,G20245,G20246,G20247,G20248,G20249,G20250,G20251,G20252,G20253,G20254,G20255,G20256,G20257,G20258,G20259,G20260,
       G20261,G20262,G20263,G20264,G20265,G20266,G20267,G20268,G20269,G20270,G20271,G20272,G20273,G20274,G20275,G20276,G20277,G20278,G20279,G20280,
       G20281,G20282,G20283,G20284,G20285,G20286,G20287,G20288,G20289,G20290,G20291,G20292,G20293,G20294,G20295,G20296,G20297,G20298,G20299,G20300,
       G20301,G20302,G20303,G20304,G20305,G20306,G20307,G20308,G20309,G20310,G20311,G20312,G20313,G20314,G20315,G20316,G20317,G20318,G20319,G20320,
       G20321,G20322,G20323,G20324,G20325,G20326,G20327,G20328,G20329,G20330,G20331,G20332,G20333,G20334,G20335,G20336,G20337,G20338,G20339,G20340,
       G20341,G20342,G20343,G20344,G20345,G20346,G20347,G20348,G20349,G20350,G20351,G20352,G20353,G20354,G20355,G20356,G20357,G20358,G20359,G20360,
       G20361,G20362,G20363,G20364,G20365,G20366,G20367,G20368,G20369,G20370,G20371,G20372,G20373,G20374,G20375,G20376,G20377,G20378,G20379,G20380,
       G20381,G20382,G20383,G20384,G20385,G20386,G20387,G20388,G20389,G20390,G20391,G20392,G20393,G20394,G20395,G20396,G20397,G20398,G20399,G20400,
       G20401,G20402,G20403,G20404,G20405,G20406,G20407,G20408,G20409,G20410,G20411,G20412,G20413,G20414,G20415,G20416,G20417,G20418,G20419,G20420,
       G20421,G20422,G20423,G20424,G20425,G20426,G20427,G20428,G20429,G20430,G20431,G20432,G20433,G20434,G20435,G20436,G20437,G20438,G20439,G20440,
       G20441,G20442,G20443,G20444,G20445,G20446,G20447,G20448,G20449,G20450,G20451,G20452,G20453,G20454,G20455,G20456,G20457,G20458,G20459,G20460,
       G20461,G20462,G20463,G20464,G20465,G20466,G20467,G20468,G20469,G20470,G20471,G20472,G20473,G20474,G20475,G20476,G20477,G20478,G20479,G20480,
       G20481,G20482,G20483,G20484,G20485,G20486,G20487,G20488,G20489,G20490,G20491,G20492,G20493,G20494,G20495,G20496,G20497,G20498,G20499,G20500,
       G20501,G20502,G20503,G20504,G20505,G20506,G20507,G20508,G20509,G20510,G20511,G20512,G20513,G20514,G20515,G20516,G20517,G20518,G20519,G20520,
       G20521,G20522,G20523,G20524,G20525,G20526,G20527,G20528,G20529,G20530,G20531,G20532,G20533,G20534,G20535,G20536,G20537,G20538,G20539,G20540,
       G20541,G20542,G20543,G20544,G20545,G20546,G20547,G20548,G20549,G20550,G20551,G20552,G20553,G20554,G20555,G20556,G20557,G20558,G20559,G20560,
       G20561,G20562,G20563,G20564,G20565,G20566,G20567,G20568,G20569,G20570,G20571,G20572,G20573,G20574,G20575,G20576,G20577,G20578,G20579,G20580,
       G20581,G20582,G20583,G20584,G20585,G20586,G20587,G20588,G20589,G20590,G20591,G20592,G20593,G20594,G20595,G20596,G20597,G20598,G20599,G20600,
       G20601,G20602,G20603,G20604,G20605,G20606,G20607,G20608,G20609,G20610,G20611,G20612,G20613,G20614,G20615,G20616,G20617,G20618,G20619,G20620,
       G20621,G20622,G20623,G20624,G20625,G20626,G20627,G20628,G20629,G20630,G20631,G20632,G20633,G20634,G20635,G20636,G20637,G20638,G20639,G20640,
       G20641,G20642,G20643,G20644,G20645,G20646,G20647,G20648,G20649,G20650,G20651,G20652,G20653,G20654,G20655,G20656,G20657,G20658,G20659,G20660,
       G20661,G20662,G20663,G20664,G20665,G20666,G20667,G20668,G20669,G20670,G20671,G20672,G20673,G20674,G20675,G20676,G20677,G20678,G20679,G20680,
       G20681,G20682,G20683,G20684,G20685,G20686,G20687,G20688,G20689,G20690,G20691,G20692,G20693,G20694,G20695,G20696,G20697,G20698,G20699,G20700,
       G20701,G20702,G20703,G20704,G20705,G20706,G20707,G20708,G20709,G20710,G20711,G20712,G20713,G20714,G20715,G20716,G20717,G20718,G20719,G20720,
       G20721,G20722,G20723,G20724,G20725,G20726,G20727,G20728,G20729,G20730,G20731,G20732,G20733,G20734,G20735,G20736,G20737,G20738,G20739,G20740,
       G20741,G20742,G20743,G20744,G20745,G20746,G20747,G20748,G20749,G20750,G20751,G20752,G20753,G20754,G20755,G20756,G20757,G20758,G20759,G20760,
       G20761,G20762,G20763,G20764,G20765,G20766,G20767,G20768,G20769,G20770,G20771,G20772,G20773,G20774,G20775,G20776,G20777,G20778,G20779,G20780,
       G20781,G20782,G20783,G20784,G20785,G20786,G20787,G20788,G20789,G20790,G20791,G20792,G20793,G20794,G20795,G20796,G20797,G20798,G20799,G20800,
       G20801,G20802,G20803,G20804,G20805,G20806,G20807,G20808,G20809,G20810,G20811,G20812,G20813,G20814,G20815,G20816,G20817,G20818,G20819,G20820,
       G20821,G20822,G20823,G20824,G20825,G20826,G20827,G20828,G20829,G20830,G20831,G20832,G20833,G20834,G20835,G20836,G20837,G20838,G20839,G20840,
       G20841,G20842,G20843,G20844,G20845,G20846,G20847,G20848,G20849,G20850,G20851,G20852,G20853,G20854,G20855,G20856,G20857,G20858,G20859,G20860,
       G20861,G20862,G20863,G20864,G20865,G20866,G20867,G20868,G20869,G20870,G20871,G20872,G20873,G20874,G20875,G20876,G20877,G20878,G20879,G20880,
       G20881,G20882,G20883,G20884,G20885,G20886,G20887,G20888,G20889,G20890,G20891,G20892,G20893,G20894,G20895,G20896,G20897,G20898,G20899,G20900,
       G20901,G20902,G20903,G20904,G20905,G20906,G20907,G20908,G20909,G20910,G20911,G20912,G20913,G20914,G20915,G20916,G20917,G20918,G20919,G20920,
       G20921,G20922,G20923,G20924,G20925,G20926,G20927,G20928,G20929,G20930,G20931,G20932,G20933,G20934,G20935,G20936,G20937,G20938,G20939,G20940,
       G20941,G20942,G20943,G20944,G20945,G20946,G20947,G20948,G20949,G20950,G20951,G20952,G20953,G20954,G20955,G20956,G20957,G20958,G20959,G20960,
       G20961,G20962,G20963,G20964,G20965,G20966,G20967,G20968,G20969,G20970,G20971,G20972,G20973,G20974,G20975,G20976,G20977,G20978,G20979,G20980,
       G20981,G20982,G20983,G20984,G20985,G20986,G20987,G20988,G20989,G20990,G20991,G20992,G20993,G20994,G20995,G20996,G20997,G20998,G20999,G21000,
       G21001,G21002,G21003,G21004,G21005,G21006,G21007,G21008,G21009,G21010,G21011,G21012,G21013,G21014,G21015,G21016,G21017,G21018,G21019,G21020,
       G21021,G21022,G21023,G21024,G21025,G21026,G21027,G21028,G21029,G21030,G21031,G21032,G21033,G21034,G21035,G21036,G21037,G21038,G21039,G21040,
       G21041,G21042,G21043,G21044,G21045,G21046,G21047,G21048,G21049,G21050,G21051,G21052,G21053,G21054,G21055,G21056,G21057,G21058,G21059,G21060,
       G21061,G21062,G21063,G21064,G21065,G21066,G21067,G21068,G21069,G21070,G21071,G21072,G21073,G21074,G21075,G21076,G21077,G21078,G21079,G21080,
       G21081,G21082,G21083,G21084,G21085,G21086,G21087,G21088,G21089,G21090,G21091,G21092,G21093,G21094,G21095,G21096,G21097,G21098,G21099,G21100,
       G21101,G21102,G21103,G21104,G21105,G21106,G21107,G21108,G21109,G21110,G21111,G21112,G21113,G21114,G21115,G21116,G21117,G21118,G21119,G21120,
       G21121,G21122,G21123,G21124,G21125,G21126,G21127,G21128,G21129,G21130,G21131,G21132,G21133,G21134,G21135,G21136,G21137,G21138,G21139,G21140,
       G21141,G21142,G21143,G21144,G21145,G21146,G21147,G21148,G21149,G21150,G21151,G21152,G21153,G21154,G21155,G21156,G21157,G21158,G21159,G21160,
       G21161,G21162,G21163,G21164,G21165,G21166,G21167,G21168,G21169,G21170,G21171,G21172,G21173,G21174,G21175,G21176,G21177,G21178,G21179,G21180,
       G21181,G21182,G21183,G21184,G21185,G21186,G21187,G21188,G21189,G21190,G21191,G21192,G21193,G21194,G21195,G21196,G21197,G21198,G21199,G21200,
       G21201,G21202,G21203,G21204,G21205,G21206,G21207,G21208,G21209,G21210,G21211,G21212,G21213,G21214,G21215,G21216,G21217,G21218,G21219,G21220,
       G21221,G21222,G21223,G21224,G21225,G21226,G21227,G21228,G21229,G21230,G21231,G21232,G21233,G21234,G21235,G21236,G21237,G21238,G21239,G21240,
       G21241,G21242,G21243,G21244,G21245,G21246,G21247,G21248,G21249,G21250,G21251,G21252,G21253,G21254,G21255,G21256,G21257,G21258,G21259,G21260,
       G21261,G21262,G21263,G21264,G21265,G21266,G21267,G21268,G21269,G21270,G21271,G21272,G21273,G21274,G21275,G21276,G21277,G21278,G21279,G21280,
       G21281,G21282,G21283,G21284,G21285,G21286,G21287,G21288,G21289,G21290,G21291,G21292,G21293,G21294,G21295,G21296,G21297,G21298,G21299,G21300,
       G21301,G21302,G21303,G21304,G21305,G21306,G21307,G21308,G21309,G21310,G21311,G21312,G21313,G21314,G21315,G21316,G21317,G21318,G21319,G21320,
       G21321,G21322,G21323,G21324,G21325,G21326,G21327,G21328,G21329,G21330,G21331,G21332,G21333,G21334,G21335,G21336,G21337,G21338,G21339,G21340,
       G21341,G21342,G21343,G21344,G21345,G21346,G21347,G21348,G21349,G21350,G21351,G21352,G21353,G21354,G21355,G21356,G21357,G21358,G21359,G21360,
       G21361,G21362,G21363,G21364,G21365,G21366,G21367,G21368,G21369,G21370,G21371,G21372,G21373,G21374,G21375,G21376,G21377,G21378,G21379,G21380,
       G21381,G21382,G21383,G21384,G21385,G21386,G21387,G21388,G21389,G21390,G21391,G21392,G21393,G21394,G21395,G21396,G21397,G21398,G21399,G21400,
       G21401,G21402,G21403,G21404,G21405,G21406,G21407,G21408,G21409,G21410,G21411,G21412,G21413,G21414,G21415,G21416,G21417,G21418,G21419,G21420,
       G21421,G21422,G21423,G21424,G21425,G21426,G21427,G21428,G21429,G21430,G21431,G21432,G21433,G21434,G21435,G21436,G21437,G21438,G21439,G21440,
       G21441,G21442,G21443,G21444,G21445,G21446,G21447,G21448,G21449,G21450,G21451,G21452,G21453,G21454,G21455,G21456,G21457,G21458,G21459,G21460,
       G21461,G21462,G21463,G21464,G21465,G21466,G21467,G21468,G21469,G21470,G21471,G21472,G21473,G21474,G21475,G21476,G21477,G21478,G21479,G21480,
       G21481,G21482,G21483,G21484,G21485,G21486,G21487,G21488,G21489,G21490,G21491,G21492,G21493,G21494,G21495,G21496,G21497,G21498,G21499,G21500,
       G21501,G21502,G21503,G21504,G21505,G21506,G21507,G21508,G21509,G21510,G21511,G21512,G21513,G21514,G21515,G21516,G21517,G21518,G21519,G21520,
       G21521,G21522,G21523,G21524,G21525,G21526,G21527,G21528,G21529,G21530,G21531,G21532,G21533,G21534,G21535,G21536,G21537,G21538,G21539,G21540,
       G21541,G21542,G21543,G21544,G21545,G21546,G21547,G21548,G21549,G21550,G21551,G21552,G21553,G21554,G21555,G21556,G21557,G21558,G21559,G21560,
       G21561,G21562,G21563,G21564,G21565,G21566,G21567,G21568,G21569,G21570,G21571,G21572,G21573,G21574,G21575,G21576,G21577,G21578,G21579,G21580,
       G21581,G21582,G21583,G21584,G21585,G21586,G21587,G21588,G21589,G21590,G21591,G21592,G21593,G21594,G21595,G21596,G21597,G21598,G21599,G21600,
       G21601,G21602,G21603,G21604,G21605,G21606,G21607,G21608,G21609,G21610,G21611,G21612,G21613,G21614,G21615,G21616,G21617,G21618,G21619,G21620,
       G21621,G21622,G21623,G21624,G21625,G21626,G21627,G21628,G21629,G21630,G21631,G21632,G21633,G21634,G21635,G21636,G21637,G21638,G21639,G21640,
       G21641,G21642,G21643,G21644,G21645,G21646,G21647,G21648,G21649,G21650,G21651,G21652,G21653,G21654,G21655,G21656,G21657,G21658,G21659,G21660,
       G21661,G21662,G21663,G21664,G21665,G21666,G21667,G21668,G21669,G21670,G21671,G21672,G21673,G21674,G21675,G21676,G21677,G21678,G21679,G21680,
       G21681,G21682,G21683,G21684,G21685,G21686,G21687,G21688,G21689,G21690,G21691,G21692,G21693,G21694,G21695,G21696,G21697,G21698,G21699,G21700,
       G21701,G21702,G21703,G21704,G21705,G21706,G21707,G21708,G21709,G21710,G21711,G21712,G21713,G21714,G21715,G21716,G21717,G21718,G21719,G21720,
       G21721,G21722,G21723,G21724,G21725,G21726,G21727,G21728,G21729,G21730,G21731,G21732,G21733,G21734,G21735,G21736,G21737,G21738,G21739,G21740,
       G21741,G21742,G21743,G21744,G21745,G21746,G21747,G21748,G21749,G21750,G21751,G21752,G21753,G21754,G21755,G21756,G21757,G21758,G21759,G21760,
       G21761,G21762,G21763,G21764,G21765,G21766,G21767,G21768,G21769,G21770,G21771,G21772,G21773,G21774,G21775,G21776,G21777,G21778,G21779,G21780,
       G21781,G21782,G21783,G21784,G21785,G21786,G21787,G21788,G21789,G21790,G21791,G21792,G21793,G21794,G21795,G21796,G21797,G21798,G21799,G21800,
       G21801,G21802,G21803,G21804,G21805,G21806,G21807,G21808,G21809,G21810,G21811,G21812,G21813,G21814,G21815,G21816,G21817,G21818,G21819,G21820,
       G21821,G21822,G21823,G21824,G21825,G21826,G21827,G21828,G21829,G21830,G21831,G21832,G21833,G21834,G21835,G21836,G21837,G21838,G21839,G21840,
       G21841,G21842,G21843,G21844,G21845,G21846,G21847,G21848,G21849,G21850,G21851,G21852,G21853,G21854,G21855,G21856,G21857,G21858,G21859,G21860,
       G21861,G21862,G21863,G21864,G21865,G21866,G21867,G21868,G21869,G21870,G21871,G21872,G21873,G21874,G21875,G21876,G21877,G21878,G21879,G21880,
       G21881,G21882,G21883,G21884,G21885,G21886,G21887,G21888,G21889,G21890,G21891,G21892,G21893,G21894,G21895,G21896,G21897,G21898,G21899,G21900,
       G21901,G21902,G21903,G21904,G21905,G21906,G21907,G21908,G21909,G21910,G21911,G21912,G21913,G21914,G21915,G21916,G21917,G21918,G21919,G21920,
       G21921,G21922,G21923,G21924,G21925,G21926,G21927,G21928,G21929,G21930,G21931,G21932,G21933,G21934,G21935,G21936,G21937,G21938,G21939,G21940,
       G21941,G21942,G21943,G21944,G21945,G21946,G21947,G21948,G21949,G21950,G21951,G21952,G21953,G21954,G21955,G21956,G21957,G21958,G21959,G21960,
       G21961,G21962,G21963,G21964,G21965,G21966,G21967,G21968,G21969,G21970,G21971,G21972,G21973,G21974,G21975,G21976,G21977,G21978,G21979,G21980,
       G21981,G21982,G21983,G21984,G21985,G21986,G21987,G21988,G21989,G21990,G21991,G21992,G21993,G21994,G21995,G21996,G21997,G21998,G21999,G22000,
       G22001,G22002,G22003,G22004,G22005,G22006,G22007,G22008,G22009,G22010,G22011,G22012,G22013,G22014,G22015,G22016,G22017,G22018,G22019,G22020,
       G22021,G22022,G22023,G22024,G22025,G22026,G22027,G22028,G22029,G22030,G22031,G22032,G22033,G22034,G22035,G22036,G22037,G22038,G22039,G22040,
       G22041,G22042,G22043,G22044,G22045,G22046,G22047,G22048,G22049,G22050,G22051,G22052,G22053,G22054,G22055,G22056,G22057,G22058,G22059,G22060,
       G22061,G22062,G22063,G22064,G22065,G22066,G22067,G22068,G22069,G22070,G22071,G22072,G22073,G22074,G22075,G22076,G22077,G22078,G22079,G22080,
       G22081,G22082,G22083,G22084,G22085,G22086,G22087,G22088,G22089,G22090,G22091,G22092,G22093,G22094,G22095,G22096,G22097,G22098,G22099,G22100,
       G22101,G22102,G22103,G22104,G22105,G22106,G22107,G22108,G22109,G22110,G22111,G22112,G22113,G22114,G22115,G22116,G22117,G22118,G22119,G22120,
       G22121,G22122,G22123,G22124,G22125,G22126,G22127,G22128,G22129,G22130,G22131,G22132,G22133,G22134,G22135,G22136,G22137,G22138,G22139,G22140,
       G22141,G22142,G22143,G22144,G22145,G22146,G22147,G22148,G22149,G22150,G22151,G22152,G22153,G22154,G22155,G22156,G22157,G22158,G22159,G22160,
       G22161,G22162,G22163,G22164,G22165,G22166,G22167,G22168,G22169,G22170,G22171,G22172,G22173,G22174,G22175,G22176,G22177,G22178,G22179,G22180,
       G22181,G22182,G22183,G22184,G22185,G22186,G22187,G22188,G22189,G22190,G22191,G22192,G22193,G22194,G22195,G22196,G22197,G22198,G22199,G22200,
       G22201,G22202,G22203,G22204,G22205,G22206,G22207,G22208,G22209,G22210,G22211,G22212,G22213,G22214,G22215,G22216,G22217,G22218,G22219,G22220,
       G22221,G22222,G22223,G22224,G22225,G22226,G22227,G22228,G22229,G22230,G22231,G22232,G22233,G22234,G22235,G22236,G22237,G22238,G22239,G22240,
       G22241,G22242,G22243,G22244,G22245,G22246,G22247,G22248,G22249,G22250,G22251,G22252,G22253,G22254,G22255,G22256,G22257,G22258,G22259,G22260,
       G22261,G22262,G22263,G22264,G22265,G22266,G22267,G22268,G22269,G22270,G22271,G22272,G22273,G22274,G22275,G22276,G22277,G22278,G22279,G22280,
       G22281,G22282,G22283,G22284,G22285,G22286,G22287,G22288,G22289,G22290,G22291,G22292,G22293,G22294,G22295,G22296,G22297,G22298,G22299,G22300,
       G22301,G22302,G22303,G22304,G22305,G22306,G22307,G22308,G22309,G22310,G22311,G22312,G22313,G22314,G22315,G22316,G22317,G22318,G22319,G22320,
       G22321,G22322,G22323,G22324,G22325,G22326,G22327,G22328,G22329,G22330,G22331,G22332,G22333,G22334,G22335,G22336,G22337,G22338,G22339,G22340,
       G22341,G22342,G22343,G22344,G22345,G22346,G22347,G22348,G22349,G22350,G22351,G22352,G22353,G22354,G22355,G22356,G22357,G22358,G22359,G22360,
       G22361,G22362,G22363,G22364,G22365,G22366,G22367,G22368,G22369,G22370,G22371,G22372,G22373,G22374,G22375,G22376,G22377,G22378,G22379,G22380,
       G22381,G22382,G22383,G22384,G22385,G22386,G22387,G22388,G22389,G22390,G22391,G22392,G22393,G22394,G22395,G22396,G22397,G22398,G22399,G22400,
       G22401,G22402,G22403,G22404,G22405,G22406,G22407,G22408,G22409,G22410,G22411,G22412,G22413,G22414,G22415,G22416,G22417,G22418,G22419,G22420,
       G22421,G22422,G22423,G22424,G22425,G22426,G22427,G22428,G22429,G22430,G22431,G22432,G22433,G22434,G22435,G22436,G22437,G22438,G22439,G22440,
       G22441,G22442,G22443,G22444,G22445,G22446,G22447,G22448,G22449,G22450,G22451,G22452,G22453,G22454,G22455,G22456,G22457,G22458,G22459,G22460,
       G22461,G22462,G22463,G22464,G22465,G22466,G22467,G22468,G22469,G22470,G22471,G22472,G22473,G22474,G22475,G22476,G22477,G22478,G22479,G22480,
       G22481,G22482,G22483,G22484,G22485,G22486,G22487,G22488,G22489,G22490,G22491,G22492,G22493,G22494,G22495,G22496,G22497,G22498,G22499,G22500,
       G22501,G22502,G22503,G22504,G22505,G22506,G22507,G22508,G22509,G22510,G22511,G22512,G22513,G22514,G22515,G22516,G22517,G22518,G22519,G22520,
       G22521,G22522,G22523,G22524,G22525,G22526,G22527,G22528,G22529,G22530,G22531,G22532,G22533,G22534,G22535,G22536,G22537,G22538,G22539,G22540,
       G22541,G22542,G22543,G22544,G22545,G22546,G22547,G22548,G22549,G22550,G22551,G22552,G22553,G22554,G22555,G22556,G22557,G22558,G22559,G22560,
       G22561,G22562,G22563,G22564,G22565,G22566,G22567,G22568,G22569,G22570,G22571,G22572,G22573,G22574,G22575,G22576,G22577,G22578,G22579,G22580,
       G22581,G22582,G22583,G22584,G22585,G22586,G22587,G22588,G22589,G22590,G22591,G22592,G22593,G22594,G22595,G22596,G22597,G22598,G22599,G22600,
       G22601,G22602,G22603,G22604,G22605,G22606,G22607,G22608,G22609,G22610,G22611,G22612,G22613,G22614,G22615,G22616,G22617,G22618,G22619,G22620,
       G22621,G22622,G22623,G22624,G22625,G22626,G22627,G22628,G22629,G22630,G22631,G22632,G22633,G22634,G22635,G22636,G22637,G22638,G22639,G22640,
       G22641,G22642,G22643,G22644,G22645,G22646,G22647,G22648,G22649,G22650,G22651,G22652,G22653,G22654,G22655,G22656,G22657,G22658,G22659,G22660,
       G22661,G22662,G22663,G22664,G22665,G22666,G22667,G22668,G22669,G22670,G22671,G22672,G22673,G22674,G22675,G22676,G22677,G22678,G22679,G22680,
       G22681,G22682,G22683,G22684,G22685,G22686,G22687,G22688,G22689,G22690,G22691,G22692,G22693,G22694,G22695,G22696,G22697,G22698,G22699,G22700,
       G22701,G22702,G22703,G22704,G22705,G22706,G22707,G22708,G22709,G22710,G22711,G22712,G22713,G22714,G22715,G22716,G22717,G22718,G22719,G22720,
       G22721,G22722,G22723,G22724,G22725,G22726,G22727,G22728,G22729,G22730,G22731,G22732,G22733,G22734,G22735,G22736,G22737,G22738,G22739,G22740,
       G22741,G22742,G22743,G22744,G22745,G22746,G22747,G22748,G22749,G22750,G22751,G22752,G22753,G22754,G22755,G22756,G22757,G22758,G22759,G22760,
       G22761,G22762,G22763,G22764,G22765,G22766,G22767,G22768,G22769,G22770,G22771,G22772,G22773,G22774,G22775,G22776,G22777,G22778,G22779,G22780,
       G22781,G22782,G22783,G22784,G22785,G22786,G22787,G22788,G22789,G22790,G22791,G22792,G22793,G22794,G22795,G22796,G22797,G22798,G22799,G22800,
       G22801,G22802,G22803,G22804,G22805,G22806,G22807,G22808,G22809,G22810,G22811,G22812,G22813,G22814,G22815,G22816,G22817,G22818,G22819,G22820,
       G22821,G22822,G22823,G22824,G22825,G22826,G22827,G22828,G22829,G22830,G22831,G22832,G22833,G22834,G22835,G22836,G22837,G22838,G22839,G22840,
       G22841,G22842,G22843,G22844,G22845,G22846,G22847,G22848,G22849,G22850,G22851,G22852,G22853,G22854,G22855,G22856,G22857,G22858,G22859,G22860,
       G22861,G22862,G22863,G22864,G22865,G22866,G22867,G22868,G22869,G22870,G22871,G22872,G22873,G22874,G22875,G22876,G22877,G22878,G22879,G22880,
       G22881,G22882,G22883,G22884,G22885,G22886,G22887,G22888,G22889,G22890,G22891,G22892,G22893,G22894,G22895,G22896,G22897,G22898,G22899,G22900,
       G22901,G22902,G22903,G22904,G22905,G22906,G22907,G22908,G22909,G22910,G22911,G22912,G22913,G22914,G22915,G22916,G22917,G22918,G22919,G22920,
       G22921,G22922,G22923,G22924,G22925,G22926,G22927,G22928,G22929,G22930,G22931,G22932,G22933,G22934,G22935,G22936,G22937,G22938,G22939,G22940,
       G22941,G22942,G22943,G22944,G22945,G22946,G22947,G22948,G22949,G22950,G22951,G22952,G22953,G22954,G22955,G22956,G22957,G22958,G22959,G22960,
       G22961,G22962,G22963,G22964,G22965,G22966,G22967,G22968,G22969,G22970,G22971,G22972,G22973,G22974,G22975,G22976,G22977,G22978,G22979,G22980,
       G22981,G22982,G22983,G22984,G22985,G22986,G22987,G22988,G22989,G22990,G22991,G22992,G22993,G22994,G22995,G22996,G22997,G22998,G22999,G23000,
       G23001,G23002,G23003,G23004,G23005,G23006,G23007,G23008,G23009,G23010,G23011,G23012,G23013,G23014,G23015,G23016,G23017,G23018,G23019,G23020,
       G23021,G23022,G23023,G23024,G23025,G23026,G23027,G23028,G23029,G23030,G23031,G23032,G23033,G23034,G23035,G23036,G23037,G23038,G23039,G23040,
       G23041,G23042,G23043,G23044,G23045;

  dff DFF_55(CK,G22556,G1067);
  dff DFF_56(CK,G22557,G1068);
  dff DFF_57(CK,G22558,G1069);
  dff DFF_58(CK,G22559,G1070);
  dff DFF_59(CK,G22560,G1071);
  dff DFF_60(CK,G22561,G1072);
  dff DFF_61(CK,G22562,G1073);
  dff DFF_62(CK,G22563,G1074);
  dff DFF_63(CK,G22564,G1075);
  dff DFF_64(CK,G22565,G1076);
  dff DFF_65(CK,G22566,G1077);
  dff DFF_66(CK,G22567,G1078);
  dff DFF_67(CK,G22568,G1079);
  dff DFF_68(CK,G22569,G1080);
  dff DFF_69(CK,G22570,G1081);
  dff DFF_70(CK,G22571,G1082);
  dff DFF_71(CK,G22572,G1083);
  dff DFF_72(CK,G22573,G1084);
  dff DFF_73(CK,G22574,G1085);
  dff DFF_74(CK,G22575,G1086);
  dff DFF_75(CK,G22576,G1087);
  dff DFF_76(CK,G22577,G1088);
  dff DFF_77(CK,G22578,G1089);
  dff DFF_78(CK,G22579,G1090);
  dff DFF_79(CK,G22580,G1091);
  dff DFF_80(CK,G22581,G1092);
  dff DFF_81(CK,G22582,G1093);
  dff DFF_82(CK,G22583,G1094);
  dff DFF_83(CK,G22584,G1095);
  dff DFF_84(CK,G22585,G1096);
  dff DFF_85(CK,G22586,G1097);
  dff DFF_86(CK,G22587,G1098);
  dff DFF_87(CK,G22588,G1523);
  dff DFF_88(CK,G22589,G1522);
  dff DFF_89(CK,G22590,G1099);
  dff DFF_90(CK,G22591,G1100);
  dff DFF_91(CK,G22592,G1101);
  dff DFF_92(CK,G22593,G1102);
  dff DFF_93(CK,G22594,G1103);
  dff DFF_94(CK,G22595,G1104);
  dff DFF_95(CK,G22596,G1105);
  dff DFF_96(CK,G22597,G1106);
  dff DFF_97(CK,G22598,G1107);
  dff DFF_98(CK,G22599,G1108);
  dff DFF_99(CK,G22600,G1109);
  dff DFF_100(CK,G22601,G1110);
  dff DFF_101(CK,G22602,G1111);
  dff DFF_102(CK,G22603,G1112);
  dff DFF_103(CK,G22604,G1113);
  dff DFF_104(CK,G22605,G1114);
  dff DFF_105(CK,G22606,G1115);
  dff DFF_106(CK,G22607,G1116);
  dff DFF_107(CK,G22608,G1117);
  dff DFF_108(CK,G22609,G1118);
  dff DFF_109(CK,G22610,G1119);
  dff DFF_110(CK,G22611,G1120);
  dff DFF_111(CK,G22612,G1121);
  dff DFF_112(CK,G22613,G1122);
  dff DFF_113(CK,G22614,G1123);
  dff DFF_114(CK,G22615,G1124);
  dff DFF_115(CK,G22616,G1125);
  dff DFF_116(CK,G22617,G1126);
  dff DFF_117(CK,G22618,G1127);
  dff DFF_118(CK,G22619,G1128);
  dff DFF_119(CK,G22620,G1521);
  dff DFF_120(CK,G22621,G1520);
  dff DFF_121(CK,G22622,G1519);
  dff DFF_122(CK,G22623,G1518);
  dff DFF_123(CK,G22624,G1517);
  dff DFF_124(CK,G22625,G1516);
  dff DFF_125(CK,G22626,G1515);
  dff DFF_126(CK,G22627,G1514);
  dff DFF_127(CK,G22628,G1513);
  dff DFF_128(CK,G22629,G1512);
  dff DFF_129(CK,G22630,G1511);
  dff DFF_130(CK,G22631,G1510);
  dff DFF_131(CK,G22632,G1509);
  dff DFF_132(CK,G22633,G1508);
  dff DFF_133(CK,G22634,G1507);
  dff DFF_134(CK,G22635,G1506);
  dff DFF_135(CK,G22636,G1505);
  dff DFF_136(CK,G22637,G1504);
  dff DFF_137(CK,G22638,G1503);
  dff DFF_138(CK,G22639,G1502);
  dff DFF_139(CK,G22640,G1501);
  dff DFF_140(CK,G22641,G1500);
  dff DFF_141(CK,G22642,G1499);
  dff DFF_142(CK,G22643,G1498);
  dff DFF_143(CK,G22644,G1497);
  dff DFF_144(CK,G22645,G1496);
  dff DFF_145(CK,G22646,G1495);
  dff DFF_146(CK,G22647,G1494);
  dff DFF_147(CK,G22648,G1493);
  dff DFF_148(CK,G22649,G1492);
  dff DFF_149(CK,G22650,G1491);
  dff DFF_150(CK,G22651,G1490);
  dff DFF_151(CK,G22652,G1489);
  dff DFF_152(CK,G22653,G1488);
  dff DFF_153(CK,G22654,G1487);
  dff DFF_154(CK,G22655,G1486);
  dff DFF_155(CK,G22656,G1485);
  dff DFF_156(CK,G22657,G1484);
  dff DFF_157(CK,G22658,G1483);
  dff DFF_158(CK,G22659,G1482);
  dff DFF_159(CK,G22660,G1481);
  dff DFF_160(CK,G22661,G1480);
  dff DFF_161(CK,G22662,G1479);
  dff DFF_162(CK,G22663,G1478);
  dff DFF_163(CK,G22664,G1477);
  dff DFF_164(CK,G22665,G1476);
  dff DFF_165(CK,G22666,G1475);
  dff DFF_166(CK,G22667,G1474);
  dff DFF_167(CK,G22668,G1473);
  dff DFF_168(CK,G22669,G1472);
  dff DFF_169(CK,G22670,G1471);
  dff DFF_170(CK,G22671,G1470);
  dff DFF_171(CK,G22672,G1469);
  dff DFF_172(CK,G22673,G1468);
  dff DFF_173(CK,G22674,G1467);
  dff DFF_174(CK,G22675,G1466);
  dff DFF_175(CK,G22676,G1465);
  dff DFF_176(CK,G22677,G1464);
  dff DFF_177(CK,G22678,G1463);
  dff DFF_178(CK,G22679,G1462);
  dff DFF_179(CK,G22680,G1461);
  dff DFF_180(CK,G22681,G1460);
  dff DFF_181(CK,G22682,G1459);
  dff DFF_182(CK,G22683,G1458);
  dff DFF_183(CK,G22684,G1129);
  dff DFF_184(CK,G22685,G1457);
  dff DFF_185(CK,G22686,G1130);
  dff DFF_186(CK,G22687,G1131);
  dff DFF_187(CK,G22688,G1132);
  dff DFF_188(CK,G22689,G1133);
  dff DFF_189(CK,G22690,G1134);
  dff DFF_190(CK,G22691,G1135);
  dff DFF_191(CK,G22692,G1136);
  dff DFF_192(CK,G22693,G1137);
  dff DFF_193(CK,G22694,G1138);
  dff DFF_194(CK,G22695,G1139);
  dff DFF_195(CK,G22696,G1140);
  dff DFF_196(CK,G22697,G1141);
  dff DFF_197(CK,G22698,G1142);
  dff DFF_198(CK,G22699,G1143);
  dff DFF_199(CK,G22700,G1144);
  dff DFF_200(CK,G22701,G1145);
  dff DFF_201(CK,G22702,G1146);
  dff DFF_202(CK,G22703,G1147);
  dff DFF_203(CK,G22704,G1148);
  dff DFF_204(CK,G22705,G1149);
  dff DFF_205(CK,G22706,G1150);
  dff DFF_206(CK,G22707,G1151);
  dff DFF_207(CK,G22708,G1152);
  dff DFF_208(CK,G22709,G1153);
  dff DFF_209(CK,G22710,G1154);
  dff DFF_210(CK,G22711,G1155);
  dff DFF_211(CK,G22712,G1156);
  dff DFF_212(CK,G22713,G1157);
  dff DFF_213(CK,G22714,G1158);
  dff DFF_214(CK,G22715,G1159);
  dff DFF_215(CK,G22716,G1160);
  dff DFF_216(CK,G22717,G1161);
  dff DFF_217(CK,G22718,G1162);
  dff DFF_218(CK,G22719,G1163);
  dff DFF_219(CK,G22720,G1164);
  dff DFF_220(CK,G22721,G1165);
  dff DFF_221(CK,G22722,G1166);
  dff DFF_222(CK,G22723,G1167);
  dff DFF_223(CK,G22724,G1168);
  dff DFF_224(CK,G22725,G1169);
  dff DFF_225(CK,G22726,G1170);
  dff DFF_226(CK,G22727,G1171);
  dff DFF_227(CK,G22728,G1172);
  dff DFF_228(CK,G22729,G1173);
  dff DFF_229(CK,G22730,G1174);
  dff DFF_230(CK,G22731,G1175);
  dff DFF_231(CK,G22732,G1176);
  dff DFF_232(CK,G22733,G1177);
  dff DFF_233(CK,G22734,G1178);
  dff DFF_234(CK,G22735,G1179);
  dff DFF_235(CK,G22736,G1456);
  dff DFF_236(CK,G22737,G1455);
  dff DFF_237(CK,G22738,G1454);
  dff DFF_238(CK,G22739,G1453);
  dff DFF_239(CK,G22740,G1452);
  dff DFF_240(CK,G22741,G1451);
  dff DFF_241(CK,G22742,G1450);
  dff DFF_242(CK,G22743,G1449);
  dff DFF_243(CK,G22744,G1448);
  dff DFF_244(CK,G22745,G1447);
  dff DFF_245(CK,G22746,G1446);
  dff DFF_246(CK,G22747,G1445);
  dff DFF_247(CK,G22748,G1444);
  dff DFF_248(CK,G22749,G1443);
  dff DFF_249(CK,G22750,G1442);
  dff DFF_250(CK,G22751,G1441);
  dff DFF_251(CK,G22752,G1440);
  dff DFF_252(CK,G22753,G1439);
  dff DFF_253(CK,G22754,G1438);
  dff DFF_254(CK,G22755,G1437);
  dff DFF_255(CK,G22756,G1436);
  dff DFF_256(CK,G22757,G1435);
  dff DFF_257(CK,G22758,G1434);
  dff DFF_258(CK,G22759,G1433);
  dff DFF_259(CK,G22760,G1432);
  dff DFF_260(CK,G22761,G1431);
  dff DFF_261(CK,G22762,G1430);
  dff DFF_262(CK,G22763,G1429);
  dff DFF_263(CK,G22764,G1428);
  dff DFF_264(CK,G22765,G1427);
  dff DFF_265(CK,G22766,G1426);
  dff DFF_266(CK,G22767,G1425);
  dff DFF_267(CK,G22768,G1180);
  dff DFF_268(CK,G22769,G1181);
  dff DFF_269(CK,G22770,G1182);
  dff DFF_270(CK,G22771,G1183);
  dff DFF_271(CK,G22772,G1184);
  dff DFF_272(CK,G22773,G1185);
  dff DFF_273(CK,G22774,G1186);
  dff DFF_274(CK,G22775,G1187);
  dff DFF_275(CK,G22776,G1188);
  dff DFF_276(CK,G22777,G1189);
  dff DFF_277(CK,G22778,G1190);
  dff DFF_278(CK,G22779,G1191);
  dff DFF_279(CK,G22780,G1192);
  dff DFF_280(CK,G22781,G1193);
  dff DFF_281(CK,G22782,G1194);
  dff DFF_282(CK,G22783,G1195);
  dff DFF_283(CK,G22784,G1196);
  dff DFF_284(CK,G22785,G1197);
  dff DFF_285(CK,G22786,G1198);
  dff DFF_286(CK,G22787,G1199);
  dff DFF_287(CK,G22788,G1200);
  dff DFF_288(CK,G22789,G1201);
  dff DFF_289(CK,G22790,G1202);
  dff DFF_290(CK,G22791,G1203);
  dff DFF_291(CK,G22792,G1204);
  dff DFF_292(CK,G22793,G1205);
  dff DFF_293(CK,G22794,G1206);
  dff DFF_294(CK,G22795,G1207);
  dff DFF_295(CK,G22796,G1208);
  dff DFF_296(CK,G22797,G1209);
  dff DFF_297(CK,G22798,G1066);
  dff DFF_298(CK,G22799,G1001);
  dff DFF_299(CK,G22800,G1290);
  dff DFF_300(CK,G22801,G3842);
  dff DFF_301(CK,G22802,G3843);
  dff DFF_302(CK,G22803,G3844);
  dff DFF_303(CK,G22804,G3845);
  dff DFF_304(CK,G22805,G3846);
  dff DFF_305(CK,G22806,G3847);
  dff DFF_306(CK,G22807,G3848);
  dff DFF_307(CK,G22808,G3849);
  dff DFF_308(CK,G22809,G3850);
  dff DFF_309(CK,G22810,G3851);
  dff DFF_310(CK,G22811,G3852);
  dff DFF_311(CK,G22812,G3853);
  dff DFF_312(CK,G22813,G3854);
  dff DFF_313(CK,G22814,G3855);
  dff DFF_314(CK,G22815,G3856);
  dff DFF_315(CK,G22816,G3857);
  dff DFF_316(CK,G22817,G3858);
  dff DFF_317(CK,G22818,G3859);
  dff DFF_318(CK,G22819,G3860);
  dff DFF_319(CK,G22820,G3861);
  dff DFF_320(CK,G22821,G3862);
  dff DFF_321(CK,G22822,G3863);
  dff DFF_322(CK,G22823,G3864);
  dff DFF_323(CK,G22824,G3865);
  dff DFF_324(CK,G22825,G3866);
  dff DFF_325(CK,G22826,G3867);
  dff DFF_326(CK,G22827,G3868);
  dff DFF_327(CK,G22828,G3869);
  dff DFF_328(CK,G22829,G3870);
  dff DFF_329(CK,G22830,G3871);
  dff DFF_330(CK,G22831,G3872);
  dff DFF_331(CK,G22832,G3873);
  dff DFF_332(CK,G22833,G4231);
  dff DFF_333(CK,G22834,G4230);
  dff DFF_334(CK,G22835,G3874);
  dff DFF_335(CK,G22836,G3875);
  dff DFF_336(CK,G22837,G3876);
  dff DFF_337(CK,G22838,G3877);
  dff DFF_338(CK,G22839,G3878);
  dff DFF_339(CK,G22840,G3879);
  dff DFF_340(CK,G22841,G3880);
  dff DFF_341(CK,G22842,G3881);
  dff DFF_342(CK,G22843,G3882);
  dff DFF_343(CK,G22844,G3883);
  dff DFF_344(CK,G22845,G3884);
  dff DFF_345(CK,G22846,G3885);
  dff DFF_346(CK,G22847,G3886);
  dff DFF_347(CK,G22848,G3887);
  dff DFF_348(CK,G22849,G3888);
  dff DFF_349(CK,G22850,G3889);
  dff DFF_350(CK,G22851,G3890);
  dff DFF_351(CK,G22852,G3891);
  dff DFF_352(CK,G22853,G3892);
  dff DFF_353(CK,G22854,G3893);
  dff DFF_354(CK,G22855,G3894);
  dff DFF_355(CK,G22856,G3895);
  dff DFF_356(CK,G22857,G3896);
  dff DFF_357(CK,G22858,G3897);
  dff DFF_358(CK,G22859,G3898);
  dff DFF_359(CK,G22860,G3899);
  dff DFF_360(CK,G22861,G3900);
  dff DFF_361(CK,G22862,G3901);
  dff DFF_362(CK,G22863,G3902);
  dff DFF_363(CK,G22864,G3903);
  dff DFF_364(CK,G22865,G3904);
  dff DFF_365(CK,G22866,G3905);
  dff DFF_366(CK,G22867,G3906);
  dff DFF_367(CK,G22868,G3907);
  dff DFF_368(CK,G22869,G3908);
  dff DFF_369(CK,G22870,G3909);
  dff DFF_370(CK,G22871,G3910);
  dff DFF_371(CK,G22872,G3911);
  dff DFF_372(CK,G22873,G3912);
  dff DFF_373(CK,G22874,G3913);
  dff DFF_374(CK,G22875,G3914);
  dff DFF_375(CK,G22876,G3915);
  dff DFF_376(CK,G22877,G3916);
  dff DFF_377(CK,G22878,G3917);
  dff DFF_378(CK,G22879,G3918);
  dff DFF_379(CK,G22880,G3919);
  dff DFF_380(CK,G22881,G3920);
  dff DFF_381(CK,G22882,G3921);
  dff DFF_382(CK,G22883,G3922);
  dff DFF_383(CK,G22884,G3923);
  dff DFF_384(CK,G22885,G3924);
  dff DFF_385(CK,G22886,G3925);
  dff DFF_386(CK,G22887,G3926);
  dff DFF_387(CK,G22888,G3927);
  dff DFF_388(CK,G22889,G3928);
  dff DFF_389(CK,G22890,G3929);
  dff DFF_390(CK,G22891,G3930);
  dff DFF_391(CK,G22892,G3931);
  dff DFF_392(CK,G22893,G3932);
  dff DFF_393(CK,G22894,G3933);
  dff DFF_394(CK,G22895,G3934);
  dff DFF_395(CK,G22896,G3935);
  dff DFF_396(CK,G22897,G3936);
  dff DFF_397(CK,G22898,G3937);
  dff DFF_398(CK,G22899,G3938);
  dff DFF_399(CK,G22900,G3939);
  dff DFF_400(CK,G22901,G3940);
  dff DFF_401(CK,G22902,G3941);
  dff DFF_402(CK,G22903,G3942);
  dff DFF_403(CK,G22904,G3943);
  dff DFF_404(CK,G22905,G3944);
  dff DFF_405(CK,G22906,G3945);
  dff DFF_406(CK,G22907,G3946);
  dff DFF_407(CK,G22908,G3947);
  dff DFF_408(CK,G22909,G3948);
  dff DFF_409(CK,G22910,G3949);
  dff DFF_410(CK,G22911,G3950);
  dff DFF_411(CK,G22912,G3951);
  dff DFF_412(CK,G22913,G3952);
  dff DFF_413(CK,G22914,G3953);
  dff DFF_414(CK,G22915,G3954);
  dff DFF_415(CK,G22916,G3955);
  dff DFF_416(CK,G22917,G3956);
  dff DFF_417(CK,G22918,G3957);
  dff DFF_418(CK,G22919,G3958);
  dff DFF_419(CK,G22920,G3959);
  dff DFF_420(CK,G22921,G3960);
  dff DFF_421(CK,G22922,G3961);
  dff DFF_422(CK,G22923,G3962);
  dff DFF_423(CK,G22924,G3963);
  dff DFF_424(CK,G22925,G3964);
  dff DFF_425(CK,G22926,G3965);
  dff DFF_426(CK,G22927,G3966);
  dff DFF_427(CK,G22928,G3967);
  dff DFF_428(CK,G22929,G3968);
  dff DFF_429(CK,G22930,G3969);
  dff DFF_430(CK,G22931,G3970);
  dff DFF_431(CK,G22932,G3971);
  dff DFF_432(CK,G22933,G3972);
  dff DFF_433(CK,G22934,G3973);
  dff DFF_434(CK,G22935,G3974);
  dff DFF_435(CK,G22936,G3975);
  dff DFF_436(CK,G22937,G3976);
  dff DFF_437(CK,G22938,G3977);
  dff DFF_438(CK,G22939,G3978);
  dff DFF_439(CK,G22940,G3979);
  dff DFF_440(CK,G22941,G3980);
  dff DFF_441(CK,G22942,G3981);
  dff DFF_442(CK,G22943,G3982);
  dff DFF_443(CK,G22944,G3983);
  dff DFF_444(CK,G22945,G3984);
  dff DFF_445(CK,G22946,G3985);
  dff DFF_446(CK,G22947,G3986);
  dff DFF_447(CK,G22948,G3987);
  dff DFF_448(CK,G22949,G3988);
  dff DFF_449(CK,G22950,G3989);
  dff DFF_450(CK,G22951,G3990);
  dff DFF_451(CK,G22952,G3991);
  dff DFF_452(CK,G22953,G3992);
  dff DFF_453(CK,G22954,G3993);
  dff DFF_454(CK,G22955,G3994);
  dff DFF_455(CK,G22956,G3995);
  dff DFF_456(CK,G22957,G3996);
  dff DFF_457(CK,G22958,G3997);
  dff DFF_458(CK,G22959,G3998);
  dff DFF_459(CK,G22960,G3999);
  dff DFF_460(CK,G22961,G4000);
  dff DFF_461(CK,G22962,G4001);
  dff DFF_462(CK,G22963,G4002);
  dff DFF_463(CK,G22964,G4003);
  dff DFF_464(CK,G22965,G4004);
  dff DFF_465(CK,G22966,G4005);
  dff DFF_466(CK,G22967,G4006);
  dff DFF_467(CK,G22968,G4007);
  dff DFF_468(CK,G22969,G4008);
  dff DFF_469(CK,G22970,G4009);
  dff DFF_470(CK,G22971,G4010);
  dff DFF_471(CK,G22972,G4011);
  dff DFF_472(CK,G22973,G4012);
  dff DFF_473(CK,G22974,G4013);
  dff DFF_474(CK,G22975,G4014);
  dff DFF_475(CK,G22976,G4015);
  dff DFF_476(CK,G22977,G4016);
  dff DFF_477(CK,G22978,G4017);
  dff DFF_478(CK,G22979,G4018);
  dff DFF_479(CK,G22980,G4019);
  dff DFF_480(CK,G22981,G4229);
  dff DFF_481(CK,G22982,G4228);
  dff DFF_482(CK,G22983,G4227);
  dff DFF_483(CK,G22984,G4226);
  dff DFF_484(CK,G22985,G4225);
  dff DFF_485(CK,G22986,G4224);
  dff DFF_486(CK,G22987,G4223);
  dff DFF_487(CK,G22988,G4222);
  dff DFF_488(CK,G22989,G4221);
  dff DFF_489(CK,G22990,G4220);
  dff DFF_490(CK,G22991,G4219);
  dff DFF_491(CK,G22992,G4218);
  dff DFF_492(CK,G22993,G4217);
  dff DFF_493(CK,G22994,G4216);
  dff DFF_494(CK,G22995,G4215);
  dff DFF_495(CK,G22996,G4214);
  dff DFF_496(CK,G22997,G4213);
  dff DFF_497(CK,G22998,G4212);
  dff DFF_498(CK,G22999,G4211);
  dff DFF_499(CK,G23000,G4210);
  dff DFF_500(CK,G23001,G4209);
  dff DFF_501(CK,G23002,G4208);
  dff DFF_502(CK,G23003,G4207);
  dff DFF_503(CK,G23004,G4206);
  dff DFF_504(CK,G23005,G4205);
  dff DFF_505(CK,G23006,G4204);
  dff DFF_506(CK,G23007,G4203);
  dff DFF_507(CK,G23008,G4202);
  dff DFF_508(CK,G23009,G4201);
  dff DFF_509(CK,G23010,G4200);
  dff DFF_510(CK,G23011,G4199);
  dff DFF_511(CK,G23012,G4198);
  dff DFF_512(CK,G23013,G4020);
  dff DFF_513(CK,G23014,G4021);
  dff DFF_514(CK,G23015,G4022);
  dff DFF_515(CK,G23016,G4023);
  dff DFF_516(CK,G23017,G4024);
  dff DFF_517(CK,G23018,G4025);
  dff DFF_518(CK,G23019,G4026);
  dff DFF_519(CK,G23020,G4027);
  dff DFF_520(CK,G23021,G4028);
  dff DFF_521(CK,G23022,G4029);
  dff DFF_522(CK,G23023,G4030);
  dff DFF_523(CK,G23024,G4031);
  dff DFF_524(CK,G23025,G4032);
  dff DFF_525(CK,G23026,G4033);
  dff DFF_526(CK,G23027,G4034);
  dff DFF_527(CK,G23028,G4035);
  dff DFF_528(CK,G23029,G4036);
  dff DFF_529(CK,G23030,G4037);
  dff DFF_530(CK,G23031,G4038);
  dff DFF_531(CK,G23032,G4039);
  dff DFF_532(CK,G23033,G4040);
  dff DFF_533(CK,G23034,G4041);
  dff DFF_534(CK,G23035,G4042);
  dff DFF_535(CK,G23036,G4043);
  dff DFF_536(CK,G23037,G4044);
  dff DFF_537(CK,G23038,G4045);
  dff DFF_538(CK,G23039,G4046);
  dff DFF_539(CK,G23040,G4047);
  dff DFF_540(CK,G23041,G4048);
  dff DFF_541(CK,G23042,G4049);
  dff DFF_542(CK,G23043,G3841);
  dff DFF_543(CK,G23044,G3840);
  dff DFF_544(CK,G23045,G4365);
  not GNAME545(G545,G3681);
  and GNAME546(G546,G545,G3683);
  nand GNAME547(G547,G656,G657);
  nand GNAME548(G548,G658,G659);
  nand GNAME549(G549,G660,G661);
  nand GNAME550(G550,G662,G663);
  nand GNAME551(G551,G664,G665);
  nand GNAME552(G552,G666,G667);
  nand GNAME553(G553,G668,G669);
  nand GNAME554(G554,G670,G671);
  nand GNAME555(G555,G672,G673);
  nand GNAME556(G556,G674,G675);
  nand GNAME557(G557,G676,G677);
  nand GNAME558(G558,G678,G679);
  nand GNAME559(G559,G680,G681);
  nand GNAME560(G560,G682,G683);
  nand GNAME561(G561,G684,G685);
  nand GNAME562(G562,G686,G687);
  nand GNAME563(G563,G688,G689);
  nand GNAME564(G564,G690,G691);
  nand GNAME565(G565,G692,G693);
  nand GNAME566(G566,G694,G695);
  nand GNAME567(G567,G696,G697);
  nand GNAME568(G568,G698,G699);
  nand GNAME569(G569,G700,G701);
  nand GNAME570(G570,G702,G703);
  nand GNAME571(G571,G704,G705);
  nand GNAME572(G572,G706,G707);
  nand GNAME573(G573,G708,G709);
  nand GNAME574(G574,G710,G711);
  nand GNAME575(G575,G712,G713);
  nand GNAME576(G576,G714,G715);
  nand GNAME577(G577,G716,G717);
  nand GNAME578(G578,G718,G719);
  nand GNAME579(G579,G720,G721);
  nand GNAME580(G580,G722,G723);
  nand GNAME581(G581,G724,G725);
  nand GNAME582(G582,G726,G727);
  nand GNAME583(G583,G728,G729);
  nand GNAME584(G584,G730,G731);
  nand GNAME585(G585,G732,G733);
  nand GNAME586(G586,G734,G735);
  nand GNAME587(G587,G736,G737);
  nand GNAME588(G588,G738,G739);
  nand GNAME589(G589,G740,G741);
  nand GNAME590(G590,G742,G743);
  nand GNAME591(G591,G744,G745);
  nand GNAME592(G592,G746,G747);
  nand GNAME593(G593,G748,G749);
  nand GNAME594(G594,G750,G751);
  nand GNAME595(G595,G752,G753);
  nand GNAME596(G596,G754,G755);
  nand GNAME597(G597,G756,G757);
  nand GNAME598(G598,G758,G759);
  nand GNAME599(G599,G760,G761);
  nand GNAME600(G600,G762,G763);
  nand GNAME601(G601,G764,G765);
  nand GNAME602(G602,G766,G767);
  nand GNAME603(G603,G768,G769);
  nand GNAME604(G604,G770,G771);
  nand GNAME605(G605,G772,G773);
  nand GNAME606(G606,G774,G775);
  nand GNAME607(G607,G776,G777);
  nand GNAME608(G608,G778,G779);
  nand GNAME609(G609,G780,G781);
  nand GNAME610(G610,G782,G783);
  nand GNAME611(G611,G784,G785);
  nand GNAME612(G612,G786,G787);
  nand GNAME613(G613,G788,G789);
  nand GNAME614(G614,G790,G791);
  nand GNAME615(G615,G792,G793);
  nand GNAME616(G616,G794,G795);
  nand GNAME617(G617,G796,G797);
  nand GNAME618(G618,G798,G799);
  nand GNAME619(G619,G800,G801);
  nand GNAME620(G620,G802,G803);
  nand GNAME621(G621,G804,G805);
  nand GNAME622(G622,G806,G807);
  nand GNAME623(G623,G808,G809);
  nand GNAME624(G624,G810,G811);
  nand GNAME625(G625,G812,G813);
  nand GNAME626(G626,G814,G815);
  nand GNAME627(G627,G816,G817);
  nand GNAME628(G628,G818,G819);
  nand GNAME629(G629,G820,G821);
  nand GNAME630(G630,G822,G823);
  nand GNAME631(G631,G824,G825);
  nand GNAME632(G632,G826,G827);
  nand GNAME633(G633,G828,G829);
  nand GNAME634(G634,G830,G831);
  nand GNAME635(G635,G832,G833);
  nand GNAME636(G636,G834,G835);
  nand GNAME637(G637,G836,G837);
  nand GNAME638(G638,G838,G839);
  nand GNAME639(G639,G840,G841);
  nand GNAME640(G640,G842,G843);
  nand GNAME641(G641,G844,G845);
  nand GNAME642(G642,G846,G847);
  not GNAME643(G643,G23045);
  and GNAME644(G644,G652,G653);
  not GNAME645(G645,G22799);
  not GNAME646(G646,G23044);
  and GNAME647(G647,G654,G655);
  and GNAME648(G648,G649,G650);
  nand GNAME649(G649,G22716,G646,G22961);
  nand GNAME650(G650,G6757,G645,G6972);
  not GNAME651(G651,G648);
  nand GNAME652(G652,G643,G22800);
  or GNAME653(G653,G22800,G643);
  or GNAME654(G654,G23044,G645);
  or GNAME655(G655,G22799,G646);
  nand GNAME656(G656,G651,G22745);
  nand GNAME657(G657,G648,G6464);
  nand GNAME658(G658,G651,G22744);
  nand GNAME659(G659,G648,G6465);
  nand GNAME660(G660,G651,G22743);
  nand GNAME661(G661,G648,G6466);
  nand GNAME662(G662,G651,G22742);
  nand GNAME663(G663,G648,G6467);
  nand GNAME664(G664,G651,G22741);
  nand GNAME665(G665,G648,G6468);
  nand GNAME666(G666,G651,G22740);
  nand GNAME667(G667,G648,G6469);
  nand GNAME668(G668,G651,G22739);
  nand GNAME669(G669,G648,G6470);
  nand GNAME670(G670,G651,G22767);
  nand GNAME671(G671,G648,G6404);
  nand GNAME672(G672,G651,G22766);
  nand GNAME673(G673,G648,G6471);
  nand GNAME674(G674,G651,G22738);
  nand GNAME675(G675,G648,G6472);
  nand GNAME676(G676,G651,G22765);
  nand GNAME677(G677,G648,G6473);
  nand GNAME678(G678,G651,G22764);
  nand GNAME679(G679,G648,G6474);
  nand GNAME680(G680,G651,G22763);
  nand GNAME681(G681,G648,G6403);
  nand GNAME682(G682,G651,G22762);
  nand GNAME683(G683,G648,G6475);
  nand GNAME684(G684,G651,G22761);
  nand GNAME685(G685,G648,G6476);
  nand GNAME686(G686,G651,G22760);
  nand GNAME687(G687,G648,G6477);
  nand GNAME688(G688,G651,G22759);
  nand GNAME689(G689,G648,G6478);
  nand GNAME690(G690,G651,G22758);
  nand GNAME691(G691,G648,G6479);
  nand GNAME692(G692,G651,G22757);
  nand GNAME693(G693,G648,G6480);
  nand GNAME694(G694,G651,G22756);
  nand GNAME695(G695,G648,G6481);
  nand GNAME696(G696,G651,G22737);
  nand GNAME697(G697,G648,G6405);
  nand GNAME698(G698,G651,G22755);
  nand GNAME699(G699,G648,G6482);
  nand GNAME700(G700,G651,G22754);
  nand GNAME701(G701,G648,G6483);
  nand GNAME702(G702,G651,G22753);
  nand GNAME703(G703,G648,G6484);
  nand GNAME704(G704,G651,G22752);
  nand GNAME705(G705,G648,G6485);
  nand GNAME706(G706,G651,G22751);
  nand GNAME707(G707,G648,G6402);
  nand GNAME708(G708,G651,G22750);
  nand GNAME709(G709,G648,G6401);
  nand GNAME710(G710,G651,G22749);
  nand GNAME711(G711,G648,G6486);
  nand GNAME712(G712,G651,G22748);
  nand GNAME713(G713,G648,G6487);
  nand GNAME714(G714,G651,G22747);
  nand GNAME715(G715,G648,G6400);
  nand GNAME716(G716,G651,G22746);
  nand GNAME717(G717,G648,G6399);
  nand GNAME718(G718,G651,G22736);
  nand GNAME719(G719,G648,G6463);
  nand GNAME720(G720,G651,G6464);
  nand GNAME721(G721,G648,G22990);
  nand GNAME722(G722,G651,G6465);
  nand GNAME723(G723,G648,G22989);
  nand GNAME724(G724,G651,G6466);
  nand GNAME725(G725,G648,G22988);
  nand GNAME726(G726,G651,G6467);
  nand GNAME727(G727,G648,G22987);
  nand GNAME728(G728,G651,G6468);
  nand GNAME729(G729,G648,G22986);
  nand GNAME730(G730,G651,G6469);
  nand GNAME731(G731,G648,G22985);
  nand GNAME732(G732,G651,G6470);
  nand GNAME733(G733,G648,G22984);
  nand GNAME734(G734,G651,G6404);
  nand GNAME735(G735,G648,G23012);
  nand GNAME736(G736,G651,G6471);
  nand GNAME737(G737,G648,G23011);
  nand GNAME738(G738,G651,G6472);
  nand GNAME739(G739,G648,G22983);
  nand GNAME740(G740,G651,G6473);
  nand GNAME741(G741,G648,G23010);
  nand GNAME742(G742,G651,G6474);
  nand GNAME743(G743,G648,G23009);
  nand GNAME744(G744,G651,G6403);
  nand GNAME745(G745,G648,G23008);
  nand GNAME746(G746,G651,G6475);
  nand GNAME747(G747,G648,G23007);
  nand GNAME748(G748,G651,G6476);
  nand GNAME749(G749,G648,G23006);
  nand GNAME750(G750,G651,G6477);
  nand GNAME751(G751,G648,G23005);
  nand GNAME752(G752,G651,G6478);
  nand GNAME753(G753,G648,G23004);
  nand GNAME754(G754,G651,G6479);
  nand GNAME755(G755,G648,G23003);
  nand GNAME756(G756,G651,G6480);
  nand GNAME757(G757,G648,G23002);
  nand GNAME758(G758,G651,G6481);
  nand GNAME759(G759,G648,G23001);
  nand GNAME760(G760,G651,G6405);
  nand GNAME761(G761,G648,G22982);
  nand GNAME762(G762,G651,G6482);
  nand GNAME763(G763,G648,G23000);
  nand GNAME764(G764,G651,G6483);
  nand GNAME765(G765,G648,G22999);
  nand GNAME766(G766,G651,G6484);
  nand GNAME767(G767,G648,G22998);
  nand GNAME768(G768,G651,G6485);
  nand GNAME769(G769,G648,G22997);
  nand GNAME770(G770,G651,G6402);
  nand GNAME771(G771,G648,G22996);
  nand GNAME772(G772,G651,G6401);
  nand GNAME773(G773,G648,G22995);
  nand GNAME774(G774,G651,G6486);
  nand GNAME775(G775,G648,G22994);
  nand GNAME776(G776,G651,G6487);
  nand GNAME777(G777,G648,G22993);
  nand GNAME778(G778,G651,G6400);
  nand GNAME779(G779,G648,G22992);
  nand GNAME780(G780,G651,G6399);
  nand GNAME781(G781,G648,G22991);
  nand GNAME782(G782,G651,G6463);
  nand GNAME783(G783,G648,G22981);
  nand GNAME784(G784,G651,G22990);
  nand GNAME785(G785,G22745,G648);
  nand GNAME786(G786,G651,G22989);
  nand GNAME787(G787,G648,G22744);
  nand GNAME788(G788,G651,G22988);
  nand GNAME789(G789,G648,G22743);
  nand GNAME790(G790,G651,G22987);
  nand GNAME791(G791,G648,G22742);
  nand GNAME792(G792,G651,G22986);
  nand GNAME793(G793,G648,G22741);
  nand GNAME794(G794,G651,G22985);
  nand GNAME795(G795,G648,G22740);
  nand GNAME796(G796,G651,G23012);
  nand GNAME797(G797,G648,G22767);
  nand GNAME798(G798,G651,G23011);
  nand GNAME799(G799,G648,G22766);
  nand GNAME800(G800,G651,G22984);
  nand GNAME801(G801,G648,G22739);
  nand GNAME802(G802,G651,G23010);
  nand GNAME803(G803,G648,G22765);
  nand GNAME804(G804,G651,G23009);
  nand GNAME805(G805,G648,G22764);
  nand GNAME806(G806,G651,G23008);
  nand GNAME807(G807,G648,G22763);
  nand GNAME808(G808,G651,G23007);
  nand GNAME809(G809,G648,G22762);
  nand GNAME810(G810,G651,G23006);
  nand GNAME811(G811,G648,G22761);
  nand GNAME812(G812,G651,G23005);
  nand GNAME813(G813,G648,G22760);
  nand GNAME814(G814,G651,G23004);
  nand GNAME815(G815,G648,G22759);
  nand GNAME816(G816,G651,G23003);
  nand GNAME817(G817,G648,G22758);
  nand GNAME818(G818,G651,G23002);
  nand GNAME819(G819,G648,G22757);
  nand GNAME820(G820,G651,G23001);
  nand GNAME821(G821,G648,G22756);
  nand GNAME822(G822,G651,G22983);
  nand GNAME823(G823,G648,G22738);
  nand GNAME824(G824,G651,G23000);
  nand GNAME825(G825,G648,G22755);
  nand GNAME826(G826,G651,G22999);
  nand GNAME827(G827,G648,G22754);
  nand GNAME828(G828,G651,G22998);
  nand GNAME829(G829,G648,G22753);
  nand GNAME830(G830,G651,G22997);
  nand GNAME831(G831,G648,G22752);
  nand GNAME832(G832,G651,G22996);
  nand GNAME833(G833,G648,G22751);
  nand GNAME834(G834,G651,G22995);
  nand GNAME835(G835,G648,G22750);
  nand GNAME836(G836,G651,G22994);
  nand GNAME837(G837,G648,G22749);
  nand GNAME838(G838,G651,G22993);
  nand GNAME839(G839,G648,G22748);
  nand GNAME840(G840,G651,G22992);
  nand GNAME841(G841,G648,G22747);
  nand GNAME842(G842,G651,G22991);
  nand GNAME843(G843,G648,G22746);
  nand GNAME844(G844,G651,G22982);
  nand GNAME845(G845,G648,G22737);
  nand GNAME846(G846,G651,G22981);
  nand GNAME847(G847,G648,G22736);
  nand GNAME848(G848,G6339,G4238);
  nand GNAME849(G849,G850,G852,G851);
  nand GNAME850(G850,G6340,G4239);
  or GNAME851(G851,G4238,G6339);
  nand GNAME852(G852,G853,G855,G854);
  nand GNAME853(G853,G6341,G4102);
  or GNAME854(G854,G4239,G6340);
  nand GNAME855(G855,G856,G858,G857);
  nand GNAME856(G856,G6342,G4242);
  or GNAME857(G857,G4102,G6341);
  nand GNAME858(G858,G859,G861,G860);
  nand GNAME859(G859,G6343,G4092);
  or GNAME860(G860,G4242,G6342);
  nand GNAME861(G861,G862,G864,G863);
  nand GNAME862(G862,G6344,G4244);
  or GNAME863(G863,G4092,G6343);
  nand GNAME864(G864,G865,G867,G866);
  nand GNAME865(G865,G6345,G4096);
  or GNAME866(G866,G4244,G6344);
  nand GNAME867(G867,G868,G3609,G3608);
  nand GNAME868(G868,G6346,G4246);
  or GNAME869(G869,G1333,G3062);
  or GNAME870(G870,G871,G3062);
  nand GNAME871(G871,G2997,G2998,G2996,G2994,G2995);
  nand GNAME872(G872,G3003,G2994,G3002);
  nand GNAME873(G873,G3005,G2994,G3004);
  nand GNAME874(G874,G3007,G2994,G3006);
  nand GNAME875(G875,G3009,G2994,G3008);
  nand GNAME876(G876,G3011,G2994,G3010);
  nand GNAME877(G877,G3013,G2994,G3012);
  nand GNAME878(G878,G3015,G2994,G3014);
  nand GNAME879(G879,G3017,G2994,G3016);
  nand GNAME880(G880,G3019,G2994,G3018);
  nand GNAME881(G881,G3024,G2994,G3023);
  nand GNAME882(G882,G3027,G3025,G3026);
  nand GNAME883(G883,G3030,G3028,G3029);
  nand GNAME884(G884,G3033,G3031,G3032);
  nand GNAME885(G885,G3036,G3034,G3035);
  nand GNAME886(G886,G3039,G3037,G3038);
  nand GNAME887(G887,G3042,G3040,G3041);
  nand GNAME888(G888,G3045,G3043,G3044);
  nand GNAME889(G889,G3048,G3046,G3047);
  nand GNAME890(G890,G3051,G3049,G3050);
  nand GNAME891(G891,G2978,G2976,G2977);
  nand GNAME892(G892,G2981,G2979,G2980);
  nand GNAME893(G893,G2984,G2982,G2983);
  nand GNAME894(G894,G2987,G2985,G2986);
  nand GNAME895(G895,G2990,G2988,G2989);
  nand GNAME896(G896,G2993,G2991,G2992);
  nand GNAME897(G897,G3001,G2999,G3000);
  nand GNAME898(G898,G3022,G3020,G3021);
  nand GNAME899(G899,G3054,G3052,G3053);
  nand GNAME900(G900,G3055,G3056,G3057,G3058);
  nand GNAME901(G901,G2899,G1340);
  nand GNAME902(G902,G1668,G1666,G1667);
  nand GNAME903(G903,G2900,G1340);
  nand GNAME904(G904,G1671,G1669,G1670);
  nand GNAME905(G905,G2905,G1340);
  nand GNAME906(G906,G1339,G2906,G2907);
  nand GNAME907(G907,G1339,G2908,G2909);
  nand GNAME908(G908,G1339,G2910,G2911);
  nand GNAME909(G909,G1339,G2912,G2913);
  nand GNAME910(G910,G1339,G2914,G2915);
  nand GNAME911(G911,G1339,G2916,G2917);
  nand GNAME912(G912,G1339,G2918,G2919);
  nand GNAME913(G913,G1339,G2920,G2921);
  nand GNAME914(G914,G1339,G2922,G2923);
  nand GNAME915(G915,G1339,G2928,G2929);
  nand GNAME916(G916,G2930,G2931,G2932,G2933);
  nand GNAME917(G917,G2934,G2935,G2936,G2937);
  nand GNAME918(G918,G2938,G2939,G2940,G2941);
  nand GNAME919(G919,G2942,G2943,G2944,G2945);
  nand GNAME920(G920,G2946,G2947,G2948,G2949);
  nand GNAME921(G921,G2950,G2951,G2952,G2953);
  nand GNAME922(G922,G2954,G2955,G2956,G2957);
  nand GNAME923(G923,G2958,G2959,G2960,G2961);
  nand GNAME924(G924,G2962,G2963,G2964,G2965);
  nand GNAME925(G925,G2869,G2870,G2871,G2872);
  nand GNAME926(G926,G2873,G2874,G2875,G2876);
  nand GNAME927(G927,G2877,G2878,G2879,G2880);
  nand GNAME928(G928,G2881,G2882,G2883,G2884);
  nand GNAME929(G929,G2885,G2886,G2887,G2888);
  nand GNAME930(G930,G2889,G2890,G2891,G2892);
  nand GNAME931(G931,G2901,G2902,G2903,G2904);
  nand GNAME932(G932,G2924,G2925,G2926,G2927);
  nand GNAME933(G933,G2966,G2967,G2968,G2969);
  nand GNAME934(G934,G2973,G2974,G2972,G2970,G2971);
  nand GNAME935(G935,G1215,G1216);
  nand GNAME936(G936,G1629,G1322,G3062,G3561,G3562);
  nand GNAME937(G937,G2766,G2764,G2765);
  nand GNAME938(G938,G2769,G2767,G2768);
  nand GNAME939(G939,G2773,G2774,G2775,G1324);
  nand GNAME940(G940,G2776,G2777,G2778,G1324);
  nand GNAME941(G941,G2779,G2780,G2781,G1324);
  nand GNAME942(G942,G2782,G2783,G2784,G1324);
  nand GNAME943(G943,G2785,G2786,G2787,G1324);
  nand GNAME944(G944,G2788,G2789,G2790,G1324);
  nand GNAME945(G945,G2791,G2792,G2793,G1324);
  nand GNAME946(G946,G2794,G2795,G2796,G1324);
  nand GNAME947(G947,G2797,G2798,G2799,G1324);
  nand GNAME948(G948,G2800,G2801,G2802,G1324);
  nand GNAME949(G949,G2806,G2807,G2808,G1324);
  nand GNAME950(G950,G2809,G2810,G2811,G1324);
  nand GNAME951(G951,G2812,G2813,G2814,G1324);
  nand GNAME952(G952,G2815,G2816,G2817,G1324);
  nand GNAME953(G953,G2818,G2819,G2820,G1324);
  nand GNAME954(G954,G2821,G2822,G2823,G1324);
  nand GNAME955(G955,G2824,G2825,G2826,G1324);
  nand GNAME956(G956,G2827,G2828,G2829,G1324);
  nand GNAME957(G957,G2830,G2831,G2832,G1324);
  nand GNAME958(G958,G2833,G2834,G2835,G1324);
  nand GNAME959(G959,G2746,G2747,G2748,G1324);
  nand GNAME960(G960,G2749,G2750,G2751,G1324);
  nand GNAME961(G961,G2752,G2753,G2754,G1324);
  nand GNAME962(G962,G2755,G2756,G2757,G1324);
  nand GNAME963(G963,G2758,G2759,G2760,G1324);
  nand GNAME964(G964,G2761,G2762,G2763,G1324);
  nand GNAME965(G965,G2770,G2771,G2772,G1324);
  nand GNAME966(G966,G2803,G2804,G2805,G1324);
  nand GNAME967(G967,G2836,G2837,G2838,G1324);
  nand GNAME968(G968,G2839,G2840,G2841,G1324);
  nand GNAME969(G969,G2643,G2641,G2642);
  nand GNAME970(G970,G2646,G2644,G2645);
  nand GNAME971(G971,G2651,G2652,G2653,G2654);
  nand GNAME972(G972,G2655,G2656,G2657,G2658);
  nand GNAME973(G973,G2659,G2660,G2661,G2662);
  nand GNAME974(G974,G2663,G2664,G2665,G2666);
  nand GNAME975(G975,G2667,G2668,G2669,G2670);
  nand GNAME976(G976,G2671,G2672,G2673,G2674);
  nand GNAME977(G977,G2675,G2676,G2677,G2678);
  nand GNAME978(G978,G2679,G2680,G2681,G2682);
  nand GNAME979(G979,G2683,G2684,G2685,G2686);
  nand GNAME980(G980,G2687,G2688,G2689,G2690);
  nand GNAME981(G981,G2695,G2696,G2697,G2698);
  nand GNAME982(G982,G2699,G2700,G2701,G2702);
  nand GNAME983(G983,G2703,G2704,G2705,G2706);
  nand GNAME984(G984,G2707,G2708,G2709,G2710);
  nand GNAME985(G985,G2711,G2712,G2713,G2714);
  nand GNAME986(G986,G2715,G2716,G2717,G2718);
  nand GNAME987(G987,G2719,G2720,G2721,G2722);
  nand GNAME988(G988,G2723,G2724,G2725,G2726);
  nand GNAME989(G989,G2727,G2728,G2729,G2730);
  nand GNAME990(G990,G2731,G2732,G2733,G2734);
  nand GNAME991(G991,G2617,G2618,G2619,G2620);
  nand GNAME992(G992,G2621,G2622,G2623,G2624);
  nand GNAME993(G993,G2625,G2626,G2627,G2628);
  nand GNAME994(G994,G2629,G2630,G2631,G2632);
  nand GNAME995(G995,G2633,G2634,G2635,G2636);
  nand GNAME996(G996,G2637,G2638,G2639,G2640);
  nand GNAME997(G997,G2647,G2648,G2649,G2650);
  nand GNAME998(G998,G2691,G2692,G2693,G2694);
  nand GNAME999(G999,G2735,G2736,G2737,G2738);
  nand GNAME1000(G1000,G2741,G2739,G2740);
  nand GNAME1001(G1001,G22798,G1637);
  nand GNAME1002(G1002,G2855,G1330);
  nand GNAME1003(G1003,G1330,G2856,G1367);
  nand GNAME1004(G1004,G2857,G1330);
  and GNAME1005(G1005,G2851,G1245);
  and GNAME1006(G1006,G2851,G1243);
  and GNAME1007(G1007,G2851,G1251);
  and GNAME1008(G1008,G2851,G1247);
  and GNAME1009(G1009,G2851,G1248);
  and GNAME1010(G1010,G2851,G1244);
  and GNAME1011(G1011,G2851,G1250);
  and GNAME1012(G1012,G2851,G1246);
  and GNAME1013(G1013,G2851,G1249);
  and GNAME1014(G1014,G2851,G1409);
  and GNAME1015(G1015,G2851,G1422);
  and GNAME1016(G1016,G2851,G1415);
  and GNAME1017(G1017,G2851,G1413);
  and GNAME1018(G1018,G2851,G1424);
  and GNAME1019(G1019,G2851,G1406);
  and GNAME1020(G1020,G2851,G1419);
  and GNAME1021(G1021,G2851,G1412);
  and GNAME1022(G1022,G2851,G1420);
  and GNAME1023(G1023,G2851,G1407);
  and GNAME1024(G1024,G2851,G1417);
  and GNAME1025(G1025,G2851,G1410);
  and GNAME1026(G1026,G2851,G1405);
  and GNAME1027(G1027,G2851,G1423);
  and GNAME1028(G1028,G2851,G1414);
  and GNAME1029(G1029,G2851,G1416);
  and GNAME1030(G1030,G2851,G1408);
  and GNAME1031(G1031,G2851,G1421);
  and GNAME1032(G1032,G2851,G1411);
  and GNAME1033(G1033,G2851,G1418);
  nand GNAME1034(G1034,G2847,G1327);
  nand GNAME1035(G1035,G2848,G1327);
  nand GNAME1036(G1036,G2849,G1327);
  and GNAME1037(G1037,G1285,G2844);
  and GNAME1038(G1038,G1284,G2844);
  and GNAME1039(G1039,G1283,G2844);
  and GNAME1040(G1040,G1282,G2844);
  and GNAME1041(G1041,G1281,G2844);
  and GNAME1042(G1042,G1280,G2844);
  and GNAME1043(G1043,G1279,G2844);
  and GNAME1044(G1044,G1278,G2844);
  and GNAME1045(G1045,G1277,G2844);
  and GNAME1046(G1046,G1276,G2844);
  and GNAME1047(G1047,G1275,G2844);
  and GNAME1048(G1048,G1274,G2844);
  and GNAME1049(G1049,G1273,G2844);
  and GNAME1050(G1050,G1272,G2844);
  and GNAME1051(G1051,G1271,G2844);
  and GNAME1052(G1052,G1270,G2844);
  and GNAME1053(G1053,G1269,G2844);
  and GNAME1054(G1054,G1268,G2844);
  and GNAME1055(G1055,G1267,G2844);
  and GNAME1056(G1056,G1266,G2844);
  and GNAME1057(G1057,G1265,G2844);
  and GNAME1058(G1058,G1264,G2844);
  and GNAME1059(G1059,G1263,G2844);
  and GNAME1060(G1060,G1262,G2844);
  and GNAME1061(G1061,G1261,G2844);
  and GNAME1062(G1062,G1260,G2844);
  and GNAME1063(G1063,G1259,G2844);
  and GNAME1064(G1064,G1258,G2844);
  and GNAME1065(G1065,G1257,G2844);
  not GNAME1066(G1066,G22798);
  nand GNAME1067(G1067,G2609,G2607,G2608);
  nand GNAME1068(G1068,G2606,G2604,G2605);
  nand GNAME1069(G1069,G2603,G2601,G2602);
  nand GNAME1070(G1070,G2600,G2598,G2599);
  nand GNAME1071(G1071,G2597,G2595,G2596);
  nand GNAME1072(G1072,G2594,G2592,G2593);
  nand GNAME1073(G1073,G2591,G2589,G2590);
  nand GNAME1074(G1074,G2588,G2586,G2587);
  nand GNAME1075(G1075,G2585,G2583,G2584);
  nand GNAME1076(G1076,G2582,G2580,G2581);
  nand GNAME1077(G1077,G2579,G2577,G2578);
  nand GNAME1078(G1078,G2576,G2574,G2575);
  nand GNAME1079(G1079,G2573,G2571,G2572);
  nand GNAME1080(G1080,G2570,G2568,G2569);
  nand GNAME1081(G1081,G2567,G2565,G2566);
  nand GNAME1082(G1082,G2564,G2562,G2563);
  nand GNAME1083(G1083,G2561,G2559,G2560);
  nand GNAME1084(G1084,G2558,G2556,G2557);
  nand GNAME1085(G1085,G2555,G2553,G2554);
  nand GNAME1086(G1086,G2552,G2550,G2551);
  nand GNAME1087(G1087,G2549,G2547,G2548);
  nand GNAME1088(G1088,G2546,G2544,G2545);
  nand GNAME1089(G1089,G2543,G2541,G2542);
  nand GNAME1090(G1090,G2540,G2538,G2539);
  nand GNAME1091(G1091,G2537,G2535,G2536);
  nand GNAME1092(G1092,G2534,G2532,G2533);
  nand GNAME1093(G1093,G2531,G2529,G2530);
  nand GNAME1094(G1094,G2528,G2526,G2527);
  nand GNAME1095(G1095,G2525,G2523,G2524);
  nand GNAME1096(G1096,G2522,G2520,G2521);
  nand GNAME1097(G1097,G2519,G2517,G2518);
  nand GNAME1098(G1098,G2516,G2514,G2515);
  and GNAME1099(G1099,G2513,G22590);
  and GNAME1100(G1100,G2513,G22591);
  and GNAME1101(G1101,G2513,G22592);
  and GNAME1102(G1102,G2513,G22593);
  and GNAME1103(G1103,G2513,G22594);
  and GNAME1104(G1104,G2513,G22595);
  and GNAME1105(G1105,G2513,G22596);
  and GNAME1106(G1106,G2513,G22597);
  and GNAME1107(G1107,G2513,G22598);
  and GNAME1108(G1108,G2513,G22599);
  and GNAME1109(G1109,G2513,G22600);
  and GNAME1110(G1110,G2513,G22601);
  and GNAME1111(G1111,G2513,G22602);
  and GNAME1112(G1112,G2513,G22603);
  and GNAME1113(G1113,G2513,G22604);
  and GNAME1114(G1114,G2513,G22605);
  and GNAME1115(G1115,G2513,G22606);
  and GNAME1116(G1116,G2513,G22607);
  and GNAME1117(G1117,G2513,G22608);
  and GNAME1118(G1118,G2513,G22609);
  and GNAME1119(G1119,G2513,G22610);
  and GNAME1120(G1120,G2513,G22611);
  and GNAME1121(G1121,G2513,G22612);
  and GNAME1122(G1122,G2513,G22613);
  and GNAME1123(G1123,G2513,G22614);
  and GNAME1124(G1124,G2513,G22615);
  and GNAME1125(G1125,G2513,G22616);
  and GNAME1126(G1126,G2513,G22617);
  and GNAME1127(G1127,G2513,G22618);
  and GNAME1128(G1128,G2513,G22619);
  nand GNAME1129(G1129,G1620,G2321,G2319,G2320);
  nand GNAME1130(G1130,G1619,G2307,G2305,G2306);
  nand GNAME1131(G1131,G1618,G2300,G2298,G2299);
  nand GNAME1132(G1132,G1617,G2293,G2291,G2292);
  nand GNAME1133(G1133,G1616,G2286,G2284,G2285);
  nand GNAME1134(G1134,G1615,G2279,G2277,G2278);
  nand GNAME1135(G1135,G1614,G2272,G2270,G2271);
  nand GNAME1136(G1136,G1613,G2265,G2263,G2264);
  nand GNAME1137(G1137,G1612,G2258,G2256,G2257);
  nand GNAME1138(G1138,G1611,G2251,G2249,G2250);
  nand GNAME1139(G1139,G1610,G2244,G2242,G2243);
  nand GNAME1140(G1140,G1609,G2237,G2235,G2236);
  nand GNAME1141(G1141,G1608,G2230,G2228,G2229);
  nand GNAME1142(G1142,G1607,G2223,G2221,G2222);
  nand GNAME1143(G1143,G1606,G2216,G2214,G2215);
  nand GNAME1144(G1144,G1605,G2209,G2207,G2208);
  nand GNAME1145(G1145,G1604,G2202,G2200,G2201);
  nand GNAME1146(G1146,G1603,G2195,G2193,G2194);
  nand GNAME1147(G1147,G1602,G2188,G2186,G2187);
  nand GNAME1148(G1148,G1601,G2181,G2179,G2180);
  nand GNAME1149(G1149,G1600,G2174,G2172,G2173);
  nand GNAME1150(G1150,G1599,G2167,G2165,G2166);
  nand GNAME1151(G1151,G1598,G2160,G2158,G2159);
  nand GNAME1152(G1152,G1597,G2153,G2151,G2152);
  nand GNAME1153(G1153,G1596,G2146,G2144,G2145);
  nand GNAME1154(G1154,G1595,G2139,G2137,G2138);
  nand GNAME1155(G1155,G1594,G2132,G2130,G2131);
  nand GNAME1156(G1156,G1593,G2125,G2123,G2124);
  nand GNAME1157(G1157,G2118,G1624,G2117,G2115,G2116);
  nand GNAME1158(G1158,G2107,G3421,G3422);
  nand GNAME1159(G1159,G2104,G3419,G3420);
  nand GNAME1160(G1160,G1592,G2097,G2095,G2096);
  nand GNAME1161(G1161,G2093,G2094,G2092,G2090,G2091);
  nand GNAME1162(G1162,G2088,G2089,G2087,G2085,G2086);
  nand GNAME1163(G1163,G2083,G2084,G2082,G2080,G2081);
  nand GNAME1164(G1164,G2078,G2079,G2077,G2075,G2076);
  nand GNAME1165(G1165,G2073,G2074,G2072,G2070,G2071);
  nand GNAME1166(G1166,G2068,G2069,G2067,G2065,G2066);
  nand GNAME1167(G1167,G2063,G2064,G2062,G2060,G2061);
  nand GNAME1168(G1168,G2058,G2059,G2057,G2055,G2056);
  nand GNAME1169(G1169,G2053,G2054,G2052,G2050,G2051);
  nand GNAME1170(G1170,G2048,G2049,G2047,G2045,G2046);
  nand GNAME1171(G1171,G2043,G2044,G2042,G2040,G2041);
  nand GNAME1172(G1172,G2038,G2039,G2037,G2035,G2036);
  nand GNAME1173(G1173,G2033,G2034,G2032,G2030,G2031);
  nand GNAME1174(G1174,G2028,G2029,G2027,G2025,G2026);
  nand GNAME1175(G1175,G1591,G2021,G2019,G2020);
  nand GNAME1176(G1176,G2017,G2018,G2016,G2014,G2015);
  nand GNAME1177(G1177,G1590,G2011,G2009,G2024);
  nand GNAME1178(G1178,G2007,G2008,G2006,G2004,G2005);
  nand GNAME1179(G1179,G2002,G2003,G2001,G1999,G2000);
  nand GNAME1180(G1180,G1991,G1989,G1990);
  nand GNAME1181(G1181,G1581,G1966,G1967,G1968,G1970);
  nand GNAME1182(G1182,G1580,G1959,G1960,G1961,G1964);
  nand GNAME1183(G1183,G1579,G1953,G1954,G1955,G1957);
  nand GNAME1184(G1184,G1578,G1947,G1948,G1949,G1951);
  nand GNAME1185(G1185,G1577,G1941,G1942,G1943,G1944);
  nand GNAME1186(G1186,G1576,G1935,G1936,G1937,G1939);
  nand GNAME1187(G1187,G1575,G1928,G1929,G1930,G1933);
  nand GNAME1188(G1188,G1574,G1922,G1923,G1924,G1926);
  nand GNAME1189(G1189,G1573,G1915,G1916,G1917,G1920);
  nand GNAME1190(G1190,G1572,G1912,G1910,G1911);
  nand GNAME1191(G1191,G1571,G1904,G1905,G1906,G1908);
  nand GNAME1192(G1192,G1570,G1898,G1899,G1900,G1901);
  nand GNAME1193(G1193,G1569,G1891,G1892,G1893,G1896);
  nand GNAME1194(G1194,G1568,G1885,G1886,G1887,G1889);
  nand GNAME1195(G1195,G1567,G1879,G1880,G1881,G1883);
  nand GNAME1196(G1196,G1566,G1873,G1874,G1875,G1877);
  nand GNAME1197(G1197,G1565,G1866,G1867,G1868,G1871);
  nand GNAME1198(G1198,G1564,G1860,G1861,G1862,G1864);
  nand GNAME1199(G1199,G1563,G1853,G1854,G1855,G1858);
  nand GNAME1200(G1200,G1562,G1847,G1848,G1849,G1850);
  nand GNAME1201(G1201,G1561,G1841,G1842,G1843,G1845);
  nand GNAME1202(G1202,G1560,G1834,G1835,G1836,G1839);
  nand GNAME1203(G1203,G1559,G1828,G1829,G1830,G1832);
  nand GNAME1204(G1204,G1558,G1822,G1823,G1824,G1825);
  nand GNAME1205(G1205,G1557,G1816,G1817,G1818,G1820);
  nand GNAME1206(G1206,G1556,G1809,G1810,G1811,G1814);
  nand GNAME1207(G1207,G1555,G1803,G1804,G1805,G1807);
  nand GNAME1208(G1208,G1554,G1796,G1797,G1798,G1801);
  nand GNAME1209(G1209,G1553,G1790,G1791,G1792,G1794);
  nor GNAME1210(G1210,G1345,G1343,G1344);
  nor GNAME1211(G1211,G3062,G1634);
  not GNAME1212(G1212,G7865);
  not GNAME1213(G1213,G22585);
  not GNAME1214(G1214,G7897);
  nor GNAME1215(G1215,G3062,G1368);
  nor GNAME1216(G1216,G3197,G1367,G3200);
  nor GNAME1217(G1217,G1766,G1343);
  and GNAME1218(G1218,G3206,G3209);
  and GNAME1219(G1219,G1769,G1770);
  and GNAME1220(G1220,G1218,G1219);
  nor GNAME1221(G1221,G1210,G935,G1066);
  and GNAME1222(G1222,G1221,G3112,G1220);
  and GNAME1223(G1223,G1221,G1220,G1366);
  and GNAME1224(G1224,G3200,G1368);
  nor GNAME1225(G1225,G3200,G3118);
  nor GNAME1226(G1226,G1368,G1403);
  nand GNAME1227(G1227,G1367,G1225);
  nor GNAME1228(G1228,G3200,G1368);
  nand GNAME1229(G1229,G1404,G1228);
  nor GNAME1230(G1230,G1403,G3197);
  nand GNAME1231(G1231,G3197,G1228);
  and GNAME1232(G1232,G1774,G1775);
  nand GNAME1233(G1233,G1232,G1778,G2862);
  nand GNAME1234(G1234,G1765,G1764);
  nor GNAME1235(G1235,G1367,G1368);
  and GNAME1236(G1236,G1342,G22798,G1634);
  and GNAME1237(G1237,G1220,G1236);
  and GNAME1238(G1238,G1233,G1237);
  and GNAME1239(G1239,G1234,G1237);
  and GNAME1240(G1240,G1779,G3197);
  nand GNAME1241(G1241,G1367,G1224);
  nor GNAME1242(G1242,G3197,G1241);
  and GNAME1243(G1243,G1632,G591);
  and GNAME1244(G1244,G1632,G595);
  and GNAME1245(G1245,G1632,G590);
  and GNAME1246(G1246,G1632,G597);
  and GNAME1247(G1247,G1632,G593);
  and GNAME1248(G1248,G1632,G594);
  and GNAME1249(G1249,G1632,G598);
  and GNAME1250(G1250,G1632,G596);
  and GNAME1251(G1251,G1632,G592);
  nor GNAME1252(G1252,G1366,G1365,G1368,G3605);
  and GNAME1253(G1253,G1632,G589);
  nand GNAME1254(G1254,G1676,G1677,G1678,G1679);
  and GNAME1255(G1255,G1632,G586);
  and GNAME1256(G1256,G1632,G587);
  nand GNAME1257(G1257,G1760,G1761,G1762,G1763);
  nand GNAME1258(G1258,G1716,G1717,G1718,G1719);
  nand GNAME1259(G1259,G1672,G1673,G1674,G1675);
  nand GNAME1260(G1260,G1662,G1663,G1664,G1665);
  nand GNAME1261(G1261,G1658,G1659,G1660,G1661);
  nand GNAME1262(G1262,G1654,G1655,G1656,G1657);
  nand GNAME1263(G1263,G1650,G1651,G1652,G1653);
  nand GNAME1264(G1264,G1646,G1647,G1648,G1649);
  nand GNAME1265(G1265,G1642,G1643,G1644,G1645);
  nand GNAME1266(G1266,G1638,G1639,G1640,G1641);
  nand GNAME1267(G1267,G1756,G1757,G1758,G1759);
  nand GNAME1268(G1268,G1752,G1753,G1754,G1755);
  nand GNAME1269(G1269,G1748,G1749,G1750,G1751);
  nand GNAME1270(G1270,G1744,G1745,G1746,G1747);
  nand GNAME1271(G1271,G1740,G1741,G1742,G1743);
  nand GNAME1272(G1272,G1736,G1737,G1738,G1739);
  nand GNAME1273(G1273,G1732,G1733,G1734,G1735);
  nand GNAME1274(G1274,G1728,G1729,G1730,G1731);
  nand GNAME1275(G1275,G1724,G1725,G1726,G1727);
  nand GNAME1276(G1276,G1720,G1721,G1722,G1723);
  nand GNAME1277(G1277,G1712,G1713,G1714,G1715);
  nand GNAME1278(G1278,G1708,G1709,G1710,G1711);
  nand GNAME1279(G1279,G1704,G1705,G1706,G1707);
  nand GNAME1280(G1280,G1700,G1701,G1702,G1703);
  nand GNAME1281(G1281,G1696,G1697,G1698,G1699);
  nand GNAME1282(G1282,G1692,G1693,G1694,G1695);
  nand GNAME1283(G1283,G1688,G1689,G1690,G1691);
  nand GNAME1284(G1284,G1684,G1685,G1686,G1687);
  nand GNAME1285(G1285,G1680,G1681,G1682,G1683);
  nor GNAME1286(G1286,G1404,G3115);
  and GNAME1287(G1287,G3062,G3200);
  nor GNAME1288(G1288,G1367,G1404);
  and GNAME1289(G1289,G1583,G1585,G1587,G1589);
  nor GNAME1290(G1290,G1066,G1628);
  or GNAME1291(G1291,G1303,G1226);
  and GNAME1292(G1292,G1992,G1236);
  and GNAME1293(G1293,G1292,G1296,G3112);
  or GNAME1294(G1294,G1066,G1342);
  and GNAME1295(G1295,G1777,G1776);
  or GNAME1296(G1296,G1291,G1240,G1242);
  nand GNAME1297(G1297,G3605,G1231,G1229,G1295);
  and GNAME1298(G1298,G1995,G1366);
  and GNAME1299(G1299,G3112,G1994);
  nor GNAME1300(G1300,G1001,G1211);
  and GNAME1301(G1301,G2099,G1236);
  and GNAME1302(G1302,G1240,G1301);
  nor GNAME1303(G1303,G3197,G1227);
  and GNAME1304(G1304,G1232,G1231,G1776);
  and GNAME1305(G1305,G2109,G1301);
  and GNAME1306(G1306,G1291,G1301);
  and GNAME1307(G1307,G1242,G1301);
  and GNAME1308(G1308,G1366,G1235);
  and GNAME1309(G1309,G1301,G1308);
  and GNAME1310(G1310,G3112,G1235);
  and GNAME1311(G1311,G1301,G1310);
  and GNAME1312(G1312,G2308,G2309);
  and GNAME1313(G1313,G1236,G2323,G1219);
  nor GNAME1314(G1314,G3115,G3118,G3197);
  nor GNAME1315(G1315,G3206,G3209);
  nor GNAME1316(G1316,G1066,G22587);
  nor GNAME1317(G1317,G1066,G1316);
  and GNAME1318(G1318,G2615,G1241);
  and GNAME1319(G1319,G2611,G1227,G1777);
  nor GNAME1320(G1320,G1321,G3606);
  and GNAME1321(G1321,G1231,G2610);
  nand GNAME1322(G1322,G3197,G1225);
  nor GNAME1323(G1323,G3606,G1322);
  and GNAME1324(G1324,G2742,G3062);
  nor GNAME1325(G1325,G2843,G1326);
  and GNAME1326(G1326,G2842,G1328);
  and GNAME1327(G1327,G2845,G2846);
  or GNAME1328(G1328,G1230,G1286);
  and GNAME1329(G1329,G2842,G1403);
  and GNAME1330(G1330,G2854,G2853);
  nor GNAME1331(G1331,G1210,G1229);
  nand GNAME1332(G1332,G2866,G2867);
  nor GNAME1333(G1333,G1776,G1210,G3062);
  nand GNAME1334(G1334,G2858,G2859);
  or GNAME1335(G1335,G2860,G1334);
  and GNAME1336(G1336,G1365,G1634,G1296);
  and GNAME1337(G1337,G3109,G1634,G1296);
  and GNAME1338(G1338,G2865,G1218);
  and GNAME1339(G1339,G2893,G2894);
  and GNAME1340(G1340,G2898,G1339,G2897,G2895,G2896);
  nand GNAME1341(G1341,G3563,G3564);
  and GNAME1342(G1342,G3060,G3061);
  and GNAME1343(G1343,G3065,G3066);
  and GNAME1344(G1344,G3067,G3068);
  nand GNAME1345(G1345,G3063,G3064);
  nand GNAME1346(G1346,G3069,G3070);
  nand GNAME1347(G1347,G3071,G3072);
  nand GNAME1348(G1348,G3073,G3074);
  nand GNAME1349(G1349,G3075,G3076);
  nand GNAME1350(G1350,G3077,G3078);
  nand GNAME1351(G1351,G3079,G3080);
  nand GNAME1352(G1352,G3081,G3082);
  nand GNAME1353(G1353,G3083,G3084);
  nand GNAME1354(G1354,G3085,G3086);
  nand GNAME1355(G1355,G3087,G3088);
  nand GNAME1356(G1356,G3089,G3090);
  nand GNAME1357(G1357,G3091,G3092);
  nand GNAME1358(G1358,G3093,G3094);
  nand GNAME1359(G1359,G3095,G3096);
  nand GNAME1360(G1360,G3097,G3098);
  nand GNAME1361(G1361,G3099,G3100);
  nand GNAME1362(G1362,G3101,G3102);
  nand GNAME1363(G1363,G3103,G3104);
  nand GNAME1364(G1364,G3105,G3106);
  and GNAME1365(G1365,G3107,G3108);
  and GNAME1366(G1366,G3110,G3111);
  and GNAME1367(G1367,G3113,G3114);
  and GNAME1368(G1368,G3116,G3117);
  nand GNAME1369(G1369,G3131,G3132);
  nand GNAME1370(G1370,G3133,G3134);
  nand GNAME1371(G1371,G3135,G3136);
  nand GNAME1372(G1372,G3137,G3138);
  nand GNAME1373(G1373,G3139,G3140);
  nand GNAME1374(G1374,G3141,G3142);
  nand GNAME1375(G1375,G3143,G3144);
  nand GNAME1376(G1376,G3145,G3146);
  nand GNAME1377(G1377,G3147,G3148);
  nand GNAME1378(G1378,G3149,G3150);
  nand GNAME1379(G1379,G3151,G3152);
  nand GNAME1380(G1380,G3153,G3154);
  nand GNAME1381(G1381,G3155,G3156);
  nand GNAME1382(G1382,G3157,G3158);
  nand GNAME1383(G1383,G3159,G3160);
  nand GNAME1384(G1384,G3161,G3162);
  nand GNAME1385(G1385,G3163,G3164);
  nand GNAME1386(G1386,G3165,G3166);
  nand GNAME1387(G1387,G3167,G3168);
  nand GNAME1388(G1388,G3169,G3170);
  nand GNAME1389(G1389,G3171,G3172);
  nand GNAME1390(G1390,G3173,G3174);
  nand GNAME1391(G1391,G3175,G3176);
  nand GNAME1392(G1392,G3177,G3178);
  nand GNAME1393(G1393,G3179,G3180);
  nand GNAME1394(G1394,G3181,G3182);
  nand GNAME1395(G1395,G3183,G3184);
  nand GNAME1396(G1396,G3185,G3186);
  nand GNAME1397(G1397,G3187,G3188);
  nand GNAME1398(G1398,G3189,G3190);
  nand GNAME1399(G1399,G3191,G3192);
  nand GNAME1400(G1400,G3193,G3194);
  and GNAME1401(G1401,G3204,G3205);
  and GNAME1402(G1402,G3207,G3208);
  and GNAME1403(G1403,G3198,G3199);
  and GNAME1404(G1404,G3195,G3196);
  nand GNAME1405(G1405,G3210,G3211);
  nand GNAME1406(G1406,G3212,G3213);
  nand GNAME1407(G1407,G3214,G3215);
  nand GNAME1408(G1408,G3216,G3217);
  nand GNAME1409(G1409,G3218,G3219);
  nand GNAME1410(G1410,G3220,G3221);
  nand GNAME1411(G1411,G3222,G3223);
  nand GNAME1412(G1412,G3224,G3225);
  nand GNAME1413(G1413,G3226,G3227);
  nand GNAME1414(G1414,G3228,G3229);
  nand GNAME1415(G1415,G3230,G3231);
  nand GNAME1416(G1416,G3232,G3233);
  nand GNAME1417(G1417,G3234,G3235);
  nand GNAME1418(G1418,G3236,G3237);
  nand GNAME1419(G1419,G3238,G3239);
  nand GNAME1420(G1420,G3240,G3241);
  nand GNAME1421(G1421,G3242,G3243);
  nand GNAME1422(G1422,G3244,G3245);
  nand GNAME1423(G1423,G3246,G3247);
  nand GNAME1424(G1424,G3248,G3249);
  nand GNAME1425(G1425,G3353,G3354);
  nand GNAME1426(G1426,G3355,G3356);
  nand GNAME1427(G1427,G3357,G3358);
  nand GNAME1428(G1428,G3359,G3360);
  nand GNAME1429(G1429,G3361,G3362);
  nand GNAME1430(G1430,G3363,G3364);
  nand GNAME1431(G1431,G3365,G3366);
  nand GNAME1432(G1432,G3367,G3368);
  nand GNAME1433(G1433,G3369,G3370);
  nand GNAME1434(G1434,G3371,G3372);
  nand GNAME1435(G1435,G3373,G3374);
  nand GNAME1436(G1436,G3375,G3376);
  nand GNAME1437(G1437,G3377,G3378);
  nand GNAME1438(G1438,G3379,G3380);
  nand GNAME1439(G1439,G3381,G3382);
  nand GNAME1440(G1440,G3383,G3384);
  nand GNAME1441(G1441,G3385,G3386);
  nand GNAME1442(G1442,G3387,G3388);
  nand GNAME1443(G1443,G3389,G3390);
  nand GNAME1444(G1444,G3391,G3392);
  nand GNAME1445(G1445,G3393,G3394);
  nand GNAME1446(G1446,G3395,G3396);
  nand GNAME1447(G1447,G3397,G3398);
  nand GNAME1448(G1448,G3399,G3400);
  nand GNAME1449(G1449,G3401,G3402);
  nand GNAME1450(G1450,G3403,G3404);
  nand GNAME1451(G1451,G3405,G3406);
  nand GNAME1452(G1452,G3407,G3408);
  nand GNAME1453(G1453,G3409,G3410);
  nand GNAME1454(G1454,G3411,G3412);
  nand GNAME1455(G1455,G3413,G3414);
  nand GNAME1456(G1456,G3415,G3416);
  nand GNAME1457(G1457,G3425,G3426);
  nand GNAME1458(G1458,G3427,G3428);
  nand GNAME1459(G1459,G3429,G3430);
  nand GNAME1460(G1460,G3431,G3432);
  nand GNAME1461(G1461,G3433,G3434);
  nand GNAME1462(G1462,G3435,G3436);
  nand GNAME1463(G1463,G3437,G3438);
  nand GNAME1464(G1464,G3439,G3440);
  nand GNAME1465(G1465,G3441,G3442);
  nand GNAME1466(G1466,G3443,G3444);
  nand GNAME1467(G1467,G3445,G3446);
  nand GNAME1468(G1468,G3447,G3448);
  nand GNAME1469(G1469,G3449,G3450);
  nand GNAME1470(G1470,G3451,G3452);
  nand GNAME1471(G1471,G3453,G3454);
  nand GNAME1472(G1472,G3455,G3456);
  nand GNAME1473(G1473,G3457,G3458);
  nand GNAME1474(G1474,G3459,G3460);
  nand GNAME1475(G1475,G3461,G3462);
  nand GNAME1476(G1476,G3463,G3464);
  nand GNAME1477(G1477,G3465,G3466);
  nand GNAME1478(G1478,G3467,G3468);
  nand GNAME1479(G1479,G3469,G3470);
  nand GNAME1480(G1480,G3471,G3472);
  nand GNAME1481(G1481,G3473,G3474);
  nand GNAME1482(G1482,G3475,G3476);
  nand GNAME1483(G1483,G3477,G3478);
  nand GNAME1484(G1484,G3479,G3480);
  nand GNAME1485(G1485,G3481,G3482);
  nand GNAME1486(G1486,G3483,G3484);
  nand GNAME1487(G1487,G3485,G3486);
  nand GNAME1488(G1488,G3487,G3488);
  nand GNAME1489(G1489,G3489,G3490);
  nand GNAME1490(G1490,G3491,G3492);
  nand GNAME1491(G1491,G3493,G3494);
  nand GNAME1492(G1492,G3495,G3496);
  nand GNAME1493(G1493,G3497,G3498);
  nand GNAME1494(G1494,G3499,G3500);
  nand GNAME1495(G1495,G3501,G3502);
  nand GNAME1496(G1496,G3503,G3504);
  nand GNAME1497(G1497,G3505,G3506);
  nand GNAME1498(G1498,G3507,G3508);
  nand GNAME1499(G1499,G3509,G3510);
  nand GNAME1500(G1500,G3511,G3512);
  nand GNAME1501(G1501,G3513,G3514);
  nand GNAME1502(G1502,G3515,G3516);
  nand GNAME1503(G1503,G3517,G3518);
  nand GNAME1504(G1504,G3519,G3520);
  nand GNAME1505(G1505,G3521,G3522);
  nand GNAME1506(G1506,G3523,G3524);
  nand GNAME1507(G1507,G3525,G3526);
  nand GNAME1508(G1508,G3527,G3528);
  nand GNAME1509(G1509,G3529,G3530);
  nand GNAME1510(G1510,G3531,G3532);
  nand GNAME1511(G1511,G3533,G3534);
  nand GNAME1512(G1512,G3535,G3536);
  nand GNAME1513(G1513,G3537,G3538);
  nand GNAME1514(G1514,G3539,G3540);
  nand GNAME1515(G1515,G3541,G3542);
  nand GNAME1516(G1516,G3543,G3544);
  nand GNAME1517(G1517,G3545,G3546);
  nand GNAME1518(G1518,G3547,G3548);
  nand GNAME1519(G1519,G3549,G3550);
  nand GNAME1520(G1520,G3551,G3552);
  nand GNAME1521(G1521,G3553,G3554);
  nand GNAME1522(G1522,G3555,G3556);
  nand GNAME1523(G1523,G3557,G3558);
  nand GNAME1524(G1524,G3559,G3560);
  nand GNAME1525(G1525,G3565,G3566);
  nand GNAME1526(G1526,G3567,G3568);
  nand GNAME1527(G1527,G3569,G3570);
  nand GNAME1528(G1528,G3571,G3572);
  nand GNAME1529(G1529,G3573,G3574);
  nand GNAME1530(G1530,G3575,G3576);
  nand GNAME1531(G1531,G3577,G3578);
  nand GNAME1532(G1532,G3579,G3580);
  nand GNAME1533(G1533,G3581,G3582);
  nand GNAME1534(G1534,G3583,G3584);
  nand GNAME1535(G1535,G3585,G3586);
  nand GNAME1536(G1536,G3587,G3588);
  nand GNAME1537(G1537,G3589,G3590);
  nand GNAME1538(G1538,G3591,G3592);
  nand GNAME1539(G1539,G3593,G3594);
  nand GNAME1540(G1540,G3595,G3596);
  nand GNAME1541(G1541,G3597,G3598);
  nand GNAME1542(G1542,G3599,G3600);
  nand GNAME1543(G1543,G3601,G3602);
  nand GNAME1544(G1544,G3603,G3604);
  or GNAME1545(G1545,G22594,G22593,G22592,G22591);
  nor GNAME1546(G1546,G1545,G22595,G22596,G22597,G22598);
  or GNAME1547(G1547,G22602,G22601,G22600,G22599);
  nor GNAME1548(G1548,G1547,G22605,G22603,G22604);
  or GNAME1549(G1549,G22609,G22608,G22607,G22606);
  nor GNAME1550(G1550,G1549,G22612,G22610,G22611);
  or GNAME1551(G1551,G22616,G22615,G22614,G22613);
  nor GNAME1552(G1552,G1551,G22619,G22617,G22618);
  and GNAME1553(G1553,G1795,G1793,G2038);
  and GNAME1554(G1554,G1802,G1800,G1799);
  and GNAME1555(G1555,G1808,G1806,G2073);
  and GNAME1556(G1556,G1815,G1813,G1812);
  and GNAME1557(G1557,G1821,G1819,G2053);
  and GNAME1558(G1558,G1827,G2017,G1826);
  and GNAME1559(G1559,G1833,G1831,G3418);
  and GNAME1560(G1560,G1840,G1838,G1837);
  and GNAME1561(G1561,G1846,G1844,G2043);
  and GNAME1562(G1562,G1852,G2007,G1851);
  and GNAME1563(G1563,G1859,G1857,G1856);
  and GNAME1564(G1564,G1865,G1863,G2063);
  and GNAME1565(G1565,G1872,G1870,G1869);
  and GNAME1566(G1566,G1878,G1876,G2083);
  and GNAME1567(G1567,G1884,G1882,G2028);
  and GNAME1568(G1568,G1890,G1888,G2088);
  and GNAME1569(G1569,G1897,G1895,G1894);
  and GNAME1570(G1570,G1903,G2022,G1902);
  and GNAME1571(G1571,G1909,G1907,G2048);
  and GNAME1572(G1572,G1914,G2002,G1913);
  and GNAME1573(G1573,G1921,G1919,G1918);
  and GNAME1574(G1574,G1927,G1925,G2068);
  and GNAME1575(G1575,G1934,G1932,G1931);
  and GNAME1576(G1576,G1940,G1938,G2058);
  and GNAME1577(G1577,G1946,G2012,G1945);
  and GNAME1578(G1578,G1952,G1950,G2093);
  and GNAME1579(G1579,G1958,G1956,G2033);
  and GNAME1580(G1580,G1965,G1963,G1962);
  and GNAME1581(G1581,G1971,G1969,G2078);
  and GNAME1582(G1582,G3255,G3258,G3261,G3264);
  and GNAME1583(G1583,G1582,G3267,G3270,G3273,G3276);
  and GNAME1584(G1584,G3279,G3282,G3285,G3288);
  and GNAME1585(G1585,G1584,G3291,G3294,G3297,G3300);
  and GNAME1586(G1586,G3303,G3306,G3309,G3312);
  and GNAME1587(G1587,G1586,G3315,G3318,G3321,G3324);
  and GNAME1588(G1588,G3327,G3330,G3333,G3336);
  and GNAME1589(G1589,G1588,G3339,G3342,G3345,G3348);
  and GNAME1590(G1590,G2010,G2012,G2013);
  and GNAME1591(G1591,G2024,G2022,G2023);
  and GNAME1592(G1592,G3059,G3417,G3418);
  and GNAME1593(G1593,G2119,G2120,G2121,G2122);
  and GNAME1594(G1594,G2126,G2127,G2128,G2129);
  and GNAME1595(G1595,G2133,G2134,G2135,G2136);
  and GNAME1596(G1596,G2140,G2141,G2142,G2143);
  and GNAME1597(G1597,G2147,G2148,G2149,G2150);
  and GNAME1598(G1598,G2154,G2155,G2156,G2157);
  and GNAME1599(G1599,G2161,G2162,G2163,G2164);
  and GNAME1600(G1600,G2168,G2169,G2170,G2171);
  and GNAME1601(G1601,G2175,G2176,G2177,G2178);
  and GNAME1602(G1602,G2182,G2183,G2184,G2185);
  and GNAME1603(G1603,G2189,G2190,G2191,G2192);
  and GNAME1604(G1604,G2196,G2197,G2198,G2199);
  and GNAME1605(G1605,G2203,G2204,G2205,G2206);
  and GNAME1606(G1606,G2210,G2211,G2212,G2213);
  and GNAME1607(G1607,G2217,G2218,G2219,G2220);
  and GNAME1608(G1608,G2224,G2225,G2226,G2227);
  and GNAME1609(G1609,G2231,G2232,G2233,G2234);
  and GNAME1610(G1610,G2238,G2239,G2240,G2241);
  and GNAME1611(G1611,G2245,G2246,G2247,G2248);
  and GNAME1612(G1612,G2252,G2253,G2254,G2255);
  and GNAME1613(G1613,G2259,G2260,G2261,G2262);
  and GNAME1614(G1614,G2266,G2267,G2268,G2269);
  and GNAME1615(G1615,G2273,G2274,G2275,G2276);
  and GNAME1616(G1616,G2280,G2281,G2282,G2283);
  and GNAME1617(G1617,G2287,G2288,G2289,G2290);
  and GNAME1618(G1618,G2294,G2295,G2296,G2297);
  and GNAME1619(G1619,G2301,G2302,G2303,G2304);
  and GNAME1620(G1620,G2318,G2316,G2317);
  not GNAME1621(G1621,G22587);
  not GNAME1622(G1622,G7729);
  nor GNAME1623(G1623,G3109,G3112);
  and GNAME1624(G1624,G3423,G3424);
  and GNAME1625(G1625,G1313,G3206,G1402);
  and GNAME1626(G1626,G1313,G1315);
  and GNAME1627(G1627,G1767,G1236);
  not GNAME1628(G1628,G1211);
  not GNAME1629(G1629,G1226);
  not GNAME1630(G1630,G1290);
  not GNAME1631(G1631,G1329);
  not GNAME1632(G1632,G1623);
  nand GNAME1633(G1633,G1783,G1235);
  not GNAME1634(G1634,G1210);
  or GNAME1635(G1635,G1235,G1210);
  nand GNAME1636(G1636,G1635,G1342);
  nand GNAME1637(G1637,G1632,G1636);
  nand GNAME1638(G1638,G3121,G22661);
  nand GNAME1639(G1639,G3124,G22693);
  nand GNAME1640(G1640,G3127,G7990);
  nand GNAME1641(G1641,G3130,G22629);
  nand GNAME1642(G1642,G3121,G22660);
  nand GNAME1643(G1643,G3124,G22692);
  nand GNAME1644(G1644,G3127,G7991);
  nand GNAME1645(G1645,G3130,G22628);
  nand GNAME1646(G1646,G3121,G22659);
  nand GNAME1647(G1647,G3124,G22691);
  nand GNAME1648(G1648,G3127,G7992);
  nand GNAME1649(G1649,G3130,G22627);
  nand GNAME1650(G1650,G3121,G22658);
  nand GNAME1651(G1651,G3124,G22690);
  nand GNAME1652(G1652,G3127,G7993);
  nand GNAME1653(G1653,G3130,G22626);
  nand GNAME1654(G1654,G3121,G22657);
  nand GNAME1655(G1655,G3124,G22689);
  nand GNAME1656(G1656,G3127,G7994);
  nand GNAME1657(G1657,G3130,G22625);
  nand GNAME1658(G1658,G3121,G22656);
  nand GNAME1659(G1659,G3124,G22688);
  nand GNAME1660(G1660,G3127,G7995);
  nand GNAME1661(G1661,G3130,G22624);
  nand GNAME1662(G1662,G3121,G22655);
  nand GNAME1663(G1663,G3124,G22687);
  nand GNAME1664(G1664,G3127,G7959);
  nand GNAME1665(G1665,G3130,G22623);
  nand GNAME1666(G1666,G3130,G22651);
  nand GNAME1667(G1667,G3121,G22683);
  nand GNAME1668(G1668,G3124,G22715);
  nand GNAME1669(G1669,G3130,G22650);
  nand GNAME1670(G1670,G3121,G22682);
  nand GNAME1671(G1671,G3124,G22714);
  nand GNAME1672(G1672,G3121,G22654);
  nand GNAME1673(G1673,G3124,G22686);
  nand GNAME1674(G1674,G3127,G22773);
  nand GNAME1675(G1675,G3130,G22622);
  nand GNAME1676(G1676,G3130,G22649);
  nand GNAME1677(G1677,G3121,G22681);
  nand GNAME1678(G1678,G3124,G22713);
  nand GNAME1679(G1679,G3127,G7960);
  nand GNAME1680(G1680,G3127,G7996);
  nand GNAME1681(G1681,G3130,G22648);
  nand GNAME1682(G1682,G3121,G22680);
  nand GNAME1683(G1683,G3124,G22712);
  nand GNAME1684(G1684,G3127,G7997);
  nand GNAME1685(G1685,G3130,G22647);
  nand GNAME1686(G1686,G3121,G22679);
  nand GNAME1687(G1687,G3124,G22711);
  nand GNAME1688(G1688,G3127,G7998);
  nand GNAME1689(G1689,G3130,G22646);
  nand GNAME1690(G1690,G3121,G22678);
  nand GNAME1691(G1691,G3124,G22710);
  nand GNAME1692(G1692,G3127,G7999);
  nand GNAME1693(G1693,G3130,G22645);
  nand GNAME1694(G1694,G3121,G22677);
  nand GNAME1695(G1695,G3124,G22709);
  nand GNAME1696(G1696,G3127,G8000);
  nand GNAME1697(G1697,G3130,G22644);
  nand GNAME1698(G1698,G3121,G22676);
  nand GNAME1699(G1699,G3124,G22708);
  nand GNAME1700(G1700,G3127,G8001);
  nand GNAME1701(G1701,G3130,G22643);
  nand GNAME1702(G1702,G3121,G22675);
  nand GNAME1703(G1703,G3124,G22707);
  nand GNAME1704(G1704,G3127,G8002);
  nand GNAME1705(G1705,G3130,G22642);
  nand GNAME1706(G1706,G3121,G22674);
  nand GNAME1707(G1707,G3124,G22706);
  nand GNAME1708(G1708,G3127,G8003);
  nand GNAME1709(G1709,G3130,G22641);
  nand GNAME1710(G1710,G3121,G22673);
  nand GNAME1711(G1711,G3124,G22705);
  nand GNAME1712(G1712,G3127,G8004);
  nand GNAME1713(G1713,G3130,G22640);
  nand GNAME1714(G1714,G3121,G22672);
  nand GNAME1715(G1715,G3124,G22704);
  nand GNAME1716(G1716,G3130,G22621);
  nand GNAME1717(G1717,G3121,G22653);
  nand GNAME1718(G1718,G3124,G22685);
  nand GNAME1719(G1719,G3127,G22788);
  nand GNAME1720(G1720,G3121,G22671);
  nand GNAME1721(G1721,G3124,G22703);
  nand GNAME1722(G1722,G3127,G8005);
  nand GNAME1723(G1723,G3130,G22639);
  nand GNAME1724(G1724,G3121,G22670);
  nand GNAME1725(G1725,G3124,G22702);
  nand GNAME1726(G1726,G3127,G8006);
  nand GNAME1727(G1727,G3130,G22638);
  nand GNAME1728(G1728,G3121,G22669);
  nand GNAME1729(G1729,G3124,G22701);
  nand GNAME1730(G1730,G3127,G8007);
  nand GNAME1731(G1731,G3130,G22637);
  nand GNAME1732(G1732,G3121,G22668);
  nand GNAME1733(G1733,G3124,G22700);
  nand GNAME1734(G1734,G3127,G8008);
  nand GNAME1735(G1735,G3130,G22636);
  nand GNAME1736(G1736,G3121,G22667);
  nand GNAME1737(G1737,G3124,G22699);
  nand GNAME1738(G1738,G3127,G8009);
  nand GNAME1739(G1739,G3130,G22635);
  nand GNAME1740(G1740,G3121,G22666);
  nand GNAME1741(G1741,G3124,G22698);
  nand GNAME1742(G1742,G3127,G8010);
  nand GNAME1743(G1743,G3130,G22634);
  nand GNAME1744(G1744,G3121,G22665);
  nand GNAME1745(G1745,G3124,G22697);
  nand GNAME1746(G1746,G3127,G8011);
  nand GNAME1747(G1747,G3130,G22633);
  nand GNAME1748(G1748,G3121,G22664);
  nand GNAME1749(G1749,G3124,G22696);
  nand GNAME1750(G1750,G3127,G8012);
  nand GNAME1751(G1751,G3130,G22632);
  nand GNAME1752(G1752,G3121,G22663);
  nand GNAME1753(G1753,G3124,G22695);
  nand GNAME1754(G1754,G3127,G8013);
  nand GNAME1755(G1755,G3130,G22631);
  nand GNAME1756(G1756,G3121,G22662);
  nand GNAME1757(G1757,G3124,G22694);
  nand GNAME1758(G1758,G3127,G8014);
  nand GNAME1759(G1759,G3130,G22630);
  nand GNAME1760(G1760,G3130,G22620);
  nand GNAME1761(G1761,G3121,G22652);
  nand GNAME1762(G1762,G3124,G22684);
  nand GNAME1763(G1763,G3127,G22778);
  not GNAME1764(G1764,G1303);
  or GNAME1765(G1765,G3115,G1629);
  and GNAME1766(G1766,G1345,G3203);
  not GNAME1767(G1767,G1217);
  nand GNAME1768(G1768,G1546,G1548,G1550,G1552);
  nand GNAME1769(G1769,G1768,G1217);
  nand GNAME1770(G1770,G1217,G22590);
  nand GNAME1771(G1771,G1343,G1344);
  nand GNAME1772(G1772,G1343,G1345);
  not GNAME1773(G1773,G1220);
  or GNAME1774(G1774,G3115,G1229);
  or GNAME1775(G1775,G3605,G3118);
  not GNAME1776(G1776,G1288);
  nand GNAME1777(G1777,G3115,G1230);
  or GNAME1778(G1778,G1295,G3118);
  nand GNAME1779(G1779,G1241,G1227);
  nand GNAME1780(G1780,G1237,G1240);
  nand GNAME1781(G1781,G1236,G1242);
  nand GNAME1782(G1782,G1780,G1781);
  or GNAME1783(G1783,G3200,G3197);
  or GNAME1784(G1784,G1234,G1240,G1233);
  nand GNAME1785(G1785,G1773,G1784);
  nand GNAME1786(G1786,G1785,G1633);
  nand GNAME1787(G1787,G1786,G1236);
  nand GNAME1788(G1788,G1773,G1221);
  nand GNAME1789(G1789,G1630,G1294,G1787,G1788);
  nand GNAME1790(G1790,G1263,G1222);
  nand GNAME1791(G1791,G1265,G1223);
  nand GNAME1792(G1792,G1789,G7992);
  nand GNAME1793(G1793,G7012,G1238);
  nand GNAME1794(G1794,G8178,G1239);
  nand GNAME1795(G1795,G1782,G1405);
  nand GNAME1796(G1796,G1283,G1222);
  nand GNAME1797(G1797,G1285,G1223);
  nand GNAME1798(G1798,G1789,G7997);
  nand GNAME1799(G1799,G1066,G22796);
  nand GNAME1800(G1800,G1238,G7068);
  nand GNAME1801(G1801,G8187,G1239);
  nand GNAME1802(G1802,G1782,G1243);
  nand GNAME1803(G1803,G1270,G1222);
  nand GNAME1804(G1804,G1272,G1223);
  nand GNAME1805(G1805,G1789,G8010);
  nand GNAME1806(G1806,G1238,G7016);
  nand GNAME1807(G1807,G8200,G1239);
  nand GNAME1808(G1808,G1782,G1406);
  nand GNAME1809(G1809,G1279,G1222);
  nand GNAME1810(G1810,G1281,G1223);
  nand GNAME1811(G1811,G1789,G8001);
  nand GNAME1812(G1812,G1066,G22794);
  nand GNAME1813(G1813,G1238,G7080);
  nand GNAME1814(G1814,G8191,G1239);
  nand GNAME1815(G1815,G1782,G1244);
  nand GNAME1816(G1816,G1266,G1222);
  nand GNAME1817(G1817,G1268,G1223);
  nand GNAME1818(G1818,G1789,G8014);
  nand GNAME1819(G1819,G1238,G6973);
  nand GNAME1820(G1820,G8204,G1239);
  nand GNAME1821(G1821,G1782,G1407);
  nand GNAME1822(G1822,G1259,G1222);
  nand GNAME1823(G1823,G1261,G1223);
  nand GNAME1824(G1824,G1789,G7959);
  nand GNAME1825(G1825,G1238,G7013);
  nand GNAME1826(G1826,G8182,G1239);
  nand GNAME1827(G1827,G1782,G1408);
  nand GNAME1828(G1828,G1275,G1222);
  nand GNAME1829(G1829,G1277,G1223);
  nand GNAME1830(G1830,G1789,G8005);
  nand GNAME1831(G1831,G1238,G7095);
  nand GNAME1832(G1832,G8195,G1239);
  nand GNAME1833(G1833,G1782,G1409);
  nand GNAME1834(G1834,G1284,G1222);
  nand GNAME1835(G1835,G1254,G1223);
  nand GNAME1836(G1836,G1789,G7996);
  nand GNAME1837(G1837,G1066,G22790);
  nand GNAME1838(G1838,G1238,G7065);
  nand GNAME1839(G1839,G8186,G1239);
  nand GNAME1840(G1840,G1782,G1245);
  nand GNAME1841(G1841,G1264,G1222);
  nand GNAME1842(G1842,G1266,G1223);
  nand GNAME1843(G1843,G1789,G7991);
  nand GNAME1844(G1844,G1238,G7031);
  nand GNAME1845(G1845,G8177,G1239);
  nand GNAME1846(G1846,G1782,G1410);
  nand GNAME1847(G1847,G1257,G1222);
  nand GNAME1848(G1848,G1259,G1223);
  nand GNAME1849(G1849,G1789,G22788);
  nand GNAME1850(G1850,G1238,G7092);
  nand GNAME1851(G1851,G8175,G1239);
  nand GNAME1852(G1852,G1782,G1411);
  nand GNAME1853(G1853,G1277,G1222);
  nand GNAME1854(G1854,G1279,G1223);
  nand GNAME1855(G1855,G1789,G8003);
  nand GNAME1856(G1856,G1066,G22787);
  nand GNAME1857(G1857,G1238,G7086);
  nand GNAME1858(G1858,G8193,G1239);
  nand GNAME1859(G1859,G1782,G1246);
  nand GNAME1860(G1860,G1268,G1222);
  nand GNAME1861(G1861,G1270,G1223);
  nand GNAME1862(G1862,G1789,G8012);
  nand GNAME1863(G1863,G1238,G7114);
  nand GNAME1864(G1864,G8202,G1239);
  nand GNAME1865(G1865,G1782,G1412);
  nand GNAME1866(G1866,G1281,G1222);
  nand GNAME1867(G1867,G1283,G1223);
  nand GNAME1868(G1868,G1789,G7999);
  nand GNAME1869(G1869,G1066,G22785);
  nand GNAME1870(G1870,G1238,G7074);
  nand GNAME1871(G1871,G8189,G1239);
  nand GNAME1872(G1872,G1782,G1247);
  nand GNAME1873(G1873,G1272,G1222);
  nand GNAME1874(G1874,G1274,G1223);
  nand GNAME1875(G1875,G1789,G8008);
  nand GNAME1876(G1876,G1238,G7104);
  nand GNAME1877(G1877,G8198,G1239);
  nand GNAME1878(G1878,G1782,G1413);
  nand GNAME1879(G1879,G1261,G1222);
  nand GNAME1880(G1880,G1263,G1223);
  nand GNAME1881(G1881,G1789,G7994);
  nand GNAME1882(G1882,G1238,G7035);
  nand GNAME1883(G1883,G8180,G1239);
  nand GNAME1884(G1884,G1782,G1414);
  nand GNAME1885(G1885,G1273,G1222);
  nand GNAME1886(G1886,G1275,G1223);
  nand GNAME1887(G1887,G1789,G8007);
  nand GNAME1888(G1888,G1238,G7101);
  nand GNAME1889(G1889,G8197,G1239);
  nand GNAME1890(G1890,G1782,G1415);
  nand GNAME1891(G1891,G1280,G1222);
  nand GNAME1892(G1892,G1282,G1223);
  nand GNAME1893(G1893,G1789,G8000);
  nand GNAME1894(G1894,G1066,G22781);
  nand GNAME1895(G1895,G1238,G7077);
  nand GNAME1896(G1896,G8190,G1239);
  nand GNAME1897(G1897,G1782,G1248);
  nand GNAME1898(G1898,G1260,G1222);
  nand GNAME1899(G1899,G1262,G1223);
  nand GNAME1900(G1900,G1789,G7995);
  nand GNAME1901(G1901,G1238,G7038);
  nand GNAME1902(G1902,G8181,G1239);
  nand GNAME1903(G1903,G1782,G1416);
  nand GNAME1904(G1904,G1265,G1222);
  nand GNAME1905(G1905,G1267,G1223);
  nand GNAME1906(G1906,G1789,G7990);
  nand GNAME1907(G1907,G1238,G7028);
  nand GNAME1908(G1908,G8176,G1239);
  nand GNAME1909(G1909,G1782,G1417);
  nand GNAME1910(G1910,G1258,G1223);
  nand GNAME1911(G1911,G1789,G22778);
  nand GNAME1912(G1912,G1238,G7011);
  nand GNAME1913(G1913,G8085,G1239);
  nand GNAME1914(G1914,G1782,G1418);
  nand GNAME1915(G1915,G1276,G1222);
  nand GNAME1916(G1916,G1278,G1223);
  nand GNAME1917(G1917,G1789,G8004);
  nand GNAME1918(G1918,G1066,G22777);
  nand GNAME1919(G1919,G1238,G7089);
  nand GNAME1920(G1920,G8194,G1239);
  nand GNAME1921(G1921,G1782,G1249);
  nand GNAME1922(G1922,G1269,G1222);
  nand GNAME1923(G1923,G1271,G1223);
  nand GNAME1924(G1924,G1789,G8011);
  nand GNAME1925(G1925,G1238,G7111);
  nand GNAME1926(G1926,G8201,G1239);
  nand GNAME1927(G1927,G1782,G1419);
  nand GNAME1928(G1928,G1278,G1222);
  nand GNAME1929(G1929,G1280,G1223);
  nand GNAME1930(G1930,G1789,G8002);
  nand GNAME1931(G1931,G1066,G22775);
  nand GNAME1932(G1932,G1238,G7083);
  nand GNAME1933(G1933,G8192,G1239);
  nand GNAME1934(G1934,G1782,G1250);
  nand GNAME1935(G1935,G1267,G1222);
  nand GNAME1936(G1936,G1269,G1223);
  nand GNAME1937(G1937,G1789,G8013);
  nand GNAME1938(G1938,G1238,G7017);
  nand GNAME1939(G1939,G8203,G1239);
  nand GNAME1940(G1940,G1782,G1420);
  nand GNAME1941(G1941,G1258,G1222);
  nand GNAME1942(G1942,G1260,G1223);
  nand GNAME1943(G1943,G1789,G22773);
  nand GNAME1944(G1944,G1238,G6974);
  nand GNAME1945(G1945,G8184,G1239);
  nand GNAME1946(G1946,G1782,G1421);
  nand GNAME1947(G1947,G1274,G1222);
  nand GNAME1948(G1948,G1276,G1223);
  nand GNAME1949(G1949,G1789,G8006);
  nand GNAME1950(G1950,G1238,G7098);
  nand GNAME1951(G1951,G8196,G1239);
  nand GNAME1952(G1952,G1782,G1422);
  nand GNAME1953(G1953,G1262,G1222);
  nand GNAME1954(G1954,G1264,G1223);
  nand GNAME1955(G1955,G1789,G7993);
  nand GNAME1956(G1956,G1238,G6975);
  nand GNAME1957(G1957,G8179,G1239);
  nand GNAME1958(G1958,G1782,G1423);
  nand GNAME1959(G1959,G1282,G1222);
  nand GNAME1960(G1960,G1284,G1223);
  nand GNAME1961(G1961,G1789,G7998);
  nand GNAME1962(G1962,G1066,G22770);
  nand GNAME1963(G1963,G1238,G7071);
  nand GNAME1964(G1964,G8188,G1239);
  nand GNAME1965(G1965,G1782,G1251);
  nand GNAME1966(G1966,G1271,G1222);
  nand GNAME1967(G1967,G1273,G1223);
  nand GNAME1968(G1968,G1789,G8009);
  nand GNAME1969(G1969,G1238,G7107);
  nand GNAME1970(G1970,G8199,G1239);
  nand GNAME1971(G1971,G1782,G1424);
  nor GNAME1972(G1972,G3197,G3118);
  or GNAME1973(G1973,G1972,G1235);
  nand GNAME1974(G1974,G1286,G1289);
  nand GNAME1975(G1975,G1974,G3349,G3350);
  or GNAME1976(G1976,G1629,G7603);
  or GNAME1977(G1977,G7729,G3118);
  nand GNAME1978(G1978,G1976,G1977);
  nand GNAME1979(G1979,G1978,G1288);
  nand GNAME1980(G1980,G1975,G1403);
  nand GNAME1981(G1981,G1979,G1980);
  nand GNAME1982(G1982,G3252,G1404);
  or GNAME1983(G1983,G1289,G3607);
  nand GNAME1984(G1984,G1982,G1983);
  nand GNAME1985(G1985,G1984,G1287);
  nand GNAME1986(G1986,G1981,G3062);
  nand GNAME1987(G1987,G1985,G1986);
  nand GNAME1988(G1988,G3351,G3352,G22798,G1628);
  nand GNAME1989(G1989,G1252,G1622,G1236);
  nand GNAME1990(G1990,G1988,G22768);
  nand GNAME1991(G1991,G22798,G1987);
  not GNAME1992(G1992,G1300);
  nand GNAME1993(G1993,G1297,G1292);
  nand GNAME1994(G1994,G1294,G1993);
  or GNAME1995(G1995,G1296,G1297);
  or GNAME1996(G1996,G1294,G1300,G3112);
  nand GNAME1997(G1997,G1292,G1298);
  nand GNAME1998(G1998,G1996,G1997);
  nand GNAME1999(G1999,G7011,G1293);
  nand GNAME2000(G2000,G1998,G1364);
  nand GNAME2001(G2001,G1299,G7433);
  nand GNAME2002(G2002,G1066,G22778);
  nand GNAME2003(G2003,G1300,G22735);
  nand GNAME2004(G2004,G7092,G1293);
  nand GNAME2005(G2005,G1998,G1354);
  nand GNAME2006(G2006,G1299,G7432);
  nand GNAME2007(G2007,G1066,G22788);
  nand GNAME2008(G2008,G1300,G22734);
  nand GNAME2009(G2009,G6974,G1293);
  nand GNAME2010(G2010,G1998,G1353);
  nand GNAME2011(G2011,G1299,G7455);
  nand GNAME2012(G2012,G1066,G22773);
  nand GNAME2013(G2013,G1300,G22733);
  nand GNAME2014(G2014,G7013,G1293);
  nand GNAME2015(G2015,G1998,G1352);
  nand GNAME2016(G2016,G1299,G7454);
  nand GNAME2017(G2017,G1066,G22792);
  nand GNAME2018(G2018,G1300,G22732);
  nand GNAME2019(G2019,G7038,G1293);
  nand GNAME2020(G2020,G1998,G1351);
  nand GNAME2021(G2021,G1299,G7431);
  nand GNAME2022(G2022,G1066,G22780);
  nand GNAME2023(G2023,G1300,G22731);
  nand GNAME2024(G2024,G1290,G1524);
  nand GNAME2025(G2025,G7035,G1293);
  nand GNAME2026(G2026,G1998,G1350);
  nand GNAME2027(G2027,G1299,G7451);
  nand GNAME2028(G2028,G1066,G22783);
  nand GNAME2029(G2029,G1300,G22730);
  nand GNAME2030(G2030,G6975,G1293);
  nand GNAME2031(G2031,G1998,G1349);
  nand GNAME2032(G2032,G1299,G7430);
  nand GNAME2033(G2033,G1066,G22771);
  nand GNAME2034(G2034,G1300,G22729);
  nand GNAME2035(G2035,G7012,G1293);
  nand GNAME2036(G2036,G1998,G1348);
  nand GNAME2037(G2037,G1299,G7450);
  nand GNAME2038(G2038,G1066,G22797);
  nand GNAME2039(G2039,G1300,G22728);
  nand GNAME2040(G2040,G7031,G1293);
  nand GNAME2041(G2041,G1998,G1347);
  nand GNAME2042(G2042,G1299,G7449);
  nand GNAME2043(G2043,G1066,G22789);
  nand GNAME2044(G2044,G1300,G22727);
  nand GNAME2045(G2045,G7028,G1293);
  nand GNAME2046(G2046,G1998,G1346);
  nand GNAME2047(G2047,G1299,G7448);
  nand GNAME2048(G2048,G1066,G22779);
  nand GNAME2049(G2049,G1300,G22726);
  nand GNAME2050(G2050,G6973,G1293);
  nand GNAME2051(G2051,G1998,G1363);
  nand GNAME2052(G2052,G1299,G7388);
  nand GNAME2053(G2053,G1066,G22793);
  nand GNAME2054(G2054,G1300,G22725);
  nand GNAME2055(G2055,G7017,G1293);
  nand GNAME2056(G2056,G1998,G1362);
  nand GNAME2057(G2057,G1299,G7434);
  nand GNAME2058(G2058,G1066,G22774);
  nand GNAME2059(G2059,G1300,G22724);
  nand GNAME2060(G2060,G7114,G1293);
  nand GNAME2061(G2061,G1998,G1361);
  nand GNAME2062(G2062,G1299,G7462);
  nand GNAME2063(G2063,G1066,G22786);
  nand GNAME2064(G2064,G1300,G22723);
  nand GNAME2065(G2065,G7111,G1293);
  nand GNAME2066(G2066,G1998,G1360);
  nand GNAME2067(G2067,G1299,G7461);
  nand GNAME2068(G2068,G1066,G22776);
  nand GNAME2069(G2069,G1300,G22722);
  nand GNAME2070(G2070,G7016,G1293);
  nand GNAME2071(G2071,G1998,G1359);
  nand GNAME2072(G2072,G1299,G7389);
  nand GNAME2073(G2073,G1066,G22795);
  nand GNAME2074(G2074,G1300,G22721);
  nand GNAME2075(G2075,G7107,G1293);
  nand GNAME2076(G2076,G1998,G1358);
  nand GNAME2077(G2077,G1299,G7390);
  nand GNAME2078(G2078,G1066,G22769);
  nand GNAME2079(G2079,G1300,G22720);
  nand GNAME2080(G2080,G7104,G1293);
  nand GNAME2081(G2081,G1998,G1357);
  nand GNAME2082(G2082,G1299,G7460);
  nand GNAME2083(G2083,G1066,G22784);
  nand GNAME2084(G2084,G1300,G22719);
  nand GNAME2085(G2085,G7101,G1293);
  nand GNAME2086(G2086,G1998,G1356);
  nand GNAME2087(G2087,G1299,G7459);
  nand GNAME2088(G2088,G1066,G22782);
  nand GNAME2089(G2089,G1300,G22718);
  nand GNAME2090(G2090,G7098,G1293);
  nand GNAME2091(G2091,G1998,G1355);
  nand GNAME2092(G2092,G1299,G7458);
  nand GNAME2093(G2093,G1066,G22772);
  nand GNAME2094(G2094,G1300,G22717);
  nand GNAME2095(G2095,G1298,G3200,G1292);
  nand GNAME2096(G2096,G7095,G1293);
  nand GNAME2097(G2097,G1299,G7391);
  and GNAME2098(G2098,G1633,G3209,G1219,G1401);
  or GNAME2099(G2099,G1242,G2098);
  not GNAME2100(G2100,G1301);
  nand GNAME2101(G2101,G1235,G902,G2111);
  nand GNAME2102(G2102,G8084,G1303);
  nand GNAME2103(G2103,G2102,G2101);
  nand GNAME2104(G2104,G1255,G1302);
  nand GNAME2105(G2105,G8183,G1303);
  nand GNAME2106(G2106,G2105,G2101);
  nand GNAME2107(G2107,G1256,G1302);
  or GNAME2108(G2108,G1367,G1403);
  nand GNAME2109(G2109,G2108,G1304);
  or GNAME2110(G2110,G22768,G3112);
  nand GNAME2111(G2111,G2110,G1632);
  nand GNAME2112(G2112,G904,G2111);
  nand GNAME2113(G2113,G1285,G3112);
  nand GNAME2114(G2114,G2112,G2113);
  nand GNAME2115(G2115,G7062,G1305);
  nand GNAME2116(G2116,G8185,G1306);
  nand GNAME2117(G2117,G7960,G1307);
  nand GNAME2118(G2118,G1253,G1302);
  nand GNAME2119(G2119,G7065,G1305);
  nand GNAME2120(G2120,G8186,G1306);
  nand GNAME2121(G2121,G7996,G1307);
  nand GNAME2122(G2122,G2100,G22712);
  nand GNAME2123(G2123,G1254,G1309);
  nand GNAME2124(G2124,G1284,G1311);
  nand GNAME2125(G2125,G1245,G1302);
  nand GNAME2126(G2126,G7068,G1305);
  nand GNAME2127(G2127,G8187,G1306);
  nand GNAME2128(G2128,G7997,G1307);
  nand GNAME2129(G2129,G2100,G22711);
  nand GNAME2130(G2130,G1283,G1311);
  nand GNAME2131(G2131,G1243,G1302);
  nand GNAME2132(G2132,G1285,G1309);
  nand GNAME2133(G2133,G7071,G1305);
  nand GNAME2134(G2134,G8188,G1306);
  nand GNAME2135(G2135,G7998,G1307);
  nand GNAME2136(G2136,G2100,G22710);
  nand GNAME2137(G2137,G1282,G1311);
  nand GNAME2138(G2138,G1251,G1302);
  nand GNAME2139(G2139,G1284,G1309);
  nand GNAME2140(G2140,G7074,G1305);
  nand GNAME2141(G2141,G8189,G1306);
  nand GNAME2142(G2142,G7999,G1307);
  nand GNAME2143(G2143,G2100,G22709);
  nand GNAME2144(G2144,G1281,G1311);
  nand GNAME2145(G2145,G1247,G1302);
  nand GNAME2146(G2146,G1283,G1309);
  nand GNAME2147(G2147,G7077,G1305);
  nand GNAME2148(G2148,G8190,G1306);
  nand GNAME2149(G2149,G8000,G1307);
  nand GNAME2150(G2150,G2100,G22708);
  nand GNAME2151(G2151,G1280,G1311);
  nand GNAME2152(G2152,G1248,G1302);
  nand GNAME2153(G2153,G1282,G1309);
  nand GNAME2154(G2154,G7080,G1305);
  nand GNAME2155(G2155,G8191,G1306);
  nand GNAME2156(G2156,G8001,G1307);
  nand GNAME2157(G2157,G2100,G22707);
  nand GNAME2158(G2158,G1279,G1311);
  nand GNAME2159(G2159,G1244,G1302);
  nand GNAME2160(G2160,G1281,G1309);
  nand GNAME2161(G2161,G7083,G1305);
  nand GNAME2162(G2162,G8192,G1306);
  nand GNAME2163(G2163,G8002,G1307);
  nand GNAME2164(G2164,G2100,G22706);
  nand GNAME2165(G2165,G1278,G1311);
  nand GNAME2166(G2166,G1250,G1302);
  nand GNAME2167(G2167,G1280,G1309);
  nand GNAME2168(G2168,G7086,G1305);
  nand GNAME2169(G2169,G8193,G1306);
  nand GNAME2170(G2170,G8003,G1307);
  nand GNAME2171(G2171,G2100,G22705);
  nand GNAME2172(G2172,G1277,G1311);
  nand GNAME2173(G2173,G1246,G1302);
  nand GNAME2174(G2174,G1279,G1309);
  nand GNAME2175(G2175,G7089,G1305);
  nand GNAME2176(G2176,G8194,G1306);
  nand GNAME2177(G2177,G8004,G1307);
  nand GNAME2178(G2178,G2100,G22704);
  nand GNAME2179(G2179,G1276,G1311);
  nand GNAME2180(G2180,G1249,G1302);
  nand GNAME2181(G2181,G1278,G1309);
  nand GNAME2182(G2182,G7095,G1305);
  nand GNAME2183(G2183,G8195,G1306);
  nand GNAME2184(G2184,G2100,G22703);
  nand GNAME2185(G2185,G8005,G1307);
  nand GNAME2186(G2186,G1275,G1311);
  nand GNAME2187(G2187,G1409,G1302);
  nand GNAME2188(G2188,G1277,G1309);
  nand GNAME2189(G2189,G7098,G1305);
  nand GNAME2190(G2190,G8196,G1306);
  nand GNAME2191(G2191,G2100,G22702);
  nand GNAME2192(G2192,G8006,G1307);
  nand GNAME2193(G2193,G1274,G1311);
  nand GNAME2194(G2194,G1422,G1302);
  nand GNAME2195(G2195,G1276,G1309);
  nand GNAME2196(G2196,G7101,G1305);
  nand GNAME2197(G2197,G8197,G1306);
  nand GNAME2198(G2198,G2100,G22701);
  nand GNAME2199(G2199,G8007,G1307);
  nand GNAME2200(G2200,G1273,G1311);
  nand GNAME2201(G2201,G1415,G1302);
  nand GNAME2202(G2202,G1275,G1309);
  nand GNAME2203(G2203,G7104,G1305);
  nand GNAME2204(G2204,G8198,G1306);
  nand GNAME2205(G2205,G2100,G22700);
  nand GNAME2206(G2206,G8008,G1307);
  nand GNAME2207(G2207,G1272,G1311);
  nand GNAME2208(G2208,G1413,G1302);
  nand GNAME2209(G2209,G1274,G1309);
  nand GNAME2210(G2210,G7107,G1305);
  nand GNAME2211(G2211,G8199,G1306);
  nand GNAME2212(G2212,G2100,G22699);
  nand GNAME2213(G2213,G8009,G1307);
  nand GNAME2214(G2214,G1271,G1311);
  nand GNAME2215(G2215,G1424,G1302);
  nand GNAME2216(G2216,G1273,G1309);
  nand GNAME2217(G2217,G7016,G1305);
  nand GNAME2218(G2218,G8200,G1306);
  nand GNAME2219(G2219,G2100,G22698);
  nand GNAME2220(G2220,G8010,G1307);
  nand GNAME2221(G2221,G1270,G1311);
  nand GNAME2222(G2222,G1406,G1302);
  nand GNAME2223(G2223,G1272,G1309);
  nand GNAME2224(G2224,G7111,G1305);
  nand GNAME2225(G2225,G8201,G1306);
  nand GNAME2226(G2226,G2100,G22697);
  nand GNAME2227(G2227,G8011,G1307);
  nand GNAME2228(G2228,G1269,G1311);
  nand GNAME2229(G2229,G1419,G1302);
  nand GNAME2230(G2230,G1271,G1309);
  nand GNAME2231(G2231,G7114,G1305);
  nand GNAME2232(G2232,G8202,G1306);
  nand GNAME2233(G2233,G2100,G22696);
  nand GNAME2234(G2234,G8012,G1307);
  nand GNAME2235(G2235,G1268,G1311);
  nand GNAME2236(G2236,G1412,G1302);
  nand GNAME2237(G2237,G1270,G1309);
  nand GNAME2238(G2238,G7017,G1305);
  nand GNAME2239(G2239,G8203,G1306);
  nand GNAME2240(G2240,G2100,G22695);
  nand GNAME2241(G2241,G8013,G1307);
  nand GNAME2242(G2242,G1267,G1311);
  nand GNAME2243(G2243,G1420,G1302);
  nand GNAME2244(G2244,G1269,G1309);
  nand GNAME2245(G2245,G6973,G1305);
  nand GNAME2246(G2246,G8204,G1306);
  nand GNAME2247(G2247,G2100,G22694);
  nand GNAME2248(G2248,G8014,G1307);
  nand GNAME2249(G2249,G1266,G1311);
  nand GNAME2250(G2250,G1407,G1302);
  nand GNAME2251(G2251,G1268,G1309);
  nand GNAME2252(G2252,G7028,G1305);
  nand GNAME2253(G2253,G8176,G1306);
  nand GNAME2254(G2254,G2100,G22693);
  nand GNAME2255(G2255,G7990,G1307);
  nand GNAME2256(G2256,G1265,G1311);
  nand GNAME2257(G2257,G1417,G1302);
  nand GNAME2258(G2258,G1267,G1309);
  nand GNAME2259(G2259,G7031,G1305);
  nand GNAME2260(G2260,G8177,G1306);
  nand GNAME2261(G2261,G2100,G22692);
  nand GNAME2262(G2262,G7991,G1307);
  nand GNAME2263(G2263,G1264,G1311);
  nand GNAME2264(G2264,G1410,G1302);
  nand GNAME2265(G2265,G1266,G1309);
  nand GNAME2266(G2266,G7012,G1305);
  nand GNAME2267(G2267,G8178,G1306);
  nand GNAME2268(G2268,G2100,G22691);
  nand GNAME2269(G2269,G7992,G1307);
  nand GNAME2270(G2270,G1263,G1311);
  nand GNAME2271(G2271,G1405,G1302);
  nand GNAME2272(G2272,G1265,G1309);
  nand GNAME2273(G2273,G6975,G1305);
  nand GNAME2274(G2274,G8179,G1306);
  nand GNAME2275(G2275,G2100,G22690);
  nand GNAME2276(G2276,G7993,G1307);
  nand GNAME2277(G2277,G1262,G1311);
  nand GNAME2278(G2278,G1423,G1302);
  nand GNAME2279(G2279,G1264,G1309);
  nand GNAME2280(G2280,G7035,G1305);
  nand GNAME2281(G2281,G8180,G1306);
  nand GNAME2282(G2282,G2100,G22689);
  nand GNAME2283(G2283,G7994,G1307);
  nand GNAME2284(G2284,G1261,G1311);
  nand GNAME2285(G2285,G1414,G1302);
  nand GNAME2286(G2286,G1263,G1309);
  nand GNAME2287(G2287,G7038,G1305);
  nand GNAME2288(G2288,G8181,G1306);
  nand GNAME2289(G2289,G2100,G22688);
  nand GNAME2290(G2290,G7995,G1307);
  nand GNAME2291(G2291,G1260,G1311);
  nand GNAME2292(G2292,G1416,G1302);
  nand GNAME2293(G2293,G1262,G1309);
  nand GNAME2294(G2294,G7013,G1305);
  nand GNAME2295(G2295,G8182,G1306);
  nand GNAME2296(G2296,G2100,G22687);
  nand GNAME2297(G2297,G7959,G1307);
  nand GNAME2298(G2298,G1259,G1311);
  nand GNAME2299(G2299,G1408,G1302);
  nand GNAME2300(G2300,G1261,G1309);
  nand GNAME2301(G2301,G6974,G1305);
  nand GNAME2302(G2302,G8184,G1306);
  nand GNAME2303(G2303,G2100,G22686);
  nand GNAME2304(G2304,G22773,G1307);
  nand GNAME2305(G2305,G1258,G1311);
  nand GNAME2306(G2306,G1421,G1302);
  nand GNAME2307(G2307,G1260,G1309);
  nand GNAME2308(G2308,G1257,G1310);
  nand GNAME2309(G2309,G1259,G1308);
  nand GNAME2310(G2310,G1777,G1304);
  nand GNAME2311(G2311,G2310,G7092);
  nand GNAME2312(G2312,G1291,G8175);
  nand GNAME2313(G2313,G22788,G1242);
  nand GNAME2314(G2314,G1411,G1240);
  nand GNAME2315(G2315,G2314,G1312,G2313,G2311,G2312);
  nand GNAME2316(G2316,G7011,G1305);
  nand GNAME2317(G2317,G8085,G1306);
  nand GNAME2318(G2318,G2100,G22684);
  nand GNAME2319(G2319,G22778,G1307);
  nand GNAME2320(G2320,G1418,G1302);
  nand GNAME2321(G2321,G1258,G1309);
  and GNAME2322(G2322,G1633,G1241);
  or GNAME2323(G2323,G1286,G2322);
  not GNAME2324(G2324,G1625);
  or GNAME2325(G2325,G1404,G1227);
  nand GNAME2326(G2326,G2325,G1241);
  nand GNAME2327(G2327,G8084,G1314);
  nand GNAME2328(G2328,G2326,G1255);
  nand GNAME2329(G2329,G2328,G2101,G2327);
  nand GNAME2330(G2330,G8183,G1314);
  nand GNAME2331(G2331,G2326,G1256);
  nand GNAME2332(G2332,G2331,G2101,G2330);
  nand GNAME2333(G2333,G1368,G1230);
  nand GNAME2334(G2334,G2333,G1304);
  or GNAME2335(G2335,G1314,G1226);
  nand GNAME2336(G2336,G2334,G7062);
  nand GNAME2337(G2337,G2335,G8185);
  nand GNAME2338(G2338,G2114,G1235);
  nand GNAME2339(G2339,G2326,G1253);
  nand GNAME2340(G2340,G2336,G2337,G2338,G2339);
  nand GNAME2341(G2341,G2334,G7065);
  nand GNAME2342(G2342,G2335,G8186);
  nand GNAME2343(G2343,G2326,G1245);
  nand GNAME2344(G2344,G1254,G1308);
  nand GNAME2345(G2345,G1284,G1310);
  nand GNAME2346(G2346,G2344,G2345,G2343,G2341,G2342);
  nand GNAME2347(G2347,G2334,G7068);
  nand GNAME2348(G2348,G2335,G8187);
  nand GNAME2349(G2349,G2326,G1243);
  nand GNAME2350(G2350,G1283,G1310);
  nand GNAME2351(G2351,G1285,G1308);
  nand GNAME2352(G2352,G2350,G2351,G2349,G2347,G2348);
  nand GNAME2353(G2353,G2334,G7071);
  nand GNAME2354(G2354,G2335,G8188);
  nand GNAME2355(G2355,G2326,G1251);
  nand GNAME2356(G2356,G1282,G1310);
  nand GNAME2357(G2357,G1284,G1308);
  nand GNAME2358(G2358,G2356,G2357,G2355,G2353,G2354);
  nand GNAME2359(G2359,G2334,G7074);
  nand GNAME2360(G2360,G2335,G8189);
  nand GNAME2361(G2361,G2326,G1247);
  nand GNAME2362(G2362,G1281,G1310);
  nand GNAME2363(G2363,G1283,G1308);
  nand GNAME2364(G2364,G2362,G2363,G2361,G2359,G2360);
  nand GNAME2365(G2365,G2334,G7077);
  nand GNAME2366(G2366,G2335,G8190);
  nand GNAME2367(G2367,G2326,G1248);
  nand GNAME2368(G2368,G1280,G1310);
  nand GNAME2369(G2369,G1282,G1308);
  nand GNAME2370(G2370,G2368,G2369,G2367,G2365,G2366);
  nand GNAME2371(G2371,G2334,G7080);
  nand GNAME2372(G2372,G2335,G8191);
  nand GNAME2373(G2373,G2326,G1244);
  nand GNAME2374(G2374,G1279,G1310);
  nand GNAME2375(G2375,G1281,G1308);
  nand GNAME2376(G2376,G2374,G2375,G2373,G2371,G2372);
  nand GNAME2377(G2377,G2334,G7083);
  nand GNAME2378(G2378,G2335,G8192);
  nand GNAME2379(G2379,G2326,G1250);
  nand GNAME2380(G2380,G1278,G1310);
  nand GNAME2381(G2381,G1280,G1308);
  nand GNAME2382(G2382,G2380,G2381,G2379,G2377,G2378);
  nand GNAME2383(G2383,G2334,G7086);
  nand GNAME2384(G2384,G2335,G8193);
  nand GNAME2385(G2385,G2326,G1246);
  nand GNAME2386(G2386,G1277,G1310);
  nand GNAME2387(G2387,G1279,G1308);
  nand GNAME2388(G2388,G2386,G2387,G2385,G2383,G2384);
  nand GNAME2389(G2389,G2334,G7089);
  nand GNAME2390(G2390,G2335,G8194);
  nand GNAME2391(G2391,G2326,G1249);
  nand GNAME2392(G2392,G1276,G1310);
  nand GNAME2393(G2393,G1278,G1308);
  nand GNAME2394(G2394,G2392,G2393,G2391,G2389,G2390);
  nand GNAME2395(G2395,G2334,G7095);
  nand GNAME2396(G2396,G2335,G8195);
  nand GNAME2397(G2397,G2326,G1409);
  nand GNAME2398(G2398,G1275,G1310);
  nand GNAME2399(G2399,G1277,G1308);
  nand GNAME2400(G2400,G2398,G2399,G2397,G2395,G2396);
  nand GNAME2401(G2401,G2334,G7098);
  nand GNAME2402(G2402,G2335,G8196);
  nand GNAME2403(G2403,G2326,G1422);
  nand GNAME2404(G2404,G1274,G1310);
  nand GNAME2405(G2405,G1276,G1308);
  nand GNAME2406(G2406,G2404,G2405,G2403,G2401,G2402);
  nand GNAME2407(G2407,G2334,G7101);
  nand GNAME2408(G2408,G2335,G8197);
  nand GNAME2409(G2409,G2326,G1415);
  nand GNAME2410(G2410,G1273,G1310);
  nand GNAME2411(G2411,G1275,G1308);
  nand GNAME2412(G2412,G2410,G2411,G2409,G2407,G2408);
  nand GNAME2413(G2413,G2334,G7104);
  nand GNAME2414(G2414,G2335,G8198);
  nand GNAME2415(G2415,G2326,G1413);
  nand GNAME2416(G2416,G1272,G1310);
  nand GNAME2417(G2417,G1274,G1308);
  nand GNAME2418(G2418,G2416,G2417,G2415,G2413,G2414);
  nand GNAME2419(G2419,G2334,G7107);
  nand GNAME2420(G2420,G2335,G8199);
  nand GNAME2421(G2421,G2326,G1424);
  nand GNAME2422(G2422,G1271,G1310);
  nand GNAME2423(G2423,G1273,G1308);
  nand GNAME2424(G2424,G2422,G2423,G2421,G2419,G2420);
  nand GNAME2425(G2425,G2334,G7016);
  nand GNAME2426(G2426,G2335,G8200);
  nand GNAME2427(G2427,G2326,G1406);
  nand GNAME2428(G2428,G1270,G1310);
  nand GNAME2429(G2429,G1272,G1308);
  nand GNAME2430(G2430,G2428,G2429,G2427,G2425,G2426);
  nand GNAME2431(G2431,G2334,G7111);
  nand GNAME2432(G2432,G2335,G8201);
  nand GNAME2433(G2433,G2326,G1419);
  nand GNAME2434(G2434,G1269,G1310);
  nand GNAME2435(G2435,G1271,G1308);
  nand GNAME2436(G2436,G2434,G2435,G2433,G2431,G2432);
  nand GNAME2437(G2437,G2334,G7114);
  nand GNAME2438(G2438,G2335,G8202);
  nand GNAME2439(G2439,G2326,G1412);
  nand GNAME2440(G2440,G1268,G1310);
  nand GNAME2441(G2441,G1270,G1308);
  nand GNAME2442(G2442,G2440,G2441,G2439,G2437,G2438);
  nand GNAME2443(G2443,G2334,G7017);
  nand GNAME2444(G2444,G2335,G8203);
  nand GNAME2445(G2445,G2326,G1420);
  nand GNAME2446(G2446,G1267,G1310);
  nand GNAME2447(G2447,G1269,G1308);
  nand GNAME2448(G2448,G2446,G2447,G2445,G2443,G2444);
  nand GNAME2449(G2449,G2334,G6973);
  nand GNAME2450(G2450,G2335,G8204);
  nand GNAME2451(G2451,G2326,G1407);
  nand GNAME2452(G2452,G1266,G1310);
  nand GNAME2453(G2453,G1268,G1308);
  nand GNAME2454(G2454,G2452,G2453,G2451,G2449,G2450);
  nand GNAME2455(G2455,G2334,G7028);
  nand GNAME2456(G2456,G2335,G8176);
  nand GNAME2457(G2457,G2326,G1417);
  nand GNAME2458(G2458,G1265,G1310);
  nand GNAME2459(G2459,G1267,G1308);
  nand GNAME2460(G2460,G2458,G2459,G2457,G2455,G2456);
  nand GNAME2461(G2461,G2334,G7031);
  nand GNAME2462(G2462,G2335,G8177);
  nand GNAME2463(G2463,G2326,G1410);
  nand GNAME2464(G2464,G1264,G1310);
  nand GNAME2465(G2465,G1266,G1308);
  nand GNAME2466(G2466,G2464,G2465,G2463,G2461,G2462);
  nand GNAME2467(G2467,G2334,G7012);
  nand GNAME2468(G2468,G2335,G8178);
  nand GNAME2469(G2469,G2326,G1405);
  nand GNAME2470(G2470,G1263,G1310);
  nand GNAME2471(G2471,G1265,G1308);
  nand GNAME2472(G2472,G2470,G2471,G2469,G2467,G2468);
  nand GNAME2473(G2473,G2334,G6975);
  nand GNAME2474(G2474,G2335,G8179);
  nand GNAME2475(G2475,G2326,G1423);
  nand GNAME2476(G2476,G1262,G1310);
  nand GNAME2477(G2477,G1264,G1308);
  nand GNAME2478(G2478,G2476,G2477,G2475,G2473,G2474);
  nand GNAME2479(G2479,G2334,G7035);
  nand GNAME2480(G2480,G2335,G8180);
  nand GNAME2481(G2481,G2326,G1414);
  nand GNAME2482(G2482,G1261,G1310);
  nand GNAME2483(G2483,G1263,G1308);
  nand GNAME2484(G2484,G2482,G2483,G2481,G2479,G2480);
  nand GNAME2485(G2485,G2334,G7038);
  nand GNAME2486(G2486,G2335,G8181);
  nand GNAME2487(G2487,G2326,G1416);
  nand GNAME2488(G2488,G1260,G1310);
  nand GNAME2489(G2489,G1262,G1308);
  nand GNAME2490(G2490,G2488,G2489,G2487,G2485,G2486);
  nand GNAME2491(G2491,G2334,G7013);
  nand GNAME2492(G2492,G2335,G8182);
  nand GNAME2493(G2493,G2326,G1408);
  nand GNAME2494(G2494,G1259,G1310);
  nand GNAME2495(G2495,G1261,G1308);
  nand GNAME2496(G2496,G2494,G2495,G2493,G2491,G2492);
  nand GNAME2497(G2497,G2334,G6974);
  nand GNAME2498(G2498,G2335,G8184);
  nand GNAME2499(G2499,G2326,G1421);
  nand GNAME2500(G2500,G1258,G1310);
  nand GNAME2501(G2501,G1260,G1308);
  nand GNAME2502(G2502,G2500,G2501,G2499,G2497,G2498);
  nand GNAME2503(G2503,G2334,G7092);
  nand GNAME2504(G2504,G2335,G8175);
  nand GNAME2505(G2505,G2326,G1411);
  nand GNAME2506(G2506,G2503,G2504,G2505,G1312);
  nand GNAME2507(G2507,G2334,G7011);
  nand GNAME2508(G2508,G2335,G8085);
  nand GNAME2509(G2509,G2326,G1418);
  nand GNAME2510(G2510,G1258,G1308);
  nand GNAME2511(G2511,G2507,G2508,G2509,G2510);
  not GNAME2512(G2512,G1626);
  not GNAME2513(G2513,G1627);
  nand GNAME2514(G2514,G22587,G1316);
  nand GNAME2515(G2515,G7896,G1317);
  nand GNAME2516(G2516,G1066,G586);
  nand GNAME2517(G2517,G22586,G1316);
  nand GNAME2518(G2518,G1066,G587);
  nand GNAME2519(G2519,G7897,G1317);
  nand GNAME2520(G2520,G1066,G589);
  nand GNAME2521(G2521,G22585,G1316);
  nand GNAME2522(G2522,G7865,G1317);
  nand GNAME2523(G2523,G22584,G1316);
  nand GNAME2524(G2524,G7870,G1317);
  nand GNAME2525(G2525,G1066,G590);
  nand GNAME2526(G2526,G22583,G1316);
  nand GNAME2527(G2527,G7898,G1317);
  nand GNAME2528(G2528,G1066,G591);
  nand GNAME2529(G2529,G22582,G1316);
  nand GNAME2530(G2530,G7864,G1317);
  nand GNAME2531(G2531,G1066,G592);
  nand GNAME2532(G2532,G1316,G22581);
  nand GNAME2533(G2533,G1317,G7899);
  nand GNAME2534(G2534,G1066,G593);
  nand GNAME2535(G2535,G22580,G1316);
  nand GNAME2536(G2536,G7871,G1317);
  nand GNAME2537(G2537,G1066,G594);
  nand GNAME2538(G2538,G22579,G1316);
  nand GNAME2539(G2539,G7900,G1317);
  nand GNAME2540(G2540,G1066,G595);
  nand GNAME2541(G2541,G22578,G1316);
  nand GNAME2542(G2542,G7863,G1317);
  nand GNAME2543(G2543,G1066,G596);
  nand GNAME2544(G2544,G22577,G1316);
  nand GNAME2545(G2545,G7901,G1317);
  nand GNAME2546(G2546,G1066,G597);
  nand GNAME2547(G2547,G22576,G1316);
  nand GNAME2548(G2548,G7872,G1317);
  nand GNAME2549(G2549,G1066,G598);
  nand GNAME2550(G2550,G22575,G1316);
  nand GNAME2551(G2551,G7903,G1317);
  nand GNAME2552(G2552,G1066,G600);
  nand GNAME2553(G2553,G22574,G1316);
  nand GNAME2554(G2554,G7862,G1317);
  nand GNAME2555(G2555,G1066,G601);
  nand GNAME2556(G2556,G22573,G1316);
  nand GNAME2557(G2557,G7904,G1317);
  nand GNAME2558(G2558,G1066,G602);
  nand GNAME2559(G2559,G22572,G1316);
  nand GNAME2560(G2560,G7873,G1317);
  nand GNAME2561(G2561,G1066,G603);
  nand GNAME2562(G2562,G22571,G1316);
  nand GNAME2563(G2563,G7905,G1317);
  nand GNAME2564(G2564,G1066,G604);
  nand GNAME2565(G2565,G22570,G1316);
  nand GNAME2566(G2566,G7861,G1317);
  nand GNAME2567(G2567,G1066,G605);
  nand GNAME2568(G2568,G22569,G1316);
  nand GNAME2569(G2569,G7906,G1317);
  nand GNAME2570(G2570,G1066,G606);
  nand GNAME2571(G2571,G22568,G1316);
  nand GNAME2572(G2572,G7874,G1317);
  nand GNAME2573(G2573,G1066,G607);
  nand GNAME2574(G2574,G22567,G1316);
  nand GNAME2575(G2575,G7907,G1317);
  nand GNAME2576(G2576,G1066,G608);
  nand GNAME2577(G2577,G22566,G1316);
  nand GNAME2578(G2578,G7860,G1317);
  nand GNAME2579(G2579,G1066,G609);
  nand GNAME2580(G2580,G22565,G1316);
  nand GNAME2581(G2581,G7892,G1317);
  nand GNAME2582(G2582,G1066,G579);
  nand GNAME2583(G2583,G22564,G1316);
  nand GNAME2584(G2584,G7868,G1317);
  nand GNAME2585(G2585,G1066,G580);
  nand GNAME2586(G2586,G22563,G1316);
  nand GNAME2587(G2587,G7893,G1317);
  nand GNAME2588(G2588,G1066,G581);
  nand GNAME2589(G2589,G22562,G1316);
  nand GNAME2590(G2590,G7867,G1317);
  nand GNAME2591(G2591,G1066,G582);
  nand GNAME2592(G2592,G22561,G1316);
  nand GNAME2593(G2593,G7894,G1317);
  nand GNAME2594(G2594,G1066,G583);
  nand GNAME2595(G2595,G22560,G1316);
  nand GNAME2596(G2596,G7869,G1317);
  nand GNAME2597(G2597,G1066,G584);
  nand GNAME2598(G2598,G22559,G1316);
  nand GNAME2599(G2599,G7895,G1317);
  nand GNAME2600(G2600,G1066,G585);
  nand GNAME2601(G2601,G22558,G1316);
  nand GNAME2602(G2602,G7866,G1317);
  nand GNAME2603(G2603,G1066,G588);
  nand GNAME2604(G2604,G22557,G1316);
  nand GNAME2605(G2605,G7890,G1317);
  nand GNAME2606(G2606,G1066,G599);
  nand GNAME2607(G2607,G22556,G1316);
  nand GNAME2608(G2608,G22556,G1317);
  nand GNAME2609(G2609,G1066,G610);
  nand GNAME2610(G2610,G3197,G1224);
  or GNAME2611(G2611,G1215,G3605);
  or GNAME2612(G2612,G1321,G7957);
  nand GNAME2613(G2613,G1319,G2612,G2742);
  or GNAME2614(G2614,G1228,G1226);
  nand GNAME2615(G2615,G2614,G1367);
  nand GNAME2616(G2616,G1322,G1318);
  nand GNAME2617(G2617,G2616,G1417);
  nand GNAME2618(G2618,G1266,G2613);
  nand GNAME2619(G2619,G7028,G1320);
  nand GNAME2620(G2620,G1265,G1342);
  nand GNAME2621(G2621,G2616,G1410);
  nand GNAME2622(G2622,G1265,G2613);
  nand GNAME2623(G2623,G7031,G1320);
  nand GNAME2624(G2624,G1264,G1342);
  nand GNAME2625(G2625,G2616,G1405);
  nand GNAME2626(G2626,G1264,G2613);
  nand GNAME2627(G2627,G7012,G1320);
  nand GNAME2628(G2628,G1263,G1342);
  nand GNAME2629(G2629,G2616,G1423);
  nand GNAME2630(G2630,G1263,G2613);
  nand GNAME2631(G2631,G6975,G1320);
  nand GNAME2632(G2632,G1262,G1342);
  nand GNAME2633(G2633,G2616,G1414);
  nand GNAME2634(G2634,G1262,G2613);
  nand GNAME2635(G2635,G7035,G1320);
  nand GNAME2636(G2636,G1261,G1342);
  nand GNAME2637(G2637,G2616,G1416);
  nand GNAME2638(G2638,G1261,G2613);
  nand GNAME2639(G2639,G7038,G1320);
  nand GNAME2640(G2640,G1260,G1342);
  nand GNAME2641(G2641,G1320,G7014);
  nand GNAME2642(G2642,G2616,G1255);
  nand GNAME2643(G2643,G902,G2613);
  nand GNAME2644(G2644,G1320,G7015);
  nand GNAME2645(G2645,G2616,G1256);
  nand GNAME2646(G2646,G904,G2613);
  nand GNAME2647(G2647,G2616,G1408);
  nand GNAME2648(G2648,G1260,G2613);
  nand GNAME2649(G2649,G7013,G1320);
  nand GNAME2650(G2650,G1259,G1342);
  nand GNAME2651(G2651,G2616,G1253);
  nand GNAME2652(G2652,G1254,G2613);
  nand GNAME2653(G2653,G7062,G1320);
  nand GNAME2654(G2654,G1285,G1342);
  nand GNAME2655(G2655,G2616,G1245);
  nand GNAME2656(G2656,G1285,G2613);
  nand GNAME2657(G2657,G7065,G1320);
  nand GNAME2658(G2658,G1284,G1342);
  nand GNAME2659(G2659,G2616,G1243);
  nand GNAME2660(G2660,G1284,G2613);
  nand GNAME2661(G2661,G7068,G1320);
  nand GNAME2662(G2662,G1283,G1342);
  nand GNAME2663(G2663,G2616,G1251);
  nand GNAME2664(G2664,G1283,G2613);
  nand GNAME2665(G2665,G7071,G1320);
  nand GNAME2666(G2666,G1282,G1342);
  nand GNAME2667(G2667,G2616,G1247);
  nand GNAME2668(G2668,G1282,G2613);
  nand GNAME2669(G2669,G7074,G1320);
  nand GNAME2670(G2670,G1281,G1342);
  nand GNAME2671(G2671,G2616,G1248);
  nand GNAME2672(G2672,G1281,G2613);
  nand GNAME2673(G2673,G7077,G1320);
  nand GNAME2674(G2674,G1280,G1342);
  nand GNAME2675(G2675,G2616,G1244);
  nand GNAME2676(G2676,G1280,G2613);
  nand GNAME2677(G2677,G7080,G1320);
  nand GNAME2678(G2678,G1279,G1342);
  nand GNAME2679(G2679,G2616,G1250);
  nand GNAME2680(G2680,G1279,G2613);
  nand GNAME2681(G2681,G7083,G1320);
  nand GNAME2682(G2682,G1278,G1342);
  nand GNAME2683(G2683,G2616,G1246);
  nand GNAME2684(G2684,G1278,G2613);
  nand GNAME2685(G2685,G7086,G1320);
  nand GNAME2686(G2686,G1277,G1342);
  nand GNAME2687(G2687,G2616,G1249);
  nand GNAME2688(G2688,G1277,G2613);
  nand GNAME2689(G2689,G7089,G1320);
  nand GNAME2690(G2690,G1276,G1342);
  nand GNAME2691(G2691,G2616,G1421);
  nand GNAME2692(G2692,G1259,G2613);
  nand GNAME2693(G2693,G6974,G1320);
  nand GNAME2694(G2694,G1258,G1342);
  nand GNAME2695(G2695,G2616,G1409);
  nand GNAME2696(G2696,G1276,G2613);
  nand GNAME2697(G2697,G7095,G1320);
  nand GNAME2698(G2698,G1275,G1342);
  nand GNAME2699(G2699,G2616,G1422);
  nand GNAME2700(G2700,G1275,G2613);
  nand GNAME2701(G2701,G7098,G1320);
  nand GNAME2702(G2702,G1274,G1342);
  nand GNAME2703(G2703,G2616,G1415);
  nand GNAME2704(G2704,G1274,G2613);
  nand GNAME2705(G2705,G7101,G1320);
  nand GNAME2706(G2706,G1273,G1342);
  nand GNAME2707(G2707,G2616,G1413);
  nand GNAME2708(G2708,G1273,G2613);
  nand GNAME2709(G2709,G7104,G1320);
  nand GNAME2710(G2710,G1272,G1342);
  nand GNAME2711(G2711,G2616,G1424);
  nand GNAME2712(G2712,G1272,G2613);
  nand GNAME2713(G2713,G7107,G1320);
  nand GNAME2714(G2714,G1271,G1342);
  nand GNAME2715(G2715,G2616,G1406);
  nand GNAME2716(G2716,G1271,G2613);
  nand GNAME2717(G2717,G7016,G1320);
  nand GNAME2718(G2718,G1270,G1342);
  nand GNAME2719(G2719,G2616,G1419);
  nand GNAME2720(G2720,G1270,G2613);
  nand GNAME2721(G2721,G7111,G1320);
  nand GNAME2722(G2722,G1269,G1342);
  nand GNAME2723(G2723,G2616,G1412);
  nand GNAME2724(G2724,G1269,G2613);
  nand GNAME2725(G2725,G7114,G1320);
  nand GNAME2726(G2726,G1268,G1342);
  nand GNAME2727(G2727,G2616,G1420);
  nand GNAME2728(G2728,G1268,G2613);
  nand GNAME2729(G2729,G7017,G1320);
  nand GNAME2730(G2730,G1267,G1342);
  nand GNAME2731(G2731,G2616,G1407);
  nand GNAME2732(G2732,G1267,G2613);
  nand GNAME2733(G2733,G6973,G1320);
  nand GNAME2734(G2734,G1266,G1342);
  nand GNAME2735(G2735,G2616,G1411);
  nand GNAME2736(G2736,G1258,G2613);
  nand GNAME2737(G2737,G7092,G1320);
  nand GNAME2738(G2738,G1257,G1342);
  nand GNAME2739(G2739,G2616,G1418);
  nand GNAME2740(G2740,G1257,G2613);
  nand GNAME2741(G2741,G7011,G1320);
  or GNAME2742(G2742,G1404,G1629);
  or GNAME2743(G2743,G7957,G1322);
  nand GNAME2744(G2744,G2743,G1318);
  nand GNAME2745(G2745,G1319,G1321);
  nand GNAME2746(G2746,G2745,G1417);
  nand GNAME2747(G2747,G1266,G2744);
  nand GNAME2748(G2748,G7028,G1323);
  nand GNAME2749(G2749,G2745,G1410);
  nand GNAME2750(G2750,G1265,G2744);
  nand GNAME2751(G2751,G7031,G1323);
  nand GNAME2752(G2752,G2745,G1405);
  nand GNAME2753(G2753,G1264,G2744);
  nand GNAME2754(G2754,G7012,G1323);
  nand GNAME2755(G2755,G2745,G1423);
  nand GNAME2756(G2756,G1263,G2744);
  nand GNAME2757(G2757,G6975,G1323);
  nand GNAME2758(G2758,G2745,G1414);
  nand GNAME2759(G2759,G1262,G2744);
  nand GNAME2760(G2760,G7035,G1323);
  nand GNAME2761(G2761,G2745,G1416);
  nand GNAME2762(G2762,G1261,G2744);
  nand GNAME2763(G2763,G7038,G1323);
  nand GNAME2764(G2764,G2745,G1255);
  nand GNAME2765(G2765,G902,G2744);
  nand GNAME2766(G2766,G7014,G1323);
  nand GNAME2767(G2767,G2745,G1256);
  nand GNAME2768(G2768,G904,G2744);
  nand GNAME2769(G2769,G7015,G1323);
  nand GNAME2770(G2770,G2745,G1408);
  nand GNAME2771(G2771,G1260,G2744);
  nand GNAME2772(G2772,G7013,G1323);
  nand GNAME2773(G2773,G2745,G1253);
  nand GNAME2774(G2774,G1254,G2744);
  nand GNAME2775(G2775,G7062,G1323);
  nand GNAME2776(G2776,G2745,G1245);
  nand GNAME2777(G2777,G1285,G2744);
  nand GNAME2778(G2778,G7065,G1323);
  nand GNAME2779(G2779,G2745,G1243);
  nand GNAME2780(G2780,G1284,G2744);
  nand GNAME2781(G2781,G7068,G1323);
  nand GNAME2782(G2782,G2745,G1251);
  nand GNAME2783(G2783,G1283,G2744);
  nand GNAME2784(G2784,G7071,G1323);
  nand GNAME2785(G2785,G2745,G1247);
  nand GNAME2786(G2786,G1282,G2744);
  nand GNAME2787(G2787,G7074,G1323);
  nand GNAME2788(G2788,G2745,G1248);
  nand GNAME2789(G2789,G1281,G2744);
  nand GNAME2790(G2790,G7077,G1323);
  nand GNAME2791(G2791,G2745,G1244);
  nand GNAME2792(G2792,G1280,G2744);
  nand GNAME2793(G2793,G7080,G1323);
  nand GNAME2794(G2794,G2745,G1250);
  nand GNAME2795(G2795,G1279,G2744);
  nand GNAME2796(G2796,G7083,G1323);
  nand GNAME2797(G2797,G2745,G1246);
  nand GNAME2798(G2798,G1278,G2744);
  nand GNAME2799(G2799,G7086,G1323);
  nand GNAME2800(G2800,G2745,G1249);
  nand GNAME2801(G2801,G1277,G2744);
  nand GNAME2802(G2802,G7089,G1323);
  nand GNAME2803(G2803,G2745,G1421);
  nand GNAME2804(G2804,G1259,G2744);
  nand GNAME2805(G2805,G6974,G1323);
  nand GNAME2806(G2806,G2745,G1409);
  nand GNAME2807(G2807,G1276,G2744);
  nand GNAME2808(G2808,G7095,G1323);
  nand GNAME2809(G2809,G2745,G1422);
  nand GNAME2810(G2810,G1275,G2744);
  nand GNAME2811(G2811,G7098,G1323);
  nand GNAME2812(G2812,G2745,G1415);
  nand GNAME2813(G2813,G1274,G2744);
  nand GNAME2814(G2814,G7101,G1323);
  nand GNAME2815(G2815,G2745,G1413);
  nand GNAME2816(G2816,G1273,G2744);
  nand GNAME2817(G2817,G7104,G1323);
  nand GNAME2818(G2818,G2745,G1424);
  nand GNAME2819(G2819,G1272,G2744);
  nand GNAME2820(G2820,G7107,G1323);
  nand GNAME2821(G2821,G2745,G1406);
  nand GNAME2822(G2822,G1271,G2744);
  nand GNAME2823(G2823,G7016,G1323);
  nand GNAME2824(G2824,G2745,G1419);
  nand GNAME2825(G2825,G1270,G2744);
  nand GNAME2826(G2826,G7111,G1323);
  nand GNAME2827(G2827,G2745,G1412);
  nand GNAME2828(G2828,G1269,G2744);
  nand GNAME2829(G2829,G7114,G1323);
  nand GNAME2830(G2830,G2745,G1420);
  nand GNAME2831(G2831,G1268,G2744);
  nand GNAME2832(G2832,G7017,G1323);
  nand GNAME2833(G2833,G2745,G1407);
  nand GNAME2834(G2834,G1267,G2744);
  nand GNAME2835(G2835,G6973,G1323);
  nand GNAME2836(G2836,G2745,G1411);
  nand GNAME2837(G2837,G1258,G2744);
  nand GNAME2838(G2838,G7092,G1323);
  nand GNAME2839(G2839,G2745,G1418);
  nand GNAME2840(G2840,G1257,G2744);
  nand GNAME2841(G2841,G7011,G1323);
  or GNAME2842(G2842,G1315,G1341);
  and GNAME2843(G2843,G1328,G1218);
  nand GNAME2844(G2844,G1367,G1325);
  nand GNAME2845(G2845,G1218,G1285,G1328);
  nand GNAME2846(G2846,G1254,G1326);
  nand GNAME2847(G2847,G902,G3115);
  nand GNAME2848(G2848,G904,G3115);
  nand GNAME2849(G2849,G1254,G3115);
  nand GNAME2850(G2850,G1403,G1218);
  nand GNAME2851(G2851,G1325,G1631,G2850);
  or GNAME2852(G2852,G1403,G1328);
  nand GNAME2853(G2853,G1245,G2852,G1218);
  nand GNAME2854(G2854,G1253,G1326);
  nand GNAME2855(G2855,G1255,G1329);
  nand GNAME2856(G2856,G1256,G1329);
  nand GNAME2857(G2857,G1253,G1329);
  nand GNAME2858(G2858,G2842,G1333);
  nand GNAME2859(G2859,G1315,G1331);
  and GNAME2860(G2860,G1218,G1333);
  or GNAME2861(G2861,G3062,G1335);
  or GNAME2862(G2862,G3115,G1231);
  nand GNAME2863(G2863,G2862,G3605,G1777);
  and GNAME2864(G2864,G1634,G2863);
  or GNAME2865(G2865,G2864,G1331);
  nand GNAME2866(G2866,G2863,G1634,G2842);
  nand GNAME2867(G2867,G1341,G1331);
  or GNAME2868(G2868,G1338,G1332);
  nand GNAME2869(G2869,G2868,G1417);
  nand GNAME2870(G2870,G1266,G2861);
  nand GNAME2871(G2871,G22661,G1336);
  nand GNAME2872(G2872,G22693,G1337);
  nand GNAME2873(G2873,G2868,G1410);
  nand GNAME2874(G2874,G1265,G2861);
  nand GNAME2875(G2875,G22660,G1336);
  nand GNAME2876(G2876,G22692,G1337);
  nand GNAME2877(G2877,G2868,G1405);
  nand GNAME2878(G2878,G1264,G2861);
  nand GNAME2879(G2879,G22659,G1336);
  nand GNAME2880(G2880,G22691,G1337);
  nand GNAME2881(G2881,G2868,G1423);
  nand GNAME2882(G2882,G1263,G2861);
  nand GNAME2883(G2883,G22658,G1336);
  nand GNAME2884(G2884,G22690,G1337);
  nand GNAME2885(G2885,G2868,G1414);
  nand GNAME2886(G2886,G1262,G2861);
  nand GNAME2887(G2887,G22657,G1336);
  nand GNAME2888(G2888,G22689,G1337);
  nand GNAME2889(G2889,G2868,G1416);
  nand GNAME2890(G2890,G1261,G2861);
  nand GNAME2891(G2891,G22656,G1336);
  nand GNAME2892(G2892,G22688,G1337);
  nand GNAME2893(G2893,G22703,G1337);
  nand GNAME2894(G2894,G22671,G1336);
  nand GNAME2895(G2895,G1333,G1285,G1218);
  nand GNAME2896(G2896,G1334,G1254);
  nand GNAME2897(G2897,G1332,G1253);
  nand GNAME2898(G2898,G1245,G1338);
  nand GNAME2899(G2899,G902,G3062);
  nand GNAME2900(G2900,G904,G3062);
  nand GNAME2901(G2901,G2868,G1408);
  nand GNAME2902(G2902,G1260,G2861);
  nand GNAME2903(G2903,G22655,G1336);
  nand GNAME2904(G2904,G22687,G1337);
  nand GNAME2905(G2905,G1254,G3062);
  nand GNAME2906(G2906,G2868,G1245);
  nand GNAME2907(G2907,G1285,G2861);
  nand GNAME2908(G2908,G2868,G1243);
  nand GNAME2909(G2909,G1284,G2861);
  nand GNAME2910(G2910,G2868,G1251);
  nand GNAME2911(G2911,G1283,G2861);
  nand GNAME2912(G2912,G2868,G1247);
  nand GNAME2913(G2913,G1282,G2861);
  nand GNAME2914(G2914,G2868,G1248);
  nand GNAME2915(G2915,G1281,G2861);
  nand GNAME2916(G2916,G2868,G1244);
  nand GNAME2917(G2917,G1280,G2861);
  nand GNAME2918(G2918,G2868,G1250);
  nand GNAME2919(G2919,G1279,G2861);
  nand GNAME2920(G2920,G2868,G1246);
  nand GNAME2921(G2921,G1278,G2861);
  nand GNAME2922(G2922,G2868,G1249);
  nand GNAME2923(G2923,G1277,G2861);
  nand GNAME2924(G2924,G2868,G1421);
  nand GNAME2925(G2925,G1259,G2861);
  nand GNAME2926(G2926,G22654,G1336);
  nand GNAME2927(G2927,G22686,G1337);
  nand GNAME2928(G2928,G2868,G1409);
  nand GNAME2929(G2929,G1276,G2861);
  nand GNAME2930(G2930,G2868,G1422);
  nand GNAME2931(G2931,G1275,G2861);
  nand GNAME2932(G2932,G22670,G1336);
  nand GNAME2933(G2933,G22702,G1337);
  nand GNAME2934(G2934,G2868,G1415);
  nand GNAME2935(G2935,G1274,G2861);
  nand GNAME2936(G2936,G22669,G1336);
  nand GNAME2937(G2937,G22701,G1337);
  nand GNAME2938(G2938,G2868,G1413);
  nand GNAME2939(G2939,G1273,G2861);
  nand GNAME2940(G2940,G22668,G1336);
  nand GNAME2941(G2941,G22700,G1337);
  nand GNAME2942(G2942,G2868,G1424);
  nand GNAME2943(G2943,G1272,G2861);
  nand GNAME2944(G2944,G22667,G1336);
  nand GNAME2945(G2945,G22699,G1337);
  nand GNAME2946(G2946,G2868,G1406);
  nand GNAME2947(G2947,G1271,G2861);
  nand GNAME2948(G2948,G22666,G1336);
  nand GNAME2949(G2949,G22698,G1337);
  nand GNAME2950(G2950,G2868,G1419);
  nand GNAME2951(G2951,G1270,G2861);
  nand GNAME2952(G2952,G22665,G1336);
  nand GNAME2953(G2953,G22697,G1337);
  nand GNAME2954(G2954,G2868,G1412);
  nand GNAME2955(G2955,G1269,G2861);
  nand GNAME2956(G2956,G22664,G1336);
  nand GNAME2957(G2957,G22696,G1337);
  nand GNAME2958(G2958,G2868,G1420);
  nand GNAME2959(G2959,G1268,G2861);
  nand GNAME2960(G2960,G22663,G1336);
  nand GNAME2961(G2961,G22695,G1337);
  nand GNAME2962(G2962,G2868,G1407);
  nand GNAME2963(G2963,G1267,G2861);
  nand GNAME2964(G2964,G22662,G1336);
  nand GNAME2965(G2965,G22694,G1337);
  nand GNAME2966(G2966,G2868,G1411);
  nand GNAME2967(G2967,G1258,G2861);
  nand GNAME2968(G2968,G22653,G1336);
  nand GNAME2969(G2969,G22685,G1337);
  nand GNAME2970(G2970,G2868,G1418);
  nand GNAME2971(G2971,G1257,G2861);
  nand GNAME2972(G2972,G22652,G1336);
  nand GNAME2973(G2973,G22684,G1337);
  nand GNAME2974(G2974,G1364,G1211);
  or GNAME2975(G2975,G1337,G1336);
  nand GNAME2976(G2976,G1266,G2868);
  nand GNAME2977(G2977,G2975,G1346);
  nand GNAME2978(G2978,G1335,G1417);
  nand GNAME2979(G2979,G1265,G2868);
  nand GNAME2980(G2980,G2975,G1347);
  nand GNAME2981(G2981,G1335,G1410);
  nand GNAME2982(G2982,G1264,G2868);
  nand GNAME2983(G2983,G2975,G1348);
  nand GNAME2984(G2984,G1335,G1405);
  nand GNAME2985(G2985,G1263,G2868);
  nand GNAME2986(G2986,G2975,G1349);
  nand GNAME2987(G2987,G1335,G1423);
  nand GNAME2988(G2988,G1262,G2868);
  nand GNAME2989(G2989,G2975,G1350);
  nand GNAME2990(G2990,G1335,G1414);
  nand GNAME2991(G2991,G1261,G2868);
  nand GNAME2992(G2992,G2975,G1351);
  nand GNAME2993(G2993,G1335,G1416);
  nand GNAME2994(G2994,G2975,G3200);
  nand GNAME2995(G2995,G1333,G1218,G1245);
  nand GNAME2996(G2996,G1334,G1253);
  nand GNAME2997(G2997,G1254,G1332);
  nand GNAME2998(G2998,G1285,G1338);
  nand GNAME2999(G2999,G1260,G2868);
  nand GNAME3000(G3000,G2975,G1352);
  nand GNAME3001(G3001,G1335,G1408);
  nand GNAME3002(G3002,G1285,G2868);
  nand GNAME3003(G3003,G1335,G1245);
  nand GNAME3004(G3004,G1284,G2868);
  nand GNAME3005(G3005,G1335,G1243);
  nand GNAME3006(G3006,G1283,G2868);
  nand GNAME3007(G3007,G1335,G1251);
  nand GNAME3008(G3008,G1282,G2868);
  nand GNAME3009(G3009,G1335,G1247);
  nand GNAME3010(G3010,G1281,G2868);
  nand GNAME3011(G3011,G1335,G1248);
  nand GNAME3012(G3012,G1280,G2868);
  nand GNAME3013(G3013,G1335,G1244);
  nand GNAME3014(G3014,G1279,G2868);
  nand GNAME3015(G3015,G1335,G1250);
  nand GNAME3016(G3016,G1278,G2868);
  nand GNAME3017(G3017,G1335,G1246);
  nand GNAME3018(G3018,G1277,G2868);
  nand GNAME3019(G3019,G1335,G1249);
  nand GNAME3020(G3020,G1259,G2868);
  nand GNAME3021(G3021,G2975,G1353);
  nand GNAME3022(G3022,G1335,G1421);
  nand GNAME3023(G3023,G1276,G2868);
  nand GNAME3024(G3024,G1335,G1409);
  nand GNAME3025(G3025,G1275,G2868);
  nand GNAME3026(G3026,G2975,G1355);
  nand GNAME3027(G3027,G1335,G1422);
  nand GNAME3028(G3028,G1274,G2868);
  nand GNAME3029(G3029,G2975,G1356);
  nand GNAME3030(G3030,G1335,G1415);
  nand GNAME3031(G3031,G1273,G2868);
  nand GNAME3032(G3032,G2975,G1357);
  nand GNAME3033(G3033,G1335,G1413);
  nand GNAME3034(G3034,G1272,G2868);
  nand GNAME3035(G3035,G2975,G1358);
  nand GNAME3036(G3036,G1335,G1424);
  nand GNAME3037(G3037,G1271,G2868);
  nand GNAME3038(G3038,G2975,G1359);
  nand GNAME3039(G3039,G1335,G1406);
  nand GNAME3040(G3040,G1270,G2868);
  nand GNAME3041(G3041,G2975,G1360);
  nand GNAME3042(G3042,G1335,G1419);
  nand GNAME3043(G3043,G1269,G2868);
  nand GNAME3044(G3044,G2975,G1361);
  nand GNAME3045(G3045,G1335,G1412);
  nand GNAME3046(G3046,G1268,G2868);
  nand GNAME3047(G3047,G2975,G1362);
  nand GNAME3048(G3048,G1335,G1420);
  nand GNAME3049(G3049,G1267,G2868);
  nand GNAME3050(G3050,G2975,G1363);
  nand GNAME3051(G3051,G1335,G1407);
  nand GNAME3052(G3052,G1258,G2868);
  nand GNAME3053(G3053,G2975,G1354);
  nand GNAME3054(G3054,G1335,G1411);
  nand GNAME3055(G3055,G1257,G2868);
  nand GNAME3056(G3056,G2975,G1364);
  nand GNAME3057(G3057,G1544,G1211);
  nand GNAME3058(G3058,G1335,G1418);
  nand GNAME3059(G3059,G1300,G22716);
  nand GNAME3060(G3060,G1621,G22579);
  nand GNAME3061(G3061,G7900,G22587);
  not GNAME3062(G3062,G1342);
  or GNAME3063(G3063,G7899,G1621);
  or GNAME3064(G3064,G22581,G22587);
  nand GNAME3065(G3065,G1621,G22582);
  nand GNAME3066(G3066,G7864,G22587);
  nand GNAME3067(G3067,G1621,G22580);
  nand GNAME3068(G3068,G7871,G22587);
  nand GNAME3069(G3069,G1621,G22565);
  nand GNAME3070(G3070,G7892,G22587);
  nand GNAME3071(G3071,G1621,G22564);
  nand GNAME3072(G3072,G7868,G22587);
  nand GNAME3073(G3073,G1621,G22563);
  nand GNAME3074(G3074,G7893,G22587);
  nand GNAME3075(G3075,G1621,G22562);
  nand GNAME3076(G3076,G7867,G22587);
  nand GNAME3077(G3077,G1621,G22561);
  nand GNAME3078(G3078,G7894,G22587);
  nand GNAME3079(G3079,G1621,G22560);
  nand GNAME3080(G3080,G7869,G22587);
  nand GNAME3081(G3081,G1621,G22559);
  nand GNAME3082(G3082,G7895,G22587);
  nand GNAME3083(G3083,G1621,G22558);
  nand GNAME3084(G3084,G7866,G22587);
  nand GNAME3085(G3085,G1621,G22557);
  nand GNAME3086(G3086,G7890,G22587);
  nand GNAME3087(G3087,G1621,G22574);
  nand GNAME3088(G3088,G7862,G22587);
  nand GNAME3089(G3089,G1621,G22573);
  nand GNAME3090(G3090,G7904,G22587);
  nand GNAME3091(G3091,G1621,G22572);
  nand GNAME3092(G3092,G7873,G22587);
  nand GNAME3093(G3093,G1621,G22571);
  nand GNAME3094(G3094,G7905,G22587);
  nand GNAME3095(G3095,G1621,G22570);
  nand GNAME3096(G3096,G7861,G22587);
  nand GNAME3097(G3097,G1621,G22569);
  nand GNAME3098(G3098,G7906,G22587);
  nand GNAME3099(G3099,G1621,G22568);
  nand GNAME3100(G3100,G7874,G22587);
  nand GNAME3101(G3101,G1621,G22567);
  nand GNAME3102(G3102,G7907,G22587);
  nand GNAME3103(G3103,G1621,G22566);
  nand GNAME3104(G3104,G7860,G22587);
  nand GNAME3105(G3105,G1621,G22556);
  nand GNAME3106(G3106,G22556,G22587);
  nand GNAME3107(G3107,G1621,G22583);
  nand GNAME3108(G3108,G7898,G22587);
  not GNAME3109(G3109,G1365);
  nand GNAME3110(G3110,G1621,G22584);
  nand GNAME3111(G3111,G7870,G22587);
  not GNAME3112(G3112,G1366);
  nand GNAME3113(G3113,G1621,G22577);
  nand GNAME3114(G3114,G7901,G22587);
  not GNAME3115(G3115,G1367);
  nand GNAME3116(G3116,G1621,G22578);
  nand GNAME3117(G3117,G7863,G22587);
  not GNAME3118(G3118,G1368);
  or GNAME3119(G3119,G22587,G22586,G1213);
  or GNAME3120(G3120,G1621,G7897,G1212);
  nand GNAME3121(G3121,G3119,G3120);
  nand GNAME3122(G3122,G1621,G1213,G22586);
  or GNAME3123(G3123,G1621,G7865,G1214);
  nand GNAME3124(G3124,G3122,G3123);
  nand GNAME3125(G3125,G1621,G22585,G22586);
  or GNAME3126(G3126,G1621,G1212,G1214);
  nand GNAME3127(G3127,G3125,G3126);
  or GNAME3128(G3128,G22587,G22586,G22585);
  or GNAME3129(G3129,G1621,G7897,G7865);
  nand GNAME3130(G3130,G3128,G3129);
  nand GNAME3131(G3131,G1622,G8176);
  nand GNAME3132(G3132,G1266,G7729);
  nand GNAME3133(G3133,G1622,G8177);
  nand GNAME3134(G3134,G1265,G7729);
  nand GNAME3135(G3135,G1622,G8178);
  nand GNAME3136(G3136,G1264,G7729);
  nand GNAME3137(G3137,G1622,G8179);
  nand GNAME3138(G3138,G1263,G7729);
  nand GNAME3139(G3139,G1622,G8180);
  nand GNAME3140(G3140,G1262,G7729);
  nand GNAME3141(G3141,G1622,G8181);
  nand GNAME3142(G3142,G1261,G7729);
  nand GNAME3143(G3143,G1622,G8182);
  nand GNAME3144(G3144,G1260,G7729);
  nand GNAME3145(G3145,G1622,G8084);
  nand GNAME3146(G3146,G902,G7729);
  nand GNAME3147(G3147,G1622,G8183);
  nand GNAME3148(G3148,G904,G7729);
  nand GNAME3149(G3149,G1622,G8184);
  nand GNAME3150(G3150,G1259,G7729);
  nand GNAME3151(G3151,G1622,G8185);
  nand GNAME3152(G3152,G1254,G7729);
  nand GNAME3153(G3153,G1622,G8186);
  nand GNAME3154(G3154,G1285,G7729);
  nand GNAME3155(G3155,G1622,G8187);
  nand GNAME3156(G3156,G1284,G7729);
  nand GNAME3157(G3157,G1622,G8188);
  nand GNAME3158(G3158,G1283,G7729);
  nand GNAME3159(G3159,G1622,G8189);
  nand GNAME3160(G3160,G1282,G7729);
  nand GNAME3161(G3161,G1622,G8190);
  nand GNAME3162(G3162,G1281,G7729);
  nand GNAME3163(G3163,G1622,G8191);
  nand GNAME3164(G3164,G1280,G7729);
  nand GNAME3165(G3165,G1622,G8192);
  nand GNAME3166(G3166,G1279,G7729);
  nand GNAME3167(G3167,G1622,G8193);
  nand GNAME3168(G3168,G1278,G7729);
  nand GNAME3169(G3169,G1622,G8194);
  nand GNAME3170(G3170,G1277,G7729);
  nand GNAME3171(G3171,G1622,G8175);
  nand GNAME3172(G3172,G1258,G7729);
  nand GNAME3173(G3173,G1622,G8195);
  nand GNAME3174(G3174,G1276,G7729);
  nand GNAME3175(G3175,G1622,G8196);
  nand GNAME3176(G3176,G1275,G7729);
  nand GNAME3177(G3177,G1622,G8197);
  nand GNAME3178(G3178,G1274,G7729);
  nand GNAME3179(G3179,G1622,G8198);
  nand GNAME3180(G3180,G1273,G7729);
  nand GNAME3181(G3181,G1622,G8199);
  nand GNAME3182(G3182,G1272,G7729);
  nand GNAME3183(G3183,G1622,G8200);
  nand GNAME3184(G3184,G1271,G7729);
  nand GNAME3185(G3185,G1622,G8201);
  nand GNAME3186(G3186,G1270,G7729);
  nand GNAME3187(G3187,G1622,G8202);
  nand GNAME3188(G3188,G1269,G7729);
  nand GNAME3189(G3189,G1622,G8203);
  nand GNAME3190(G3190,G1268,G7729);
  nand GNAME3191(G3191,G1622,G8204);
  nand GNAME3192(G3192,G1267,G7729);
  nand GNAME3193(G3193,G1622,G8085);
  nand GNAME3194(G3194,G1257,G7729);
  nand GNAME3195(G3195,G1621,G22576);
  nand GNAME3196(G3196,G7872,G22587);
  not GNAME3197(G3197,G1404);
  nand GNAME3198(G3198,G1621,G22575);
  nand GNAME3199(G3199,G7903,G22587);
  not GNAME3200(G3200,G1403);
  nand GNAME3201(G3201,G22768,G1344);
  or GNAME3202(G3202,G22768,G1344);
  nand GNAME3203(G3203,G3201,G3202);
  nand GNAME3204(G3204,G1217,G22588);
  nand GNAME3205(G3205,G1767,G1771);
  not GNAME3206(G3206,G1401);
  nand GNAME3207(G3207,G1217,G22589);
  nand GNAME3208(G3208,G1767,G1772);
  not GNAME3209(G3209,G1402);
  nand GNAME3210(G3210,G1632,G581);
  nand GNAME3211(G3211,G1348,G1623);
  nand GNAME3212(G3212,G1632,G605);
  nand GNAME3213(G3213,G1359,G1623);
  nand GNAME3214(G3214,G1632,G609);
  nand GNAME3215(G3215,G1363,G1623);
  nand GNAME3216(G3216,G1632,G585);
  nand GNAME3217(G3217,G1352,G1623);
  nand GNAME3218(G3218,G1632,G600);
  or GNAME3219(G3219,G1403,G1632);
  nand GNAME3220(G3220,G1632,G580);
  nand GNAME3221(G3221,G1347,G1623);
  nand GNAME3222(G3222,G1632,G599);
  nand GNAME3223(G3223,G1354,G1623);
  nand GNAME3224(G3224,G1632,G607);
  nand GNAME3225(G3225,G1361,G1623);
  nand GNAME3226(G3226,G1632,G603);
  nand GNAME3227(G3227,G1357,G1623);
  nand GNAME3228(G3228,G1632,G583);
  nand GNAME3229(G3229,G1350,G1623);
  nand GNAME3230(G3230,G1632,G602);
  nand GNAME3231(G3231,G1356,G1623);
  nand GNAME3232(G3232,G1632,G584);
  nand GNAME3233(G3233,G1351,G1623);
  nand GNAME3234(G3234,G1632,G579);
  nand GNAME3235(G3235,G1346,G1623);
  nand GNAME3236(G3236,G1632,G610);
  nand GNAME3237(G3237,G1364,G1623);
  nand GNAME3238(G3238,G1632,G606);
  nand GNAME3239(G3239,G1360,G1623);
  nand GNAME3240(G3240,G1632,G608);
  nand GNAME3241(G3241,G1362,G1623);
  nand GNAME3242(G3242,G1632,G588);
  nand GNAME3243(G3243,G1353,G1623);
  nand GNAME3244(G3244,G1632,G601);
  nand GNAME3245(G3245,G1355,G1623);
  nand GNAME3246(G3246,G1632,G582);
  nand GNAME3247(G3247,G1349,G1623);
  nand GNAME3248(G3248,G1632,G604);
  nand GNAME3249(G3249,G1358,G1623);
  or GNAME3250(G3250,G3115,G1622);
  or GNAME3251(G3251,G7729,G1367);
  nand GNAME3252(G3252,G3250,G3251);
  nand GNAME3253(G3253,G1254,G1253);
  or GNAME3254(G3254,G1253,G1254);
  nand GNAME3255(G3255,G3253,G3254);
  nand GNAME3256(G3256,G902,G1255);
  or GNAME3257(G3257,G902,G1255);
  nand GNAME3258(G3258,G3256,G3257);
  nand GNAME3259(G3259,G904,G1256);
  or GNAME3260(G3260,G904,G1256);
  nand GNAME3261(G3261,G3259,G3260);
  or GNAME3262(G3262,G1257,G1418);
  nand GNAME3263(G3263,G1257,G1418);
  nand GNAME3264(G3264,G3262,G3263);
  or GNAME3265(G3265,G1258,G1411);
  nand GNAME3266(G3266,G1258,G1411);
  nand GNAME3267(G3267,G3265,G3266);
  or GNAME3268(G3268,G1259,G1421);
  nand GNAME3269(G3269,G1259,G1421);
  nand GNAME3270(G3270,G3268,G3269);
  or GNAME3271(G3271,G1260,G1408);
  nand GNAME3272(G3272,G1260,G1408);
  nand GNAME3273(G3273,G3271,G3272);
  or GNAME3274(G3274,G1261,G1416);
  nand GNAME3275(G3275,G1261,G1416);
  nand GNAME3276(G3276,G3274,G3275);
  or GNAME3277(G3277,G1262,G1414);
  nand GNAME3278(G3278,G1262,G1414);
  nand GNAME3279(G3279,G3277,G3278);
  or GNAME3280(G3280,G1263,G1423);
  nand GNAME3281(G3281,G1263,G1423);
  nand GNAME3282(G3282,G3280,G3281);
  or GNAME3283(G3283,G1264,G1405);
  nand GNAME3284(G3284,G1264,G1405);
  nand GNAME3285(G3285,G3283,G3284);
  or GNAME3286(G3286,G1265,G1410);
  nand GNAME3287(G3287,G1265,G1410);
  nand GNAME3288(G3288,G3286,G3287);
  or GNAME3289(G3289,G1266,G1417);
  nand GNAME3290(G3290,G1266,G1417);
  nand GNAME3291(G3291,G3289,G3290);
  or GNAME3292(G3292,G1267,G1407);
  nand GNAME3293(G3293,G1267,G1407);
  nand GNAME3294(G3294,G3292,G3293);
  or GNAME3295(G3295,G1268,G1420);
  nand GNAME3296(G3296,G1268,G1420);
  nand GNAME3297(G3297,G3295,G3296);
  or GNAME3298(G3298,G1269,G1412);
  nand GNAME3299(G3299,G1269,G1412);
  nand GNAME3300(G3300,G3298,G3299);
  or GNAME3301(G3301,G1270,G1419);
  nand GNAME3302(G3302,G1270,G1419);
  nand GNAME3303(G3303,G3301,G3302);
  or GNAME3304(G3304,G1271,G1406);
  nand GNAME3305(G3305,G1271,G1406);
  nand GNAME3306(G3306,G3304,G3305);
  or GNAME3307(G3307,G1272,G1424);
  nand GNAME3308(G3308,G1272,G1424);
  nand GNAME3309(G3309,G3307,G3308);
  or GNAME3310(G3310,G1273,G1413);
  nand GNAME3311(G3311,G1273,G1413);
  nand GNAME3312(G3312,G3310,G3311);
  or GNAME3313(G3313,G1274,G1415);
  nand GNAME3314(G3314,G1274,G1415);
  nand GNAME3315(G3315,G3313,G3314);
  or GNAME3316(G3316,G1275,G1422);
  nand GNAME3317(G3317,G1275,G1422);
  nand GNAME3318(G3318,G3316,G3317);
  nand GNAME3319(G3319,G1277,G1249);
  or GNAME3320(G3320,G1249,G1277);
  nand GNAME3321(G3321,G3319,G3320);
  or GNAME3322(G3322,G1276,G1409);
  nand GNAME3323(G3323,G1276,G1409);
  nand GNAME3324(G3324,G3322,G3323);
  nand GNAME3325(G3325,G1278,G1246);
  or GNAME3326(G3326,G1246,G1278);
  nand GNAME3327(G3327,G3325,G3326);
  nand GNAME3328(G3328,G1279,G1250);
  or GNAME3329(G3329,G1250,G1279);
  nand GNAME3330(G3330,G3328,G3329);
  nand GNAME3331(G3331,G1280,G1244);
  or GNAME3332(G3332,G1244,G1280);
  nand GNAME3333(G3333,G3331,G3332);
  nand GNAME3334(G3334,G1281,G1248);
  or GNAME3335(G3335,G1248,G1281);
  nand GNAME3336(G3336,G3334,G3335);
  nand GNAME3337(G3337,G1282,G1247);
  or GNAME3338(G3338,G1247,G1282);
  nand GNAME3339(G3339,G3337,G3338);
  nand GNAME3340(G3340,G1283,G1251);
  or GNAME3341(G3341,G1251,G1283);
  nand GNAME3342(G3342,G3340,G3341);
  nand GNAME3343(G3343,G1284,G1243);
  or GNAME3344(G3344,G1243,G1284);
  nand GNAME3345(G3345,G3343,G3344);
  nand GNAME3346(G3346,G1285,G1245);
  or GNAME3347(G3347,G1245,G1285);
  nand GNAME3348(G3348,G3346,G3347);
  nand GNAME3349(G3349,G1973,G7729);
  or GNAME3350(G3350,G7729,G1368,G3115,G3197);
  or GNAME3351(G3351,G1252,G3062);
  or GNAME3352(G3352,G1342,G1368);
  nand GNAME3353(G3353,G1630,G22767);
  nand GNAME3354(G3354,G902,G1290);
  nand GNAME3355(G3355,G1630,G22766);
  nand GNAME3356(G3356,G904,G1290);
  nand GNAME3357(G3357,G1630,G22765);
  nand GNAME3358(G3358,G1254,G1290);
  nand GNAME3359(G3359,G1630,G22764);
  nand GNAME3360(G3360,G1285,G1290);
  nand GNAME3361(G3361,G1630,G22763);
  nand GNAME3362(G3362,G1284,G1290);
  nand GNAME3363(G3363,G1630,G22762);
  nand GNAME3364(G3364,G1283,G1290);
  nand GNAME3365(G3365,G1630,G22761);
  nand GNAME3366(G3366,G1282,G1290);
  nand GNAME3367(G3367,G1630,G22760);
  nand GNAME3368(G3368,G1281,G1290);
  nand GNAME3369(G3369,G1630,G22759);
  nand GNAME3370(G3370,G1280,G1290);
  nand GNAME3371(G3371,G1630,G22758);
  nand GNAME3372(G3372,G1279,G1290);
  nand GNAME3373(G3373,G1630,G22757);
  nand GNAME3374(G3374,G1278,G1290);
  nand GNAME3375(G3375,G1630,G22756);
  nand GNAME3376(G3376,G1277,G1290);
  nand GNAME3377(G3377,G1630,G22755);
  nand GNAME3378(G3378,G1276,G1290);
  nand GNAME3379(G3379,G1630,G22754);
  nand GNAME3380(G3380,G1275,G1290);
  nand GNAME3381(G3381,G1630,G22753);
  nand GNAME3382(G3382,G1274,G1290);
  nand GNAME3383(G3383,G1630,G22752);
  nand GNAME3384(G3384,G1273,G1290);
  nand GNAME3385(G3385,G1630,G22751);
  nand GNAME3386(G3386,G1272,G1290);
  nand GNAME3387(G3387,G1630,G22750);
  nand GNAME3388(G3388,G1271,G1290);
  nand GNAME3389(G3389,G1630,G22749);
  nand GNAME3390(G3390,G1270,G1290);
  nand GNAME3391(G3391,G1630,G22748);
  nand GNAME3392(G3392,G1269,G1290);
  nand GNAME3393(G3393,G1630,G22747);
  nand GNAME3394(G3394,G1268,G1290);
  nand GNAME3395(G3395,G1630,G22746);
  nand GNAME3396(G3396,G1267,G1290);
  nand GNAME3397(G3397,G1630,G22745);
  nand GNAME3398(G3398,G1266,G1290);
  nand GNAME3399(G3399,G1630,G22744);
  nand GNAME3400(G3400,G1265,G1290);
  nand GNAME3401(G3401,G1630,G22743);
  nand GNAME3402(G3402,G1264,G1290);
  nand GNAME3403(G3403,G1630,G22742);
  nand GNAME3404(G3404,G1263,G1290);
  nand GNAME3405(G3405,G1630,G22741);
  nand GNAME3406(G3406,G1262,G1290);
  nand GNAME3407(G3407,G1630,G22740);
  nand GNAME3408(G3408,G1261,G1290);
  nand GNAME3409(G3409,G1630,G22739);
  nand GNAME3410(G3410,G1260,G1290);
  nand GNAME3411(G3411,G1630,G22738);
  nand GNAME3412(G3412,G1259,G1290);
  nand GNAME3413(G3413,G1630,G22737);
  nand GNAME3414(G3414,G1258,G1290);
  nand GNAME3415(G3415,G1630,G22736);
  nand GNAME3416(G3416,G1257,G1290);
  nand GNAME3417(G3417,G22798,G1287,G1992,G1366);
  nand GNAME3418(G3418,G1066,G22791);
  nand GNAME3419(G3419,G2100,G22715);
  nand GNAME3420(G3420,G2103,G1301);
  nand GNAME3421(G3421,G2100,G22714);
  nand GNAME3422(G3422,G2106,G1301);
  nand GNAME3423(G3423,G2100,G22713);
  nand GNAME3424(G3424,G1301,G2114,G1235);
  nand GNAME3425(G3425,G2100,G22685);
  nand GNAME3426(G3426,G2315,G1301);
  nand GNAME3427(G3427,G2324,G22683);
  nand GNAME3428(G3428,G2329,G1625);
  nand GNAME3429(G3429,G2324,G22682);
  nand GNAME3430(G3430,G2332,G1625);
  nand GNAME3431(G3431,G2324,G22681);
  nand GNAME3432(G3432,G2340,G1625);
  nand GNAME3433(G3433,G2324,G22680);
  nand GNAME3434(G3434,G2346,G1625);
  nand GNAME3435(G3435,G2324,G22679);
  nand GNAME3436(G3436,G2352,G1625);
  nand GNAME3437(G3437,G2324,G22678);
  nand GNAME3438(G3438,G2358,G1625);
  nand GNAME3439(G3439,G2324,G22677);
  nand GNAME3440(G3440,G2364,G1625);
  nand GNAME3441(G3441,G2324,G22676);
  nand GNAME3442(G3442,G2370,G1625);
  nand GNAME3443(G3443,G2324,G22675);
  nand GNAME3444(G3444,G2376,G1625);
  nand GNAME3445(G3445,G2324,G22674);
  nand GNAME3446(G3446,G2382,G1625);
  nand GNAME3447(G3447,G2324,G22673);
  nand GNAME3448(G3448,G2388,G1625);
  nand GNAME3449(G3449,G2324,G22672);
  nand GNAME3450(G3450,G2394,G1625);
  nand GNAME3451(G3451,G2324,G22671);
  nand GNAME3452(G3452,G2400,G1625);
  nand GNAME3453(G3453,G2324,G22670);
  nand GNAME3454(G3454,G2406,G1625);
  nand GNAME3455(G3455,G2324,G22669);
  nand GNAME3456(G3456,G2412,G1625);
  nand GNAME3457(G3457,G2324,G22668);
  nand GNAME3458(G3458,G2418,G1625);
  nand GNAME3459(G3459,G2324,G22667);
  nand GNAME3460(G3460,G2424,G1625);
  nand GNAME3461(G3461,G2324,G22666);
  nand GNAME3462(G3462,G2430,G1625);
  nand GNAME3463(G3463,G2324,G22665);
  nand GNAME3464(G3464,G2436,G1625);
  nand GNAME3465(G3465,G2324,G22664);
  nand GNAME3466(G3466,G2442,G1625);
  nand GNAME3467(G3467,G2324,G22663);
  nand GNAME3468(G3468,G2448,G1625);
  nand GNAME3469(G3469,G2324,G22662);
  nand GNAME3470(G3470,G2454,G1625);
  nand GNAME3471(G3471,G2324,G22661);
  nand GNAME3472(G3472,G2460,G1625);
  nand GNAME3473(G3473,G2324,G22660);
  nand GNAME3474(G3474,G2466,G1625);
  nand GNAME3475(G3475,G2324,G22659);
  nand GNAME3476(G3476,G2472,G1625);
  nand GNAME3477(G3477,G2324,G22658);
  nand GNAME3478(G3478,G2478,G1625);
  nand GNAME3479(G3479,G2324,G22657);
  nand GNAME3480(G3480,G2484,G1625);
  nand GNAME3481(G3481,G2324,G22656);
  nand GNAME3482(G3482,G2490,G1625);
  nand GNAME3483(G3483,G2324,G22655);
  nand GNAME3484(G3484,G2496,G1625);
  nand GNAME3485(G3485,G2324,G22654);
  nand GNAME3486(G3486,G2502,G1625);
  nand GNAME3487(G3487,G2324,G22653);
  nand GNAME3488(G3488,G2506,G1625);
  nand GNAME3489(G3489,G2324,G22652);
  nand GNAME3490(G3490,G2511,G1625);
  nand GNAME3491(G3491,G2329,G1626);
  nand GNAME3492(G3492,G2512,G22651);
  nand GNAME3493(G3493,G2332,G1626);
  nand GNAME3494(G3494,G2512,G22650);
  nand GNAME3495(G3495,G2340,G1626);
  nand GNAME3496(G3496,G2512,G22649);
  nand GNAME3497(G3497,G2346,G1626);
  nand GNAME3498(G3498,G2512,G22648);
  nand GNAME3499(G3499,G2352,G1626);
  nand GNAME3500(G3500,G2512,G22647);
  nand GNAME3501(G3501,G2358,G1626);
  nand GNAME3502(G3502,G2512,G22646);
  nand GNAME3503(G3503,G2364,G1626);
  nand GNAME3504(G3504,G2512,G22645);
  nand GNAME3505(G3505,G2370,G1626);
  nand GNAME3506(G3506,G2512,G22644);
  nand GNAME3507(G3507,G2376,G1626);
  nand GNAME3508(G3508,G2512,G22643);
  nand GNAME3509(G3509,G2382,G1626);
  nand GNAME3510(G3510,G2512,G22642);
  nand GNAME3511(G3511,G2388,G1626);
  nand GNAME3512(G3512,G2512,G22641);
  nand GNAME3513(G3513,G2394,G1626);
  nand GNAME3514(G3514,G2512,G22640);
  nand GNAME3515(G3515,G2400,G1626);
  nand GNAME3516(G3516,G2512,G22639);
  nand GNAME3517(G3517,G2406,G1626);
  nand GNAME3518(G3518,G2512,G22638);
  nand GNAME3519(G3519,G2412,G1626);
  nand GNAME3520(G3520,G2512,G22637);
  nand GNAME3521(G3521,G2418,G1626);
  nand GNAME3522(G3522,G2512,G22636);
  nand GNAME3523(G3523,G2424,G1626);
  nand GNAME3524(G3524,G2512,G22635);
  nand GNAME3525(G3525,G2430,G1626);
  nand GNAME3526(G3526,G2512,G22634);
  nand GNAME3527(G3527,G2436,G1626);
  nand GNAME3528(G3528,G2512,G22633);
  nand GNAME3529(G3529,G2442,G1626);
  nand GNAME3530(G3530,G2512,G22632);
  nand GNAME3531(G3531,G2448,G1626);
  nand GNAME3532(G3532,G2512,G22631);
  nand GNAME3533(G3533,G2454,G1626);
  nand GNAME3534(G3534,G2512,G22630);
  nand GNAME3535(G3535,G2460,G1626);
  nand GNAME3536(G3536,G2512,G22629);
  nand GNAME3537(G3537,G2466,G1626);
  nand GNAME3538(G3538,G2512,G22628);
  nand GNAME3539(G3539,G2472,G1626);
  nand GNAME3540(G3540,G2512,G22627);
  nand GNAME3541(G3541,G2478,G1626);
  nand GNAME3542(G3542,G2512,G22626);
  nand GNAME3543(G3543,G2484,G1626);
  nand GNAME3544(G3544,G2512,G22625);
  nand GNAME3545(G3545,G2490,G1626);
  nand GNAME3546(G3546,G2512,G22624);
  nand GNAME3547(G3547,G2496,G1626);
  nand GNAME3548(G3548,G2512,G22623);
  nand GNAME3549(G3549,G2502,G1626);
  nand GNAME3550(G3550,G2512,G22622);
  nand GNAME3551(G3551,G2506,G1626);
  nand GNAME3552(G3552,G2512,G22621);
  nand GNAME3553(G3553,G2511,G1626);
  nand GNAME3554(G3554,G2512,G22620);
  nand GNAME3555(G3555,G1772,G1627);
  nand GNAME3556(G3556,G2513,G22589);
  nand GNAME3557(G3557,G1771,G1627);
  nand GNAME3558(G3558,G2513,G22588);
  nand GNAME3559(G3559,G1366,G1364);
  nand GNAME3560(G3560,G7011,G3112);
  or GNAME3561(G3561,G1225,G3115);
  or GNAME3562(G3562,G3197,G1367);
  or GNAME3563(G3563,G3209,G1401);
  or GNAME3564(G3564,G3206,G1402);
  nand GNAME3565(G3565,G22661,G1365);
  nand GNAME3566(G3566,G22693,G3109);
  nand GNAME3567(G3567,G22660,G1365);
  nand GNAME3568(G3568,G22692,G3109);
  nand GNAME3569(G3569,G22659,G1365);
  nand GNAME3570(G3570,G22691,G3109);
  nand GNAME3571(G3571,G22658,G1365);
  nand GNAME3572(G3572,G22690,G3109);
  nand GNAME3573(G3573,G22657,G1365);
  nand GNAME3574(G3574,G22689,G3109);
  nand GNAME3575(G3575,G22656,G1365);
  nand GNAME3576(G3576,G22688,G3109);
  nand GNAME3577(G3577,G22655,G1365);
  nand GNAME3578(G3578,G22687,G3109);
  nand GNAME3579(G3579,G22654,G1365);
  nand GNAME3580(G3580,G22686,G3109);
  nand GNAME3581(G3581,G22671,G1365);
  nand GNAME3582(G3582,G22703,G3109);
  nand GNAME3583(G3583,G22670,G1365);
  nand GNAME3584(G3584,G22702,G3109);
  nand GNAME3585(G3585,G22669,G1365);
  nand GNAME3586(G3586,G22701,G3109);
  nand GNAME3587(G3587,G22668,G1365);
  nand GNAME3588(G3588,G22700,G3109);
  nand GNAME3589(G3589,G22667,G1365);
  nand GNAME3590(G3590,G22699,G3109);
  nand GNAME3591(G3591,G22666,G1365);
  nand GNAME3592(G3592,G22698,G3109);
  nand GNAME3593(G3593,G22665,G1365);
  nand GNAME3594(G3594,G22697,G3109);
  nand GNAME3595(G3595,G22664,G1365);
  nand GNAME3596(G3596,G22696,G3109);
  nand GNAME3597(G3597,G22663,G1365);
  nand GNAME3598(G3598,G22695,G3109);
  nand GNAME3599(G3599,G22662,G1365);
  nand GNAME3600(G3600,G22694,G3109);
  nand GNAME3601(G3601,G22653,G1365);
  nand GNAME3602(G3602,G22685,G3109);
  nand GNAME3603(G3603,G22652,G1365);
  nand GNAME3604(G3604,G22684,G3109);
  not GNAME3605(G3605,G1216);
  not GNAME3606(G3606,G7957);
  not GNAME3607(G3607,G1286);
  or GNAME3608(G3608,G4096,G6345);
  nand GNAME3609(G3609,G3610,G3612,G3611);
  nand GNAME3610(G3610,G6347,G4093);
  or GNAME3611(G3611,G4246,G6346);
  nand GNAME3612(G3612,G3613,G3615,G3614);
  nand GNAME3613(G3613,G6348,G4248);
  or GNAME3614(G3614,G4093,G6347);
  nand GNAME3615(G3615,G3616,G3618,G3617);
  nand GNAME3616(G3616,G6349,G4095);
  or GNAME3617(G3617,G4248,G6348);
  nand GNAME3618(G3618,G3619,G3621,G3620);
  nand GNAME3619(G3619,G6350,G4250);
  or GNAME3620(G3620,G4095,G6349);
  nand GNAME3621(G3621,G3622,G3624,G3623);
  nand GNAME3622(G3622,G6351,G4182);
  or GNAME3623(G3623,G4250,G6350);
  nand GNAME3624(G3624,G3625,G3627,G3626);
  nand GNAME3625(G3625,G6352,G4253);
  or GNAME3626(G3626,G4182,G6351);
  nand GNAME3627(G3627,G3628,G3630,G3629);
  nand GNAME3628(G3628,G6353,G4188);
  or GNAME3629(G3629,G4253,G6352);
  nand GNAME3630(G3630,G3631,G3633,G3632);
  nand GNAME3631(G3631,G6354,G4255);
  or GNAME3632(G3632,G4188,G6353);
  nand GNAME3633(G3633,G3634,G3636,G3635);
  nand GNAME3634(G3634,G6355,G4197);
  or GNAME3635(G3635,G4255,G6354);
  nand GNAME3636(G3636,G3637,G3639,G3638);
  nand GNAME3637(G3637,G6356,G4257);
  or GNAME3638(G3638,G4197,G6355);
  nand GNAME3639(G3639,G3640,G3642,G3641);
  nand GNAME3640(G3640,G6357,G4192);
  or GNAME3641(G3641,G4257,G6356);
  nand GNAME3642(G3642,G3643,G3645,G3644);
  nand GNAME3643(G3643,G6358,G4259);
  or GNAME3644(G3644,G4192,G6357);
  nand GNAME3645(G3645,G3646,G3648,G3647);
  nand GNAME3646(G3646,G6359,G4193);
  or GNAME3647(G3647,G4259,G6358);
  nand GNAME3648(G3648,G3649,G3651,G3650);
  nand GNAME3649(G3649,G6360,G4261);
  or GNAME3650(G3650,G4193,G6359);
  nand GNAME3651(G3651,G3652,G3654,G3653);
  nand GNAME3652(G3652,G6361,G4190);
  or GNAME3653(G3653,G4261,G6360);
  nand GNAME3654(G3654,G3655,G3657,G3656);
  nand GNAME3655(G3655,G6362,G4233);
  or GNAME3656(G3656,G4190,G6361);
  nand GNAME3657(G3657,G3658,G3660,G3659);
  nand GNAME3658(G3658,G6363,G4178);
  or GNAME3659(G3659,G4233,G6362);
  nand GNAME3660(G3660,G3661,G3663,G3662);
  nand GNAME3661(G3661,G6364,G4235);
  or GNAME3662(G3662,G4178,G6363);
  nand GNAME3663(G3663,G3664,G3666,G3665);
  nand GNAME3664(G3664,G6365,G4187);
  or GNAME3665(G3665,G4235,G6364);
  nand GNAME3666(G3666,G3667,G3669,G3668);
  nand GNAME3667(G3667,G6366,G4237);
  or GNAME3668(G3668,G4187,G6365);
  nand GNAME3669(G3669,G3670,G3672,G3671);
  nand GNAME3670(G3670,G6367,G4181);
  or GNAME3671(G3671,G4237,G6366);
  nand GNAME3672(G3672,G3673,G3675,G3674);
  nand GNAME3673(G3673,G6368,G4251);
  or GNAME3674(G3674,G4181,G6367);
  nand GNAME3675(G3675,G3676,G3678,G3677);
  nand GNAME3676(G3676,G6369,G4184);
  or GNAME3677(G3677,G4251,G6368);
  nand GNAME3678(G3678,G4191,G6338,G3679);
  or GNAME3679(G3679,G4184,G6369);
  nand GNAME3680(G3680,G5809,G5807,G5808);
  nand GNAME3681(G3681,G4371,G4766,G4767,G4768);
  nand GNAME3682(G3682,G5812,G5810,G5811);
  nand GNAME3683(G3683,G4371,G4769,G4770,G4771);
  nand GNAME3684(G3684,G5816,G5817,G5818,G4146);
  nand GNAME3685(G3685,G4371,G4530,G4531,G4532);
  nand GNAME3686(G3686,G5819,G5820,G5821,G4146);
  nand GNAME3687(G3687,G4430,G4431,G4432,G4433);
  nand GNAME3688(G3688,G5822,G5823,G5824,G4146);
  nand GNAME3689(G3689,G4533,G4534,G4535,G4536);
  nand GNAME3690(G3690,G5825,G5826,G5827,G4146);
  nand GNAME3691(G3691,G4434,G4435,G4436,G4437);
  nand GNAME3692(G3692,G5828,G5829,G5830,G4146);
  nand GNAME3693(G3693,G4623,G4624,G4625,G4626);
  nand GNAME3694(G3694,G5831,G5832,G5833,G4146);
  nand GNAME3695(G3695,G4463,G4464,G4465,G4466);
  nand GNAME3696(G3696,G5834,G5835,G5836,G4146);
  nand GNAME3697(G3697,G4627,G4628,G4629,G4630);
  nand GNAME3698(G3698,G5837,G5838,G5839,G4146);
  nand GNAME3699(G3699,G4467,G4468,G4469,G4470);
  nand GNAME3700(G3700,G5840,G5841,G5842,G4146);
  nand GNAME3701(G3701,G4680,G4681,G4682,G4683);
  nand GNAME3702(G3702,G5843,G5844,G5845,G4146);
  nand GNAME3703(G3703,G4513,G4514,G4515,G4516);
  nand GNAME3704(G3704,G5849,G5850,G5851,G4146);
  nand GNAME3705(G3705,G4684,G4685,G4686,G4687);
  nand GNAME3706(G3706,G5852,G5853,G5854,G4146);
  nand GNAME3707(G3707,G4517,G4518,G4519,G4520);
  nand GNAME3708(G3708,G5855,G5856,G5857,G4146);
  nand GNAME3709(G3709,G4589,G4590,G4591,G4592);
  nand GNAME3710(G3710,G5858,G5859,G5860,G4146);
  nand GNAME3711(G3711,G4610,G4611,G4612,G4613);
  nand GNAME3712(G3712,G5861,G5862,G5863,G4146);
  nand GNAME3713(G3713,G4445,G4446,G4447,G4448);
  nand GNAME3714(G3714,G5864,G5865,G5866,G4146);
  nand GNAME3715(G3715,G4695,G4696,G4697,G4698);
  nand GNAME3716(G3716,G5867,G5868,G5869,G4146);
  nand GNAME3717(G3717,G4450,G4451,G4452,G4453);
  nand GNAME3718(G3718,G5870,G5871,G5872,G4146);
  nand GNAME3719(G3719,G4700,G4701,G4702,G4703);
  nand GNAME3720(G3720,G5873,G5874,G5875,G4146);
  nand GNAME3721(G3721,G4477,G4478,G4479,G4480);
  nand GNAME3722(G3722,G5876,G5877,G5878,G4146);
  nand GNAME3723(G3723,G4655,G4656,G4657,G4658);
  nand GNAME3724(G3724,G5789,G5790,G5791,G4146);
  nand GNAME3725(G3725,G4482,G4483,G4484,G4485);
  nand GNAME3726(G3726,G5792,G5793,G5794,G4146);
  nand GNAME3727(G3727,G4380,G4381,G4382,G4383);
  nand GNAME3728(G3728,G5795,G5796,G5797,G4146);
  nand GNAME3729(G3729,G4543,G4544,G4545,G4546);
  nand GNAME3730(G3730,G5798,G5799,G5800,G4146);
  nand GNAME3731(G3731,G4385,G4386,G4387,G4388);
  nand GNAME3732(G3732,G5801,G5802,G5803,G4146);
  nand GNAME3733(G3733,G4637,G4638,G4639,G4640);
  nand GNAME3734(G3734,G5804,G5805,G5806,G4146);
  nand GNAME3735(G3735,G4495,G4496,G4497,G4498);
  nand GNAME3736(G3736,G5813,G5814,G5815,G4146);
  nand GNAME3737(G3737,G4642,G4643,G4644,G4645);
  nand GNAME3738(G3738,G5846,G5847,G5848,G4146);
  nand GNAME3739(G3739,G4500,G4501,G4502,G4503);
  nand GNAME3740(G3740,G5879,G5880,G5881,G4146);
  nand GNAME3741(G3741,G4668,G4669,G4670,G4671);
  nand GNAME3742(G3742,G5882,G5883,G5884,G4146);
  nand GNAME3743(G3743,G4556,G4557,G4558,G4559);
  nand GNAME3744(G3744,G5712,G5713);
  nand GNAME3745(G3745,G5714,G5715);
  nand GNAME3746(G3746,G5721,G5719,G5720);
  nand GNAME3747(G3747,G5724,G5722,G5723);
  nand GNAME3748(G3748,G5727,G5725,G5726);
  nand GNAME3749(G3749,G5730,G5728,G5729);
  nand GNAME3750(G3750,G5733,G5731,G5732);
  nand GNAME3751(G3751,G5736,G5734,G5735);
  nand GNAME3752(G3752,G5739,G5737,G5738);
  nand GNAME3753(G3753,G5742,G5740,G5741);
  nand GNAME3754(G3754,G5745,G5743,G5744);
  nand GNAME3755(G3755,G5748,G5746,G5747);
  nand GNAME3756(G3756,G5754,G5752,G5753);
  nand GNAME3757(G3757,G5757,G5755,G5756);
  nand GNAME3758(G3758,G5760,G5758,G5759);
  nand GNAME3759(G3759,G5763,G5761,G5762);
  nand GNAME3760(G3760,G5766,G5764,G5765);
  nand GNAME3761(G3761,G5769,G5767,G5768);
  nand GNAME3762(G3762,G5772,G5770,G5771);
  nand GNAME3763(G3763,G5775,G5773,G5774);
  nand GNAME3764(G3764,G5778,G5776,G5777);
  nand GNAME3765(G3765,G5781,G5779,G5780);
  nand GNAME3766(G3766,G5696,G5694,G5695);
  nand GNAME3767(G3767,G5699,G5697,G5698);
  nand GNAME3768(G3768,G5702,G5700,G5701);
  nand GNAME3769(G3769,G5705,G5703,G5704);
  nand GNAME3770(G3770,G5708,G5706,G5707);
  nand GNAME3771(G3771,G5711,G5709,G5710);
  nand GNAME3772(G3772,G5718,G5716,G5717);
  nand GNAME3773(G3773,G5751,G5749,G5750);
  nand GNAME3774(G3774,G5784,G5782,G5783);
  nand GNAME3775(G3775,G5785,G5786);
  nand GNAME3776(G3776,G4375,G4053,G5689,G5891);
  or GNAME3777(G3777,G3778,G4147);
  nand GNAME3778(G3778,G5628,G5629,G5627,G5625,G5626);
  nand GNAME3779(G3779,G5634,G5625,G5633);
  nand GNAME3780(G3780,G5636,G5625,G5635);
  nand GNAME3781(G3781,G5638,G5625,G5637);
  nand GNAME3782(G3782,G5640,G5625,G5639);
  nand GNAME3783(G3783,G5642,G5625,G5641);
  nand GNAME3784(G3784,G5644,G5625,G5643);
  nand GNAME3785(G3785,G5646,G5625,G5645);
  nand GNAME3786(G3786,G5648,G5625,G5647);
  nand GNAME3787(G3787,G5650,G5625,G5649);
  nand GNAME3788(G3788,G5655,G5625,G5654);
  nand GNAME3789(G3789,G5658,G5656,G5657);
  nand GNAME3790(G3790,G5661,G5659,G5660);
  nand GNAME3791(G3791,G5664,G5662,G5663);
  nand GNAME3792(G3792,G5667,G5665,G5666);
  nand GNAME3793(G3793,G5670,G5668,G5669);
  nand GNAME3794(G3794,G5673,G5671,G5672);
  nand GNAME3795(G3795,G5676,G5674,G5675);
  nand GNAME3796(G3796,G5679,G5677,G5678);
  nand GNAME3797(G3797,G5682,G5680,G5681);
  nand GNAME3798(G3798,G5609,G5607,G5608);
  nand GNAME3799(G3799,G5612,G5610,G5611);
  nand GNAME3800(G3800,G5615,G5613,G5614);
  nand GNAME3801(G3801,G5618,G5616,G5617);
  nand GNAME3802(G3802,G5621,G5619,G5620);
  nand GNAME3803(G3803,G5624,G5622,G5623);
  nand GNAME3804(G3804,G5632,G5630,G5631);
  nand GNAME3805(G3805,G5653,G5651,G5652);
  nand GNAME3806(G3806,G5685,G5683,G5684);
  nand GNAME3807(G3807,G5688,G5686,G5687);
  nand GNAME3808(G3808,G5531,G4142);
  nand GNAME3809(G3809,G5532,G4142);
  nand GNAME3810(G3810,G5537,G4142);
  nand GNAME3811(G3811,G4141,G5538,G5539);
  nand GNAME3812(G3812,G4141,G5540,G5541);
  nand GNAME3813(G3813,G4141,G5542,G5543);
  nand GNAME3814(G3814,G4141,G5544,G5545);
  nand GNAME3815(G3815,G4141,G5546,G5547);
  nand GNAME3816(G3816,G4141,G5548,G5549);
  nand GNAME3817(G3817,G4141,G5550,G5551);
  nand GNAME3818(G3818,G4141,G5552,G5553);
  nand GNAME3819(G3819,G4141,G5554,G5555);
  nand GNAME3820(G3820,G4141,G5560,G5561);
  nand GNAME3821(G3821,G5562,G5563,G5564,G5565);
  nand GNAME3822(G3822,G5566,G5567,G5568,G5569);
  nand GNAME3823(G3823,G5570,G5571,G5572,G5573);
  nand GNAME3824(G3824,G5574,G5575,G5576,G5577);
  nand GNAME3825(G3825,G5578,G5579,G5580,G5581);
  nand GNAME3826(G3826,G5582,G5583,G5584,G5585);
  nand GNAME3827(G3827,G5586,G5587,G5588,G5589);
  nand GNAME3828(G3828,G5590,G5591,G5592,G5593);
  nand GNAME3829(G3829,G5594,G5595,G5596,G5597);
  nand GNAME3830(G3830,G5501,G5502,G5503,G5504);
  nand GNAME3831(G3831,G5505,G5506,G5507,G5508);
  nand GNAME3832(G3832,G5509,G5510,G5511,G5512);
  nand GNAME3833(G3833,G5513,G5514,G5515,G5516);
  nand GNAME3834(G3834,G5517,G5518,G5519,G5520);
  nand GNAME3835(G3835,G5521,G5522,G5523,G5524);
  nand GNAME3836(G3836,G5533,G5534,G5535,G5536);
  nand GNAME3837(G3837,G5556,G5557,G5558,G5559);
  nand GNAME3838(G3838,G5598,G5599,G5600,G5601);
  nand GNAME3839(G3839,G5602,G5603,G5604,G5605);
  nand GNAME3840(G3840,G4379,G4058);
  not GNAME3841(G3841,G23043);
  nand GNAME3842(G3842,G5488,G5486,G5487);
  nand GNAME3843(G3843,G5485,G5483,G5484);
  nand GNAME3844(G3844,G5482,G5480,G5481);
  nand GNAME3845(G3845,G5479,G5477,G5478);
  nand GNAME3846(G3846,G5476,G5474,G5475);
  nand GNAME3847(G3847,G5473,G5471,G5472);
  nand GNAME3848(G3848,G5470,G5468,G5469);
  nand GNAME3849(G3849,G5467,G5465,G5466);
  nand GNAME3850(G3850,G5464,G5462,G5463);
  nand GNAME3851(G3851,G5461,G5459,G5460);
  nand GNAME3852(G3852,G5458,G5456,G5457);
  nand GNAME3853(G3853,G5455,G5453,G5454);
  nand GNAME3854(G3854,G5452,G5450,G5451);
  nand GNAME3855(G3855,G5449,G5447,G5448);
  nand GNAME3856(G3856,G5446,G5444,G5445);
  nand GNAME3857(G3857,G5443,G5441,G5442);
  nand GNAME3858(G3858,G5440,G5438,G5439);
  nand GNAME3859(G3859,G5437,G5435,G5436);
  nand GNAME3860(G3860,G5434,G5432,G5433);
  nand GNAME3861(G3861,G5431,G5429,G5430);
  nand GNAME3862(G3862,G5428,G5426,G5427);
  nand GNAME3863(G3863,G5425,G5423,G5424);
  nand GNAME3864(G3864,G5422,G5420,G5421);
  nand GNAME3865(G3865,G5419,G5417,G5418);
  nand GNAME3866(G3866,G5416,G5414,G5415);
  nand GNAME3867(G3867,G5413,G5411,G5412);
  nand GNAME3868(G3868,G5410,G5408,G5409);
  nand GNAME3869(G3869,G5407,G5405,G5406);
  nand GNAME3870(G3870,G5404,G5402,G5403);
  nand GNAME3871(G3871,G5401,G5399,G5400);
  nand GNAME3872(G3872,G5398,G5396,G5397);
  nand GNAME3873(G3873,G5395,G5393,G5394);
  and GNAME3874(G3874,G5392,G22835);
  and GNAME3875(G3875,G5392,G22836);
  and GNAME3876(G3876,G5392,G22837);
  and GNAME3877(G3877,G5392,G22838);
  and GNAME3878(G3878,G5392,G22839);
  and GNAME3879(G3879,G5392,G22840);
  and GNAME3880(G3880,G5392,G22841);
  and GNAME3881(G3881,G5392,G22842);
  and GNAME3882(G3882,G5392,G22843);
  and GNAME3883(G3883,G5392,G22844);
  and GNAME3884(G3884,G5392,G22845);
  and GNAME3885(G3885,G5392,G22846);
  and GNAME3886(G3886,G5392,G22847);
  and GNAME3887(G3887,G5392,G22848);
  and GNAME3888(G3888,G5392,G22849);
  and GNAME3889(G3889,G5392,G22850);
  and GNAME3890(G3890,G5392,G22851);
  and GNAME3891(G3891,G5392,G22852);
  and GNAME3892(G3892,G5392,G22853);
  and GNAME3893(G3893,G5392,G22854);
  and GNAME3894(G3894,G5392,G22855);
  and GNAME3895(G3895,G5392,G22856);
  and GNAME3896(G3896,G5392,G22857);
  and GNAME3897(G3897,G5392,G22858);
  and GNAME3898(G3898,G5392,G22859);
  and GNAME3899(G3899,G5392,G22860);
  and GNAME3900(G3900,G5392,G22861);
  and GNAME3901(G3901,G5392,G22862);
  and GNAME3902(G3902,G5392,G22863);
  and GNAME3903(G3903,G5392,G22864);
  nand GNAME3904(G3904,G5388,G5389,G5390,G5391);
  nand GNAME3905(G3905,G5386,G5387,G5385,G5383,G5384);
  nand GNAME3906(G3906,G5381,G5382,G5380,G5378,G5379);
  nand GNAME3907(G3907,G5376,G5377,G5375,G5373,G5374);
  nand GNAME3908(G3908,G5371,G5372,G5370,G5368,G5369);
  nand GNAME3909(G3909,G5366,G5367,G5365,G5363,G5364);
  nand GNAME3910(G3910,G5361,G5362,G5360,G5358,G5359);
  nand GNAME3911(G3911,G5356,G5357,G5355,G5353,G5354);
  nand GNAME3912(G3912,G5351,G5352,G5350,G5348,G5349);
  nand GNAME3913(G3913,G5346,G5347,G5345,G5343,G5344);
  nand GNAME3914(G3914,G5341,G5342,G5340,G5338,G5339);
  nand GNAME3915(G3915,G5336,G5337,G5335,G5333,G5334);
  nand GNAME3916(G3916,G5331,G5332,G5330,G5328,G5329);
  nand GNAME3917(G3917,G5326,G5327,G5325,G5323,G5324);
  nand GNAME3918(G3918,G5321,G5322,G5320,G5318,G5319);
  nand GNAME3919(G3919,G5316,G5317,G5315,G5313,G5314);
  nand GNAME3920(G3920,G5311,G5312,G5310,G5308,G5309);
  nand GNAME3921(G3921,G5306,G5307,G5305,G5303,G5304);
  nand GNAME3922(G3922,G5301,G5302,G5300,G5298,G5299);
  nand GNAME3923(G3923,G5296,G5297,G5295,G5293,G5294);
  nand GNAME3924(G3924,G5291,G5292,G5290,G5288,G5289);
  nand GNAME3925(G3925,G5286,G5287,G5285,G5283,G5284);
  nand GNAME3926(G3926,G5281,G5282,G5280,G5278,G5279);
  nand GNAME3927(G3927,G5276,G5277,G5275,G5273,G5274);
  nand GNAME3928(G3928,G5271,G5272,G5270,G5268,G5269);
  nand GNAME3929(G3929,G5266,G5267,G5265,G5263,G5264);
  nand GNAME3930(G3930,G5261,G5262,G5260,G5258,G5259);
  nand GNAME3931(G3931,G5256,G5257,G5255,G5253,G5254);
  nand GNAME3932(G3932,G5251,G5252,G5250,G5248,G5249);
  nand GNAME3933(G3933,G5245,G5246,G5247,G6226,G6227);
  nand GNAME3934(G3934,G5244,G4372,G5243);
  nand GNAME3935(G3935,G5242,G4372,G5241);
  nand GNAME3936(G3936,G5231,G5232,G5233,G5234);
  nand GNAME3937(G3937,G5229,G5230,G5228,G5226,G5227);
  nand GNAME3938(G3938,G5224,G5225,G5223,G5221,G5222);
  nand GNAME3939(G3939,G5219,G5220,G5218,G5216,G5217);
  nand GNAME3940(G3940,G5214,G5215,G5213,G5211,G5212);
  nand GNAME3941(G3941,G5209,G5210,G5208,G5206,G5207);
  nand GNAME3942(G3942,G5204,G5205,G5203,G5201,G5202);
  nand GNAME3943(G3943,G5199,G5200,G5198,G5196,G5197);
  nand GNAME3944(G3944,G5194,G5195,G5193,G5191,G5192);
  nand GNAME3945(G3945,G5189,G5190,G5188,G5186,G5187);
  nand GNAME3946(G3946,G5184,G5185,G5183,G5181,G5182);
  nand GNAME3947(G3947,G5179,G5180,G5178,G5176,G5177);
  nand GNAME3948(G3948,G5174,G5175,G5173,G5171,G5172);
  nand GNAME3949(G3949,G5169,G5170,G5168,G5166,G5167);
  nand GNAME3950(G3950,G5164,G5165,G5163,G5161,G5162);
  nand GNAME3951(G3951,G5159,G5160,G5158,G5156,G5157);
  nand GNAME3952(G3952,G5154,G5155,G5153,G5151,G5152);
  nand GNAME3953(G3953,G5149,G5150,G5148,G5146,G5147);
  nand GNAME3954(G3954,G5144,G5145,G5143,G5141,G5142);
  nand GNAME3955(G3955,G5139,G5140,G5138,G5136,G5137);
  nand GNAME3956(G3956,G5134,G5135,G5133,G5131,G5132);
  nand GNAME3957(G3957,G5129,G5130,G5128,G5126,G5127);
  nand GNAME3958(G3958,G5124,G5125,G5123,G5121,G5122);
  nand GNAME3959(G3959,G5119,G5120,G5118,G5116,G5117);
  nand GNAME3960(G3960,G5114,G5115,G5113,G5111,G5112);
  nand GNAME3961(G3961,G5109,G5110,G5108,G5106,G5107);
  nand GNAME3962(G3962,G5104,G5105,G5103,G5101,G5102);
  nand GNAME3963(G3963,G5099,G5100,G5098,G5096,G5097);
  nand GNAME3964(G3964,G5094,G5095,G5093,G5091,G5092);
  nand GNAME3965(G3965,G5088,G5089,G5090,G6221,G6222);
  nand GNAME3966(G3966,G5085,G4373,G5084);
  nand GNAME3967(G3967,G5083,G4373,G5082);
  nand GNAME3968(G3968,G5076,G5077,G5075,G5073,G5074);
  nand GNAME3969(G3969,G5072,G4362,G5071,G5069,G5070);
  nand GNAME3970(G3970,G4355,G5064,G5062,G5063);
  nand GNAME3971(G3971,G4354,G5058,G5056,G5057);
  nand GNAME3972(G3972,G4353,G5052,G5050,G5051);
  nand GNAME3973(G3973,G4352,G5046,G5044,G5045);
  nand GNAME3974(G3974,G4351,G5040,G5038,G5039);
  nand GNAME3975(G3975,G4350,G5034,G5032,G5033);
  nand GNAME3976(G3976,G4349,G5028,G5026,G5027);
  nand GNAME3977(G3977,G4348,G5022,G5020,G5021);
  nand GNAME3978(G3978,G4347,G5016,G5014,G5015);
  nand GNAME3979(G3979,G4346,G5010,G5008,G5009);
  nand GNAME3980(G3980,G4345,G5004,G5002,G5003);
  nand GNAME3981(G3981,G4344,G4998,G4996,G4997);
  nand GNAME3982(G3982,G4343,G4992,G4990,G4991);
  nand GNAME3983(G3983,G4342,G4986,G4984,G4985);
  nand GNAME3984(G3984,G4341,G4980,G4978,G4979);
  nand GNAME3985(G3985,G4340,G4974,G4972,G4973);
  nand GNAME3986(G3986,G4339,G4968,G4966,G4967);
  nand GNAME3987(G3987,G4338,G4962,G4960,G4961);
  nand GNAME3988(G3988,G4337,G4956,G4954,G4955);
  nand GNAME3989(G3989,G4336,G4950,G4948,G4949);
  nand GNAME3990(G3990,G4335,G4944,G4942,G4943);
  nand GNAME3991(G3991,G4334,G4938,G4936,G4937);
  nand GNAME3992(G3992,G4333,G4932,G4930,G4931);
  nand GNAME3993(G3993,G4332,G4926,G4924,G4925);
  nand GNAME3994(G3994,G4331,G4920,G4918,G4919);
  nand GNAME3995(G3995,G4330,G4914,G4912,G4913);
  nand GNAME3996(G3996,G4329,G4908,G4906,G4907);
  nand GNAME3997(G3997,G4902,G4361,G4901,G4899,G4900);
  nand GNAME3998(G3998,G4116,G4895,G4896);
  nand GNAME3999(G3999,G4116,G4893,G4894);
  nand GNAME4000(G4000,G4880,G4881,G4879,G4877,G4878);
  nand GNAME4001(G4001,G4875,G4876,G4874,G4872,G4873);
  nand GNAME4002(G4002,G4870,G4871,G4869,G4867,G4868);
  nand GNAME4003(G4003,G4865,G4866,G4864,G4862,G4863);
  nand GNAME4004(G4004,G4860,G4861,G4859,G4857,G4858);
  nand GNAME4005(G4005,G4855,G4856,G4854,G4852,G4853);
  nand GNAME4006(G4006,G4850,G4851,G4849,G4847,G4848);
  nand GNAME4007(G4007,G4845,G4846,G4844,G4842,G4843);
  nand GNAME4008(G4008,G4840,G4841,G4839,G4837,G4838);
  nand GNAME4009(G4009,G4835,G4836,G4834,G4832,G4833);
  nand GNAME4010(G4010,G4830,G4831,G4829,G4827,G4828);
  nand GNAME4011(G4011,G4825,G4826,G4824,G4822,G4823);
  nand GNAME4012(G4012,G4820,G4821,G4819,G4817,G4818);
  nand GNAME4013(G4013,G4815,G4816,G4814,G4812,G4813);
  nand GNAME4014(G4014,G4810,G4811,G4809,G4807,G4808);
  nand GNAME4015(G4015,G4805,G4806,G4804,G4802,G4803);
  nand GNAME4016(G4016,G4800,G4801,G4799,G4797,G4798);
  nand GNAME4017(G4017,G4795,G4796,G4794,G4792,G4793);
  nand GNAME4018(G4018,G4790,G4791,G4789,G4787,G4788);
  nand GNAME4019(G4019,G4785,G4786,G4784,G4782,G4783);
  nand GNAME4020(G4020,G6038,G6039,G4776,G4777);
  nand GNAME4021(G4021,G4320,G4759,G4760,G4761,G4762);
  nand GNAME4022(G4022,G4319,G4753,G4755,G4752);
  nand GNAME4023(G4023,G4318,G4745,G4746,G4747,G4748);
  nand GNAME4024(G4024,G4317,G4737,G4738,G4739,G4740);
  nand GNAME4025(G4025,G4316,G4729,G4730,G4731,G4732);
  nand GNAME4026(G4026,G4315,G4721,G4722,G4723,G4724);
  nand GNAME4027(G4027,G4314,G4715,G4713,G4714);
  nand GNAME4028(G4028,G4313,G4707,G4708,G4709,G4710);
  nand GNAME4029(G4029,G4312,G4691,G4689,G4690);
  nand GNAME4030(G4030,G4311,G4677,G4675,G4676);
  nand GNAME4031(G4031,G4310,G4662,G4663,G4664,G4665);
  nand GNAME4032(G4032,G4309,G4649,G4650,G4651,G4652);
  nand GNAME4033(G4033,G4308,G4633,G4631,G4632);
  nand GNAME4034(G4034,G4307,G4617,G4618,G4619,G4620);
  nand GNAME4035(G4035,G4306,G4604,G4605,G4606,G4607);
  nand GNAME4036(G4036,G4305,G4596,G4597,G4598,G4599);
  nand GNAME4037(G4037,G4304,G4585,G4583,G4584);
  nand GNAME4038(G4038,G4303,G4577,G4578,G4579,G4580);
  nand GNAME4039(G4039,G4302,G4571,G4569,G4570);
  nand GNAME4040(G4040,G4301,G4563,G4564,G4565,G4566);
  nand GNAME4041(G4041,G4300,G4550,G4551,G4552,G4553);
  nand GNAME4042(G4042,G4299,G4539,G4537,G4538);
  nand GNAME4043(G4043,G4298,G4524,G4525,G4526,G4527);
  nand GNAME4044(G4044,G4297,G4507,G4508,G4509,G4510);
  nand GNAME4045(G4045,G4296,G4489,G4490,G4491,G4492);
  nand GNAME4046(G4046,G4295,G4473,G4471,G4472);
  nand GNAME4047(G4047,G4294,G4457,G4458,G4459,G4460);
  nand GNAME4048(G4048,G4293,G4441,G4443,G4440);
  nand GNAME4049(G4049,G4292,G4424,G4425,G4426,G4427);
  nand GNAME4050(G4050,G5891,G4061);
  nand GNAME4051(G4051,G4176,G5938);
  not GNAME4052(G4052,G22832);
  nand GNAME4053(G4053,G4150,G4148,G4149);
  or GNAME4054(G4054,G4147,G4053);
  not GNAME4055(G4055,G8894);
  not GNAME4056(G4056,G22828);
  or GNAME4057(G4057,G4065,G4066);
  and GNAME4058(G4058,G23043,G4378);
  and GNAME4059(G4059,G5959,G5962);
  and GNAME4060(G4060,G4170,G4171);
  and GNAME4061(G4061,G4059,G4060);
  and GNAME4062(G4062,G5891,G23043,G4053);
  nand GNAME4063(G4063,G4148,G5967,G5968);
  and GNAME4064(G4064,G4395,G4396);
  and GNAME4065(G4065,G4052,G22829);
  and GNAME4066(G4066,G22832,G8866);
  nand GNAME4067(G4067,G4064,G5971,G5974);
  nor GNAME4068(G4068,G4411,G4366);
  not GNAME4069(G4069,G8861);
  not GNAME4070(G4070,G22830);
  not GNAME4071(G4071,G8893);
  and GNAME4072(G4072,G4068,G4423,G4400);
  and GNAME4073(G4073,G4420,G4421);
  and GNAME4074(G4074,G4068,G4422,G4400);
  and GNAME4075(G4075,G4174,G4173);
  and GNAME4076(G4076,G5941,G5938);
  nor GNAME4077(G4077,G5962,G5959);
  and GNAME4078(G4078,G5938,G4077);
  and GNAME4079(G4079,G5959,G5941);
  nand GNAME4080(G4080,G5941,G4170,G4175);
  nand GNAME4081(G4081,G4175,G5962);
  or GNAME4082(G4082,G5941,G4081);
  and GNAME4083(G4083,G4401,G4402);
  nand GNAME4084(G4084,G4403,G4404,G4405,G4083);
  nand GNAME4085(G4085,G4391,G4392);
  or GNAME4086(G4086,G5962,G4080);
  and GNAME4087(G4087,G4064,G4075);
  and GNAME4088(G4088,G4408,G4062);
  and GNAME4089(G4089,G4087,G4085,G4062);
  and GNAME4090(G4090,G4076,G4175,G5962);
  and GNAME4091(G4091,G4062,G4090);
  and GNAME4092(G4092,G4370,G559);
  and GNAME4093(G4093,G4370,G563);
  and GNAME4094(G4094,G4370,G558);
  and GNAME4095(G4095,G4370,G565);
  and GNAME4096(G4096,G4370,G561);
  and GNAME4097(G4097,G4370,G562);
  and GNAME4098(G4098,G4370,G566);
  and GNAME4099(G4099,G4370,G564);
  and GNAME4100(G4100,G4370,G560);
  and GNAME4101(G4101,G4370,G554);
  and GNAME4102(G4102,G4370,G557);
  and GNAME4103(G4103,G4370,G555);
  not GNAME4104(G4104,G8728);
  and GNAME4105(G4105,G23043,G4147);
  or GNAME4106(G4106,G3841,G4054);
  and GNAME4107(G4107,G4058,G4054,G4778);
  and GNAME4108(G4108,G4057,G4780);
  nor GNAME4109(G4109,G4057,G4106);
  and GNAME4110(G4110,G4891,G4060);
  and GNAME4111(G4111,G4176,G4170,G5959);
  nand GNAME4112(G4112,G4888,G4062);
  and GNAME4113(G4113,G3681,G4110);
  and GNAME4114(G4114,G4090,G4889);
  and GNAME4115(G4115,G4085,G4889);
  and GNAME4116(G4116,G4892,G4900);
  and GNAME4117(G4117,G4898,G4889);
  and GNAME4118(G4118,G4423,G4060);
  and GNAME4119(G4119,G4889,G4118);
  and GNAME4120(G4120,G4422,G4060);
  and GNAME4121(G4121,G4889,G4120);
  nand GNAME4122(G4122,G4062,G6219,G6220);
  nor GNAME4123(G4123,G4390,G4122);
  and GNAME4124(G4124,G5087,G5081);
  and GNAME4125(G4125,G4118,G5081);
  and GNAME4126(G4126,G4120,G5081);
  nand GNAME4127(G4127,G5239,G4062);
  nor GNAME4128(G4128,G4390,G4127);
  and GNAME4129(G4129,G5087,G5240);
  and GNAME4130(G4130,G4118,G5240);
  and GNAME4131(G4131,G4120,G5240);
  and GNAME4132(G4132,G23043,G4052);
  nor GNAME4133(G4133,G3841,G4132);
  nand GNAME4134(G4134,G5499,G5498);
  or GNAME4135(G4135,G4139,G4138);
  nor GNAME4136(G4136,G4054,G4172);
  nor GNAME4137(G4137,G5944,G4054);
  and GNAME4138(G4138,G4075,G4053,G5489);
  and GNAME4139(G4139,G5489,G4053,G4399);
  and GNAME4140(G4140,G4053,G5496);
  and GNAME4141(G4141,G5525,G5526);
  and GNAME4142(G4142,G5530,G4141,G5529,G5527,G5528);
  nand GNAME4143(G4143,G5691,G4082,G4402);
  and GNAME4144(G4144,G4390,G4080,G4401);
  and GNAME4145(G4145,G4111,G546);
  and GNAME4146(G4146,G4147,G4051,G5065);
  nand GNAME4147(G4147,G5889,G5890);
  nand GNAME4148(G4148,G5894,G5895);
  nand GNAME4149(G4149,G5896,G5897);
  and GNAME4150(G4150,G5892,G5893);
  nand GNAME4151(G4151,G5898,G5899);
  nand GNAME4152(G4152,G5900,G5901);
  nand GNAME4153(G4153,G5902,G5903);
  nand GNAME4154(G4154,G5904,G5905);
  nand GNAME4155(G4155,G5906,G5907);
  nand GNAME4156(G4156,G5908,G5909);
  nand GNAME4157(G4157,G5910,G5911);
  nand GNAME4158(G4158,G5912,G5913);
  nand GNAME4159(G4159,G5914,G5915);
  nand GNAME4160(G4160,G5916,G5917);
  nand GNAME4161(G4161,G5918,G5919);
  nand GNAME4162(G4162,G5920,G5921);
  nand GNAME4163(G4163,G5922,G5923);
  nand GNAME4164(G4164,G5924,G5925);
  nand GNAME4165(G4165,G5926,G5927);
  nand GNAME4166(G4166,G5928,G5929);
  nand GNAME4167(G4167,G5930,G5931);
  nand GNAME4168(G4168,G5932,G5933);
  nand GNAME4169(G4169,G5934,G5935);
  nand GNAME4170(G4170,G5936,G5937);
  nand GNAME4171(G4171,G5939,G5940);
  nand GNAME4172(G4172,G5942,G5943);
  nand GNAME4173(G4173,G5969,G5970);
  nand GNAME4174(G4174,G5972,G5973);
  nand GNAME4175(G4175,G5957,G5958);
  nand GNAME4176(G4176,G5960,G5961);
  nand GNAME4177(G4177,G5975,G5976);
  nand GNAME4178(G4178,G5978,G5979);
  nand GNAME4179(G4179,G5981,G5982);
  nand GNAME4180(G4180,G5984,G5985);
  nand GNAME4181(G4181,G5987,G5988);
  nand GNAME4182(G4182,G5990,G5991);
  nand GNAME4183(G4183,G5993,G5994);
  nand GNAME4184(G4184,G5996,G5997);
  nand GNAME4185(G4185,G5999,G6000);
  nand GNAME4186(G4186,G6002,G6003);
  nand GNAME4187(G4187,G6005,G6006);
  nand GNAME4188(G4188,G6008,G6009);
  nand GNAME4189(G4189,G6011,G6012);
  nand GNAME4190(G4190,G6014,G6015);
  nand GNAME4191(G4191,G6017,G6018);
  nand GNAME4192(G4192,G6020,G6021);
  nand GNAME4193(G4193,G6023,G6024);
  nand GNAME4194(G4194,G6026,G6027);
  nand GNAME4195(G4195,G6029,G6030);
  nand GNAME4196(G4196,G6032,G6033);
  nand GNAME4197(G4197,G6035,G6036);
  nand GNAME4198(G4198,G6146,G6147);
  nand GNAME4199(G4199,G6148,G6149);
  nand GNAME4200(G4200,G6150,G6151);
  nand GNAME4201(G4201,G6152,G6153);
  nand GNAME4202(G4202,G6154,G6155);
  nand GNAME4203(G4203,G6156,G6157);
  nand GNAME4204(G4204,G6158,G6159);
  nand GNAME4205(G4205,G6160,G6161);
  nand GNAME4206(G4206,G6162,G6163);
  nand GNAME4207(G4207,G6164,G6165);
  nand GNAME4208(G4208,G6166,G6167);
  nand GNAME4209(G4209,G6168,G6169);
  nand GNAME4210(G4210,G6170,G6171);
  nand GNAME4211(G4211,G6172,G6173);
  nand GNAME4212(G4212,G6174,G6175);
  nand GNAME4213(G4213,G6176,G6177);
  nand GNAME4214(G4214,G6178,G6179);
  nand GNAME4215(G4215,G6180,G6181);
  nand GNAME4216(G4216,G6182,G6183);
  nand GNAME4217(G4217,G6184,G6185);
  nand GNAME4218(G4218,G6186,G6187);
  nand GNAME4219(G4219,G6188,G6189);
  nand GNAME4220(G4220,G6190,G6191);
  nand GNAME4221(G4221,G6192,G6193);
  nand GNAME4222(G4222,G6194,G6195);
  nand GNAME4223(G4223,G6196,G6197);
  nand GNAME4224(G4224,G6198,G6199);
  nand GNAME4225(G4225,G6200,G6201);
  nand GNAME4226(G4226,G6202,G6203);
  nand GNAME4227(G4227,G6204,G6205);
  nand GNAME4228(G4228,G6206,G6207);
  nand GNAME4229(G4229,G6208,G6209);
  nand GNAME4230(G4230,G6228,G6229);
  nand GNAME4231(G4231,G6230,G6231);
  nand GNAME4232(G4232,G6232,G6233);
  nand GNAME4233(G4233,G6234,G6235);
  nand GNAME4234(G4234,G6236,G6237);
  nand GNAME4235(G4235,G6238,G6239);
  nand GNAME4236(G4236,G6240,G6241);
  nand GNAME4237(G4237,G6242,G6243);
  nand GNAME4238(G4238,G6244,G6245);
  nand GNAME4239(G4239,G6246,G6247);
  nand GNAME4240(G4240,G6248,G6249);
  nand GNAME4241(G4241,G6250,G6251);
  nand GNAME4242(G4242,G6252,G6253);
  nand GNAME4243(G4243,G6254,G6255);
  nand GNAME4244(G4244,G6256,G6257);
  nand GNAME4245(G4245,G6258,G6259);
  nand GNAME4246(G4246,G6260,G6261);
  nand GNAME4247(G4247,G6262,G6263);
  nand GNAME4248(G4248,G6264,G6265);
  nand GNAME4249(G4249,G6266,G6267);
  nand GNAME4250(G4250,G6268,G6269);
  nand GNAME4251(G4251,G6270,G6271);
  nand GNAME4252(G4252,G6272,G6273);
  nand GNAME4253(G4253,G6274,G6275);
  nand GNAME4254(G4254,G6276,G6277);
  nand GNAME4255(G4255,G6278,G6279);
  nand GNAME4256(G4256,G6280,G6281);
  nand GNAME4257(G4257,G6282,G6283);
  nand GNAME4258(G4258,G6284,G6285);
  nand GNAME4259(G4259,G6286,G6287);
  nand GNAME4260(G4260,G6288,G6289);
  nand GNAME4261(G4261,G6290,G6291);
  nand GNAME4262(G4262,G6292,G6293);
  nand GNAME4263(G4263,G6294,G6295);
  nand GNAME4264(G4264,G6296,G6297);
  nand GNAME4265(G4265,G6298,G6299);
  nand GNAME4266(G4266,G6300,G6301);
  nand GNAME4267(G4267,G6302,G6303);
  nand GNAME4268(G4268,G6304,G6305);
  nand GNAME4269(G4269,G6306,G6307);
  nand GNAME4270(G4270,G6308,G6309);
  nand GNAME4271(G4271,G6310,G6311);
  nand GNAME4272(G4272,G6312,G6313);
  nand GNAME4273(G4273,G6314,G6315);
  nand GNAME4274(G4274,G6316,G6317);
  nand GNAME4275(G4275,G6318,G6319);
  nand GNAME4276(G4276,G6320,G6321);
  nand GNAME4277(G4277,G6322,G6323);
  nand GNAME4278(G4278,G6324,G6325);
  nand GNAME4279(G4279,G6326,G6327);
  nand GNAME4280(G4280,G6328,G6329);
  nand GNAME4281(G4281,G6330,G6331);
  nand GNAME4282(G4282,G6332,G6333);
  nand GNAME4283(G4283,G6334,G6335);
  or GNAME4284(G4284,G22839,G22838,G22837,G22836);
  nor GNAME4285(G4285,G4284,G22840,G22841,G22842,G22843);
  or GNAME4286(G4286,G22847,G22846,G22845,G22844);
  nor GNAME4287(G4287,G4286,G22850,G22848,G22849);
  or GNAME4288(G4288,G22854,G22853,G22852,G22851);
  nor GNAME4289(G4289,G4288,G22857,G22855,G22856);
  or GNAME4290(G4290,G22861,G22860,G22859,G22858);
  nor GNAME4291(G4291,G4290,G22864,G22862,G22863);
  and GNAME4292(G4292,G4429,G4818,G4428);
  and GNAME4293(G4293,G4444,G4442,G4439);
  and GNAME4294(G4294,G4462,G4853,G4461);
  and GNAME4295(G4295,G4476,G4474,G4475);
  and GNAME4296(G4296,G4494,G4833,G4493);
  and GNAME4297(G4297,G4512,G4798,G4511);
  and GNAME4298(G4298,G4529,G4878,G4528);
  and GNAME4299(G4299,G4542,G4540,G4541);
  and GNAME4300(G4300,G4555,G4823,G4554);
  and GNAME4301(G4301,G4568,G4788,G4567);
  and GNAME4302(G4302,G4574,G4572,G4573);
  and GNAME4303(G4303,G4582,G4843,G4581);
  and GNAME4304(G4304,G4588,G4586,G4587);
  and GNAME4305(G4305,G4601,G4863,G4600);
  and GNAME4306(G4306,G4609,G4808,G4608);
  and GNAME4307(G4307,G4622,G4868,G4621);
  and GNAME4308(G4308,G4636,G4634,G4635);
  and GNAME4309(G4309,G4654,G4803,G4653);
  and GNAME4310(G4310,G4667,G4828,G4666);
  and GNAME4311(G4311,G4679,G4783,G4678);
  and GNAME4312(G4312,G4694,G4692,G4693);
  and GNAME4313(G4313,G4712,G4848,G4711);
  and GNAME4314(G4314,G4718,G4716,G4717);
  and GNAME4315(G4315,G4726,G4838,G4725);
  and GNAME4316(G4316,G4734,G4793,G4733);
  and GNAME4317(G4317,G4742,G4873,G4741);
  and GNAME4318(G4318,G4750,G4813,G4749);
  and GNAME4319(G4319,G4756,G4754,G4751);
  and GNAME4320(G4320,G4764,G4858,G4763);
  and GNAME4321(G4321,G6042,G6045,G6048,G6051);
  and GNAME4322(G4322,G4321,G6054,G6057,G6060,G6063);
  and GNAME4323(G4323,G6066,G6069,G6072,G6081);
  and GNAME4324(G4324,G4323,G6078,G6075,G6084,G6087);
  and GNAME4325(G4325,G6102,G6105,G6099,G6111);
  and GNAME4326(G4326,G4325,G6090,G6093,G6096,G6108);
  and GNAME4327(G4327,G6114,G6117,G6120,G6123);
  and GNAME4328(G4328,G4327,G6126,G6129,G6132,G6135);
  and GNAME4329(G4329,G4905,G4903,G4904);
  and GNAME4330(G4330,G4911,G4909,G4910);
  and GNAME4331(G4331,G4917,G4915,G4916);
  and GNAME4332(G4332,G4923,G4921,G4922);
  and GNAME4333(G4333,G4929,G4927,G4928);
  and GNAME4334(G4334,G4935,G4933,G4934);
  and GNAME4335(G4335,G4941,G4939,G4940);
  and GNAME4336(G4336,G4947,G4945,G4946);
  and GNAME4337(G4337,G4953,G4951,G4952);
  and GNAME4338(G4338,G4959,G4957,G4958);
  and GNAME4339(G4339,G4965,G4963,G4964);
  and GNAME4340(G4340,G4971,G4969,G4970);
  and GNAME4341(G4341,G4977,G4975,G4976);
  and GNAME4342(G4342,G4983,G4981,G4982);
  and GNAME4343(G4343,G4989,G4987,G4988);
  and GNAME4344(G4344,G4995,G4993,G4994);
  and GNAME4345(G4345,G5001,G4999,G5000);
  and GNAME4346(G4346,G5007,G5005,G5006);
  and GNAME4347(G4347,G5013,G5011,G5012);
  and GNAME4348(G4348,G5019,G5017,G5018);
  and GNAME4349(G4349,G5025,G5023,G5024);
  and GNAME4350(G4350,G5031,G5029,G5030);
  and GNAME4351(G4351,G5037,G5035,G5036);
  and GNAME4352(G4352,G5043,G5041,G5042);
  and GNAME4353(G4353,G5049,G5047,G5048);
  and GNAME4354(G4354,G5055,G5053,G5054);
  and GNAME4355(G4355,G5061,G5059,G5060);
  and GNAME4356(G4356,G5944,G4377);
  nand GNAME4357(G4357,G4068,G4057,G5944);
  nand GNAME4358(G4358,G4322,G4324,G4326,G4328);
  or GNAME4359(G4359,G4171,G4081);
  and GNAME4360(G4360,G3683,G4110);
  and GNAME4361(G4361,G6215,G6216);
  and GNAME4362(G4362,G6217,G6218);
  and GNAME4363(G4363,G5962,G5941);
  and GNAME4364(G4364,G4063,G4062);
  not GNAME4365(G4365,G4106);
  not GNAME4366(G4366,G4062);
  not GNAME4367(G4367,G4060);
  not GNAME4368(G4368,G4082);
  not GNAME4369(G4369,G4111);
  not GNAME4370(G4370,G4356);
  nand GNAME4371(G4371,G5953,G6396);
  nand GNAME4372(G4372,G4113,G5240);
  nand GNAME4373(G4373,G4113,G5081);
  not GNAME4374(G4374,G4105);
  not GNAME4375(G4375,G4079);
  not GNAME4376(G4376,G4086);
  not GNAME4377(G4377,G4057);
  nand GNAME4378(G4378,G4370,G4147);
  nand GNAME4379(G4379,G4053,G4367,G4370);
  nand GNAME4380(G4380,G5947,G22905);
  nand GNAME4381(G4381,G5950,G22937);
  nand GNAME4382(G4382,G5953,G9378);
  nand GNAME4383(G4383,G5956,G22873);
  not GNAME4384(G4384,G3727);
  nand GNAME4385(G4385,G5947,G22903);
  nand GNAME4386(G4386,G5950,G22935);
  nand GNAME4387(G4387,G5953,G9374);
  nand GNAME4388(G4388,G5956,G22871);
  not GNAME4389(G4389,G3731);
  not GNAME4390(G4390,G4076);
  nand GNAME4391(G4391,G5959,G4076);
  nand GNAME4392(G4392,G5941,G4078);
  not GNAME4393(G4393,G4063);
  nand GNAME4394(G4394,G4285,G4287,G4289,G4291);
  nand GNAME4395(G4395,G4394,G4393);
  nand GNAME4396(G4396,G4393,G22835);
  or GNAME4397(G4397,G4148,G4149);
  or GNAME4398(G4398,G4148,G4150);
  not GNAME4399(G4399,G4075);
  not GNAME4400(G4400,G4067);
  nand GNAME4401(G4401,G4170,G4079);
  nand GNAME4402(G4402,G5938,G4171,G4059);
  or GNAME4403(G4403,G4051,G5941);
  or GNAME4404(G4404,G4176,G4080);
  nand GNAME4405(G4405,G5938,G4368);
  nand GNAME4406(G4406,G4400,G4376);
  nand GNAME4407(G4407,G4084,G4087);
  nand GNAME4408(G4408,G4406,G4407);
  nand GNAME4409(G4409,G4153,G4177);
  nand GNAME4410(G4410,G5978,G4409);
  not GNAME4411(G4411,G4061);
  nor GNAME4412(G4412,G4084,G4085);
  or GNAME4413(G4413,G4087,G4412);
  nand GNAME4414(G4414,G4067,G4376);
  or GNAME4415(G4415,G4059,G4367);
  nand GNAME4416(G4416,G4415,G4413,G4414);
  nand GNAME4417(G4417,G4416,G4062);
  nand GNAME4418(G4418,G4067,G4068);
  nand GNAME4419(G4419,G4106,G4374,G4417,G4418);
  nand GNAME4420(G4420,G22828,G4065);
  nand GNAME4421(G4421,G8894,G4066);
  nand GNAME4422(G4422,G5977,G4073);
  nand GNAME4423(G4423,G5963,G5964,G5965,G5966);
  nand GNAME4424(G4424,G3731,G4072);
  nand GNAME4425(G4425,G3727,G4074);
  nand GNAME4426(G4426,G4419,G9384);
  nand GNAME4427(G4427,G8992,G4088);
  nand GNAME4428(G4428,G4410,G4089);
  nand GNAME4429(G4429,G4178,G4091);
  nand GNAME4430(G4430,G5953,G9395);
  nand GNAME4431(G4431,G5956,G22893);
  nand GNAME4432(G4432,G5947,G22925);
  nand GNAME4433(G4433,G5950,G22957);
  nand GNAME4434(G4434,G5953,G9393);
  nand GNAME4435(G4435,G5956,G22891);
  nand GNAME4436(G4436,G5947,G22923);
  nand GNAME4437(G4437,G5950,G22955);
  or GNAME4438(G4438,G4091,G4089);
  nand GNAME4439(G4439,G3691,G4072);
  nand GNAME4440(G4440,G3687,G4074);
  nand GNAME4441(G4441,G4419,G9389);
  nand GNAME4442(G4442,G3841,G23041);
  nand GNAME4443(G4443,G4088,G9048);
  nand GNAME4444(G4444,G4438,G4092);
  nand GNAME4445(G4445,G5947,G22912);
  nand GNAME4446(G4446,G5950,G22944);
  nand GNAME4447(G4447,G5953,G9387);
  nand GNAME4448(G4448,G5956,G22880);
  not GNAME4449(G4449,G3713);
  nand GNAME4450(G4450,G5947,G22910);
  nand GNAME4451(G4451,G5950,G22942);
  nand GNAME4452(G4452,G5953,G9391);
  nand GNAME4453(G4453,G5956,G22878);
  not GNAME4454(G4454,G3717);
  nand GNAME4455(G4455,G4164,G4177);
  nand GNAME4456(G4456,G5981,G4455);
  nand GNAME4457(G4457,G3717,G4072);
  nand GNAME4458(G4458,G3713,G4074);
  nand GNAME4459(G4459,G4419,G9397);
  nand GNAME4460(G4460,G4088,G8996);
  nand GNAME4461(G4461,G4456,G4089);
  nand GNAME4462(G4462,G4179,G4091);
  nand GNAME4463(G4463,G5953,G9376);
  nand GNAME4464(G4464,G5956,G22889);
  nand GNAME4465(G4465,G5947,G22921);
  nand GNAME4466(G4466,G5950,G22953);
  nand GNAME4467(G4467,G5953,G9383);
  nand GNAME4468(G4468,G5956,G22887);
  nand GNAME4469(G4469,G5947,G22919);
  nand GNAME4470(G4470,G5950,G22951);
  nand GNAME4471(G4471,G3699,G4072);
  nand GNAME4472(G4472,G3695,G4074);
  nand GNAME4473(G4473,G4419,G9372);
  nand GNAME4474(G4474,G3841,G23039);
  nand GNAME4475(G4475,G4088,G9060);
  nand GNAME4476(G4476,G4438,G4093);
  nand GNAME4477(G4477,G5947,G22908);
  nand GNAME4478(G4478,G5950,G22940);
  nand GNAME4479(G4479,G5953,G9375);
  nand GNAME4480(G4480,G5956,G22876);
  not GNAME4481(G4481,G3721);
  nand GNAME4482(G4482,G5947,G22906);
  nand GNAME4483(G4483,G5950,G22938);
  nand GNAME4484(G4484,G5953,G9380);
  nand GNAME4485(G4485,G5956,G22874);
  not GNAME4486(G4486,G3725);
  nand GNAME4487(G4487,G4168,G4177);
  nand GNAME4488(G4488,G5984,G4487);
  nand GNAME4489(G4489,G3725,G4072);
  nand GNAME4490(G4490,G3721,G4074);
  nand GNAME4491(G4491,G4419,G9379);
  nand GNAME4492(G4492,G4088,G8953);
  nand GNAME4493(G4493,G4488,G4089);
  nand GNAME4494(G4494,G4180,G4091);
  nand GNAME4495(G4495,G5947,G22901);
  nand GNAME4496(G4496,G5950,G22933);
  nand GNAME4497(G4497,G5953,G9396);
  nand GNAME4498(G4498,G5956,G22869);
  not GNAME4499(G4499,G3735);
  nand GNAME4500(G4500,G5947,G22899);
  nand GNAME4501(G4501,G5950,G22931);
  nand GNAME4502(G4502,G5953,G23018);
  nand GNAME4503(G4503,G5956,G22867);
  not GNAME4504(G4504,G3739);
  nand GNAME4505(G4505,G4157,G4177);
  nand GNAME4506(G4506,G5987,G4505);
  nand GNAME4507(G4507,G3739,G4072);
  nand GNAME4508(G4508,G3735,G4074);
  nand GNAME4509(G4509,G4419,G9392);
  nand GNAME4510(G4510,G4088,G8993);
  nand GNAME4511(G4511,G4506,G4089);
  nand GNAME4512(G4512,G4181,G4091);
  nand GNAME4513(G4513,G5953,G9386);
  nand GNAME4514(G4514,G5956,G22885);
  nand GNAME4515(G4515,G5947,G22917);
  nand GNAME4516(G4516,G5950,G22949);
  nand GNAME4517(G4517,G5947,G22915);
  nand GNAME4518(G4518,G5950,G22947);
  nand GNAME4519(G4519,G5953,G9377);
  nand GNAME4520(G4520,G5956,G22883);
  not GNAME4521(G4521,G3707);
  nand GNAME4522(G4522,G4175,G4177);
  nand GNAME4523(G4523,G5990,G4522);
  nand GNAME4524(G4524,G3707,G4072);
  nand GNAME4525(G4525,G3703,G4074);
  nand GNAME4526(G4526,G4419,G9381);
  nand GNAME4527(G4527,G4088,G9075);
  nand GNAME4528(G4528,G4523,G4089);
  nand GNAME4529(G4529,G4182,G4091);
  nand GNAME4530(G4530,G5956,G22894);
  nand GNAME4531(G4531,G5947,G22926);
  nand GNAME4532(G4532,G5950,G22958);
  nand GNAME4533(G4533,G5953,G9389);
  nand GNAME4534(G4534,G5956,G22892);
  nand GNAME4535(G4535,G5947,G22924);
  nand GNAME4536(G4536,G5950,G22956);
  nand GNAME4537(G4537,G3689,G4072);
  nand GNAME4538(G4538,G3685,G4074);
  nand GNAME4539(G4539,G4419,G9395);
  nand GNAME4540(G4540,G3841,G23035);
  nand GNAME4541(G4541,G4088,G9045);
  nand GNAME4542(G4542,G4438,G4094);
  nand GNAME4543(G4543,G5947,G22904);
  nand GNAME4544(G4544,G5950,G22936);
  nand GNAME4545(G4545,G5953,G9384);
  nand GNAME4546(G4546,G5956,G22872);
  not GNAME4547(G4547,G3729);
  nand GNAME4548(G4548,G4152,G4177);
  nand GNAME4549(G4549,G5993,G4548);
  nand GNAME4550(G4550,G3729,G4072);
  nand GNAME4551(G4551,G3725,G4074);
  nand GNAME4552(G4552,G4419,G9378);
  nand GNAME4553(G4553,G4088,G9011);
  nand GNAME4554(G4554,G4549,G4089);
  nand GNAME4555(G4555,G4183,G4091);
  nand GNAME4556(G4556,G5956,G22865);
  nand GNAME4557(G4557,G5947,G22897);
  nand GNAME4558(G4558,G5950,G22929);
  nand GNAME4559(G4559,G5953,G23023);
  not GNAME4560(G4560,G3743);
  nand GNAME4561(G4561,G4159,G4177);
  nand GNAME4562(G4562,G5996,G4561);
  nand GNAME4563(G4563,G3743,G4072);
  nand GNAME4564(G4564,G3739,G4074);
  nand GNAME4565(G4565,G4419,G23033);
  nand GNAME4566(G4566,G4088,G9072);
  nand GNAME4567(G4567,G4562,G4089);
  nand GNAME4568(G4568,G4184,G4091);
  nand GNAME4569(G4569,G3703,G4072);
  nand GNAME4570(G4570,G3699,G4074);
  nand GNAME4571(G4571,G4419,G9394);
  nand GNAME4572(G4572,G3841,G23032);
  nand GNAME4573(G4573,G4088,G9066);
  nand GNAME4574(G4574,G4438,G4095);
  nand GNAME4575(G4575,G4166,G4177);
  nand GNAME4576(G4576,G5999,G4575);
  nand GNAME4577(G4577,G3721,G4072);
  nand GNAME4578(G4578,G3717,G4074);
  nand GNAME4579(G4579,G4419,G9390);
  nand GNAME4580(G4580,G4088,G9094);
  nand GNAME4581(G4581,G4576,G4089);
  nand GNAME4582(G4582,G4185,G4091);
  nand GNAME4583(G4583,G3695,G4072);
  nand GNAME4584(G4584,G3691,G4074);
  nand GNAME4585(G4585,G4419,G9382);
  nand GNAME4586(G4586,G3841,G23030);
  nand GNAME4587(G4587,G4088,G9054);
  nand GNAME4588(G4588,G4438,G4096);
  nand GNAME4589(G4589,G5947,G22914);
  nand GNAME4590(G4590,G5950,G22946);
  nand GNAME4591(G4591,G5953,G9385);
  nand GNAME4592(G4592,G5956,G22882);
  not GNAME4593(G4593,G3709);
  nand GNAME4594(G4594,G4162,G4177);
  nand GNAME4595(G4595,G6002,G4594);
  nand GNAME4596(G4596,G3713,G4072);
  nand GNAME4597(G4597,G3709,G4074);
  nand GNAME4598(G4598,G4419,G9373);
  nand GNAME4599(G4599,G4088,G9084);
  nand GNAME4600(G4600,G4595,G4089);
  nand GNAME4601(G4601,G4186,G4091);
  nand GNAME4602(G4602,G4155,G4177);
  nand GNAME4603(G4603,G6005,G4602);
  nand GNAME4604(G4604,G3735,G4072);
  nand GNAME4605(G4605,G3731,G4074);
  nand GNAME4606(G4606,G4419,G9388);
  nand GNAME4607(G4607,G4088,G9015);
  nand GNAME4608(G4608,G4603,G4089);
  nand GNAME4609(G4609,G4187,G4091);
  nand GNAME4610(G4610,G5947,G22913);
  nand GNAME4611(G4611,G5950,G22945);
  nand GNAME4612(G4612,G5953,G9373);
  nand GNAME4613(G4613,G5956,G22881);
  not GNAME4614(G4614,G3711);
  nand GNAME4615(G4615,G4161,G4177);
  nand GNAME4616(G4616,G6008,G4615);
  nand GNAME4617(G4617,G3711,G4072);
  nand GNAME4618(G4618,G3707,G4074);
  nand GNAME4619(G4619,G4419,G9385);
  nand GNAME4620(G4620,G4088,G9081);
  nand GNAME4621(G4621,G4616,G4089);
  nand GNAME4622(G4622,G4188,G4091);
  nand GNAME4623(G4623,G5953,G9382);
  nand GNAME4624(G4624,G5956,G22890);
  nand GNAME4625(G4625,G5947,G22922);
  nand GNAME4626(G4626,G5950,G22954);
  nand GNAME4627(G4627,G5953,G9372);
  nand GNAME4628(G4628,G5956,G22888);
  nand GNAME4629(G4629,G5947,G22920);
  nand GNAME4630(G4630,G5950,G22952);
  nand GNAME4631(G4631,G3697,G4072);
  nand GNAME4632(G4632,G3693,G4074);
  nand GNAME4633(G4633,G4419,G9376);
  nand GNAME4634(G4634,G3841,G23026);
  nand GNAME4635(G4635,G4088,G9057);
  nand GNAME4636(G4636,G4438,G4097);
  nand GNAME4637(G4637,G5947,G22902);
  nand GNAME4638(G4638,G5950,G22934);
  nand GNAME4639(G4639,G5953,G9388);
  nand GNAME4640(G4640,G5956,G22870);
  not GNAME4641(G4641,G3733);
  nand GNAME4642(G4642,G5947,G22900);
  nand GNAME4643(G4643,G5950,G22932);
  nand GNAME4644(G4644,G5953,G9392);
  nand GNAME4645(G4645,G5956,G22868);
  not GNAME4646(G4646,G3737);
  nand GNAME4647(G4647,G4156,G4177);
  nand GNAME4648(G4648,G6011,G4647);
  nand GNAME4649(G4649,G3737,G4072);
  nand GNAME4650(G4650,G3733,G4074);
  nand GNAME4651(G4651,G4419,G9396);
  nand GNAME4652(G4652,G4088,G9018);
  nand GNAME4653(G4653,G4648,G4089);
  nand GNAME4654(G4654,G4189,G4091);
  nand GNAME4655(G4655,G5947,G22907);
  nand GNAME4656(G4656,G5950,G22939);
  nand GNAME4657(G4657,G5953,G9379);
  nand GNAME4658(G4658,G5956,G22875);
  not GNAME4659(G4659,G3723);
  nand GNAME4660(G4660,G4151,G4177);
  nand GNAME4661(G4661,G6014,G4660);
  nand GNAME4662(G4662,G3727,G4072);
  nand GNAME4663(G4663,G3723,G4074);
  nand GNAME4664(G4664,G4419,G9380);
  nand GNAME4665(G4665,G4088,G9008);
  nand GNAME4666(G4666,G4661,G4089);
  nand GNAME4667(G4667,G4190,G4091);
  nand GNAME4668(G4668,G5956,G22866);
  nand GNAME4669(G4669,G5947,G22898);
  nand GNAME4670(G4670,G5950,G22930);
  nand GNAME4671(G4671,G5953,G23033);
  not GNAME4672(G4672,G3741);
  nand GNAME4673(G4673,G4169,G4177);
  nand GNAME4674(G4674,G6017,G4673);
  nand GNAME4675(G4675,G3741,G4074);
  nand GNAME4676(G4676,G4419,G23023);
  nand GNAME4677(G4677,G4088,G8991);
  nand GNAME4678(G4678,G4674,G4089);
  nand GNAME4679(G4679,G4191,G4091);
  nand GNAME4680(G4680,G5953,G9394);
  nand GNAME4681(G4681,G5956,G22886);
  nand GNAME4682(G4682,G5947,G22918);
  nand GNAME4683(G4683,G5950,G22950);
  nand GNAME4684(G4684,G5947,G22916);
  nand GNAME4685(G4685,G5950,G22948);
  nand GNAME4686(G4686,G5953,G9381);
  nand GNAME4687(G4687,G5956,G22884);
  not GNAME4688(G4688,G3705);
  nand GNAME4689(G4689,G3705,G4072);
  nand GNAME4690(G4690,G3701,G4074);
  nand GNAME4691(G4691,G4419,G9386);
  nand GNAME4692(G4692,G3841,G23022);
  nand GNAME4693(G4693,G4088,G9069);
  nand GNAME4694(G4694,G4438,G4098);
  nand GNAME4695(G4695,G5947,G22911);
  nand GNAME4696(G4696,G5950,G22943);
  nand GNAME4697(G4697,G5953,G9397);
  nand GNAME4698(G4698,G5956,G22879);
  not GNAME4699(G4699,G3715);
  nand GNAME4700(G4700,G5947,G22909);
  nand GNAME4701(G4701,G5950,G22941);
  nand GNAME4702(G4702,G5953,G9390);
  nand GNAME4703(G4703,G5956,G22877);
  not GNAME4704(G4704,G3719);
  nand GNAME4705(G4705,G4165,G4177);
  nand GNAME4706(G4706,G6020,G4705);
  nand GNAME4707(G4707,G3719,G4072);
  nand GNAME4708(G4708,G3715,G4074);
  nand GNAME4709(G4709,G4419,G9391);
  nand GNAME4710(G4710,G4088,G9091);
  nand GNAME4711(G4711,G4706,G4089);
  nand GNAME4712(G4712,G4192,G4091);
  nand GNAME4713(G4713,G3701,G4072);
  nand GNAME4714(G4714,G3697,G4074);
  nand GNAME4715(G4715,G4419,G9383);
  nand GNAME4716(G4716,G3841,G23020);
  nand GNAME4717(G4717,G4088,G9063);
  nand GNAME4718(G4718,G4438,G4099);
  nand GNAME4719(G4719,G4167,G4177);
  nand GNAME4720(G4720,G6023,G4719);
  nand GNAME4721(G4721,G3723,G4072);
  nand GNAME4722(G4722,G3719,G4074);
  nand GNAME4723(G4723,G4419,G9375);
  nand GNAME4724(G4724,G4088,G8997);
  nand GNAME4725(G4725,G4720,G4089);
  nand GNAME4726(G4726,G4193,G4091);
  nand GNAME4727(G4727,G4158,G4177);
  nand GNAME4728(G4728,G6026,G4727);
  nand GNAME4729(G4729,G3741,G4072);
  nand GNAME4730(G4730,G3737,G4074);
  nand GNAME4731(G4731,G4419,G23018);
  nand GNAME4732(G4732,G4088,G8954);
  nand GNAME4733(G4733,G4728,G4089);
  nand GNAME4734(G4734,G4194,G4091);
  nand GNAME4735(G4735,G4160,G4177);
  nand GNAME4736(G4736,G6029,G4735);
  nand GNAME4737(G4737,G3709,G4072);
  nand GNAME4738(G4738,G3705,G4074);
  nand GNAME4739(G4739,G4419,G9377);
  nand GNAME4740(G4740,G4088,G9078);
  nand GNAME4741(G4741,G4736,G4089);
  nand GNAME4742(G4742,G4195,G4091);
  nand GNAME4743(G4743,G4154,G4177);
  nand GNAME4744(G4744,G6032,G4743);
  nand GNAME4745(G4745,G3733,G4072);
  nand GNAME4746(G4746,G3729,G4074);
  nand GNAME4747(G4747,G4419,G9374);
  nand GNAME4748(G4748,G4088,G8955);
  nand GNAME4749(G4749,G4744,G4089);
  nand GNAME4750(G4750,G4196,G4091);
  nand GNAME4751(G4751,G3693,G4072);
  nand GNAME4752(G4752,G3689,G4074);
  nand GNAME4753(G4753,G4419,G9393);
  nand GNAME4754(G4754,G3841,G23015);
  nand GNAME4755(G4755,G4088,G9051);
  nand GNAME4756(G4756,G4438,G4100);
  nand GNAME4757(G4757,G4163,G4177);
  nand GNAME4758(G4758,G6035,G4757);
  nand GNAME4759(G4759,G3715,G4072);
  nand GNAME4760(G4760,G3711,G4074);
  nand GNAME4761(G4761,G4419,G9387);
  nand GNAME4762(G4762,G4088,G9087);
  nand GNAME4763(G4763,G4758,G4089);
  nand GNAME4764(G4764,G4197,G4091);
  nand GNAME4765(G4765,G5938,G4105);
  nand GNAME4766(G4766,G5956,G22896);
  nand GNAME4767(G4767,G5947,G22928);
  nand GNAME4768(G4768,G5950,G22960);
  nand GNAME4769(G4769,G5956,G22895);
  nand GNAME4770(G4770,G5947,G22927);
  nand GNAME4771(G4771,G5950,G22959);
  not GNAME4772(G4772,G4358);
  nand GNAME4773(G4773,G4060,G8728);
  nand GNAME4774(G4774,G5959,G6142,G6143);
  nand GNAME4775(G4775,G6136,G6137,G4774,G6144,G6145);
  nand GNAME4776(G4776,G23043,G4358,G4147,G4376);
  nand GNAME4777(G4777,G4775,G4105);
  nand GNAME4778(G4778,G4367,G4370);
  or GNAME4779(G4779,G4107,G4366);
  nand GNAME4780(G4780,G4779,G4374);
  and GNAME4781(G4781,G4374,G4366);
  nand GNAME4782(G4782,G4107,G22980);
  nand GNAME4783(G4783,G3841,G23023);
  nand GNAME4784(G4784,G8485,G4108);
  nand GNAME4785(G4785,G4169,G6212);
  nand GNAME4786(G4786,G8991,G4109);
  nand GNAME4787(G4787,G4107,G22979);
  nand GNAME4788(G4788,G3841,G23033);
  nand GNAME4789(G4789,G4108,G8539);
  nand GNAME4790(G4790,G4159,G6212);
  nand GNAME4791(G4791,G9072,G4109);
  nand GNAME4792(G4792,G4107,G22978);
  nand GNAME4793(G4793,G3841,G23018);
  nand GNAME4794(G4794,G4108,G8547);
  nand GNAME4795(G4795,G4158,G6212);
  nand GNAME4796(G4796,G8954,G4109);
  nand GNAME4797(G4797,G4107,G22977);
  nand GNAME4798(G4798,G3841,G23037);
  nand GNAME4799(G4799,G4108,G8546);
  nand GNAME4800(G4800,G4157,G6212);
  nand GNAME4801(G4801,G8993,G4109);
  nand GNAME4802(G4802,G4107,G22976);
  nand GNAME4803(G4803,G3841,G23025);
  nand GNAME4804(G4804,G4108,G8545);
  nand GNAME4805(G4805,G4156,G6212);
  nand GNAME4806(G4806,G9018,G4109);
  nand GNAME4807(G4807,G4107,G22975);
  nand GNAME4808(G4808,G3841,G23028);
  nand GNAME4809(G4809,G4108,G8544);
  nand GNAME4810(G4810,G4155,G6212);
  nand GNAME4811(G4811,G9015,G4109);
  nand GNAME4812(G4812,G4107,G22974);
  nand GNAME4813(G4813,G3841,G23016);
  nand GNAME4814(G4814,G4108,G8543);
  nand GNAME4815(G4815,G4154,G6212);
  nand GNAME4816(G4816,G8955,G4109);
  nand GNAME4817(G4817,G4107,G22973);
  nand GNAME4818(G4818,G3841,G23042);
  nand GNAME4819(G4819,G4108,G8542);
  nand GNAME4820(G4820,G4153,G6212);
  nand GNAME4821(G4821,G8992,G4109);
  nand GNAME4822(G4822,G4107,G22972);
  nand GNAME4823(G4823,G3841,G23034);
  nand GNAME4824(G4824,G4108,G8541);
  nand GNAME4825(G4825,G4152,G6212);
  nand GNAME4826(G4826,G9011,G4109);
  nand GNAME4827(G4827,G4107,G22971);
  nand GNAME4828(G4828,G3841,G23024);
  nand GNAME4829(G4829,G4108,G8540);
  nand GNAME4830(G4830,G4151,G6212);
  nand GNAME4831(G4831,G9008,G4109);
  nand GNAME4832(G4832,G4107,G22970);
  nand GNAME4833(G4833,G3841,G23038);
  nand GNAME4834(G4834,G4108,G8556);
  nand GNAME4835(G4835,G4168,G6212);
  nand GNAME4836(G4836,G8953,G4109);
  nand GNAME4837(G4837,G4107,G22969);
  nand GNAME4838(G4838,G3841,G23019);
  nand GNAME4839(G4839,G4108,G8555);
  nand GNAME4840(G4840,G4167,G6212);
  nand GNAME4841(G4841,G8997,G4109);
  nand GNAME4842(G4842,G4107,G22968);
  nand GNAME4843(G4843,G3841,G23031);
  nand GNAME4844(G4844,G4108,G8554);
  nand GNAME4845(G4845,G4166,G6212);
  nand GNAME4846(G4846,G9094,G4109);
  nand GNAME4847(G4847,G4107,G22967);
  nand GNAME4848(G4848,G3841,G23021);
  nand GNAME4849(G4849,G4108,G8553);
  nand GNAME4850(G4850,G4165,G6212);
  nand GNAME4851(G4851,G9091,G4109);
  nand GNAME4852(G4852,G4107,G22966);
  nand GNAME4853(G4853,G3841,G23040);
  nand GNAME4854(G4854,G4108,G8552);
  nand GNAME4855(G4855,G4164,G6212);
  nand GNAME4856(G4856,G8996,G4109);
  nand GNAME4857(G4857,G4107,G22965);
  nand GNAME4858(G4858,G3841,G23014);
  nand GNAME4859(G4859,G4108,G8551);
  nand GNAME4860(G4860,G4163,G6212);
  nand GNAME4861(G4861,G9087,G4109);
  nand GNAME4862(G4862,G4107,G22964);
  nand GNAME4863(G4863,G3841,G23029);
  nand GNAME4864(G4864,G4108,G8550);
  nand GNAME4865(G4865,G4162,G6212);
  nand GNAME4866(G4866,G9084,G4109);
  nand GNAME4867(G4867,G4107,G22963);
  nand GNAME4868(G4868,G3841,G23027);
  nand GNAME4869(G4869,G4108,G8549);
  nand GNAME4870(G4870,G4161,G6212);
  nand GNAME4871(G4871,G9081,G4109);
  nand GNAME4872(G4872,G4107,G22962);
  nand GNAME4873(G4873,G3841,G23017);
  nand GNAME4874(G4874,G4108,G8548);
  nand GNAME4875(G4875,G4160,G6212);
  nand GNAME4876(G4876,G9078,G4109);
  nand GNAME4877(G4877,G4107,G22961);
  nand GNAME4878(G4878,G3841,G23036);
  nand GNAME4879(G4879,G4175,G6212);
  nand GNAME4880(G4880,G4108,G8484);
  nand GNAME4881(G4881,G9075,G4109);
  nand GNAME4882(G4882,G5959,G4176);
  nand GNAME4883(G4883,G4882,G5941);
  nand GNAME4884(G4884,G4883,G4170);
  nand GNAME4885(G4885,G5941,G4111);
  nand GNAME4886(G4886,G4885,G4411);
  and GNAME4887(G4887,G4064,G6213,G6214);
  or GNAME4888(G4888,G4887,G4090);
  not GNAME4889(G4889,G4112);
  or GNAME4890(G4890,G23013,G4073);
  nand GNAME4891(G4891,G4890,G5977);
  nand GNAME4892(G4892,G4889,G4113);
  nand GNAME4893(G4893,G4112,G22960);
  nand GNAME4894(G4894,G4101,G4115);
  nand GNAME4895(G4895,G4112,G22959);
  nand GNAME4896(G4896,G4103,G4115);
  or GNAME4897(G4897,G4076,G4059);
  nand GNAME4898(G4898,G4897,G4083);
  nand GNAME4899(G4899,G9042,G4117);
  nand GNAME4900(G4900,G6396,G4114);
  nand GNAME4901(G4901,G3687,G4119);
  nand GNAME4902(G4902,G4102,G4115);
  nand GNAME4903(G4903,G9045,G4117);
  nand GNAME4904(G4904,G9395,G4114);
  nand GNAME4905(G4905,G4112,G22957);
  nand GNAME4906(G4906,G3689,G4119);
  nand GNAME4907(G4907,G4094,G4115);
  nand GNAME4908(G4908,G3685,G4121);
  nand GNAME4909(G4909,G9048,G4117);
  nand GNAME4910(G4910,G9389,G4114);
  nand GNAME4911(G4911,G4112,G22956);
  nand GNAME4912(G4912,G3691,G4119);
  nand GNAME4913(G4913,G4092,G4115);
  nand GNAME4914(G4914,G3687,G4121);
  nand GNAME4915(G4915,G9051,G4117);
  nand GNAME4916(G4916,G9393,G4114);
  nand GNAME4917(G4917,G4112,G22955);
  nand GNAME4918(G4918,G3693,G4119);
  nand GNAME4919(G4919,G4100,G4115);
  nand GNAME4920(G4920,G3689,G4121);
  nand GNAME4921(G4921,G9054,G4117);
  nand GNAME4922(G4922,G9382,G4114);
  nand GNAME4923(G4923,G4112,G22954);
  nand GNAME4924(G4924,G3695,G4119);
  nand GNAME4925(G4925,G4096,G4115);
  nand GNAME4926(G4926,G3691,G4121);
  nand GNAME4927(G4927,G9057,G4117);
  nand GNAME4928(G4928,G9376,G4114);
  nand GNAME4929(G4929,G4112,G22953);
  nand GNAME4930(G4930,G3697,G4119);
  nand GNAME4931(G4931,G4097,G4115);
  nand GNAME4932(G4932,G3693,G4121);
  nand GNAME4933(G4933,G9060,G4117);
  nand GNAME4934(G4934,G9372,G4114);
  nand GNAME4935(G4935,G4112,G22952);
  nand GNAME4936(G4936,G3699,G4119);
  nand GNAME4937(G4937,G4093,G4115);
  nand GNAME4938(G4938,G3695,G4121);
  nand GNAME4939(G4939,G9063,G4117);
  nand GNAME4940(G4940,G9383,G4114);
  nand GNAME4941(G4941,G4112,G22951);
  nand GNAME4942(G4942,G3701,G4119);
  nand GNAME4943(G4943,G4099,G4115);
  nand GNAME4944(G4944,G3697,G4121);
  nand GNAME4945(G4945,G9066,G4117);
  nand GNAME4946(G4946,G9394,G4114);
  nand GNAME4947(G4947,G4112,G22950);
  nand GNAME4948(G4948,G3703,G4119);
  nand GNAME4949(G4949,G4095,G4115);
  nand GNAME4950(G4950,G3699,G4121);
  nand GNAME4951(G4951,G9069,G4117);
  nand GNAME4952(G4952,G9386,G4114);
  nand GNAME4953(G4953,G4112,G22949);
  nand GNAME4954(G4954,G3705,G4119);
  nand GNAME4955(G4955,G4098,G4115);
  nand GNAME4956(G4956,G3701,G4121);
  nand GNAME4957(G4957,G9075,G4117);
  nand GNAME4958(G4958,G4523,G4115);
  nand GNAME4959(G4959,G4112,G22948);
  nand GNAME4960(G4960,G9381,G4114);
  nand GNAME4961(G4961,G3707,G4119);
  nand GNAME4962(G4962,G3703,G4121);
  nand GNAME4963(G4963,G9078,G4117);
  nand GNAME4964(G4964,G4736,G4115);
  nand GNAME4965(G4965,G4112,G22947);
  nand GNAME4966(G4966,G9377,G4114);
  nand GNAME4967(G4967,G3709,G4119);
  nand GNAME4968(G4968,G3705,G4121);
  nand GNAME4969(G4969,G9081,G4117);
  nand GNAME4970(G4970,G4616,G4115);
  nand GNAME4971(G4971,G4112,G22946);
  nand GNAME4972(G4972,G9385,G4114);
  nand GNAME4973(G4973,G3711,G4119);
  nand GNAME4974(G4974,G3707,G4121);
  nand GNAME4975(G4975,G9084,G4117);
  nand GNAME4976(G4976,G4595,G4115);
  nand GNAME4977(G4977,G4112,G22945);
  nand GNAME4978(G4978,G9373,G4114);
  nand GNAME4979(G4979,G3713,G4119);
  nand GNAME4980(G4980,G3709,G4121);
  nand GNAME4981(G4981,G9087,G4117);
  nand GNAME4982(G4982,G4758,G4115);
  nand GNAME4983(G4983,G4112,G22944);
  nand GNAME4984(G4984,G9387,G4114);
  nand GNAME4985(G4985,G3715,G4119);
  nand GNAME4986(G4986,G3711,G4121);
  nand GNAME4987(G4987,G8996,G4117);
  nand GNAME4988(G4988,G4456,G4115);
  nand GNAME4989(G4989,G4112,G22943);
  nand GNAME4990(G4990,G9397,G4114);
  nand GNAME4991(G4991,G3717,G4119);
  nand GNAME4992(G4992,G3713,G4121);
  nand GNAME4993(G4993,G9091,G4117);
  nand GNAME4994(G4994,G4706,G4115);
  nand GNAME4995(G4995,G4112,G22942);
  nand GNAME4996(G4996,G9391,G4114);
  nand GNAME4997(G4997,G3719,G4119);
  nand GNAME4998(G4998,G3715,G4121);
  nand GNAME4999(G4999,G9094,G4117);
  nand GNAME5000(G5000,G4576,G4115);
  nand GNAME5001(G5001,G4112,G22941);
  nand GNAME5002(G5002,G9390,G4114);
  nand GNAME5003(G5003,G3721,G4119);
  nand GNAME5004(G5004,G3717,G4121);
  nand GNAME5005(G5005,G8997,G4117);
  nand GNAME5006(G5006,G4720,G4115);
  nand GNAME5007(G5007,G4112,G22940);
  nand GNAME5008(G5008,G9375,G4114);
  nand GNAME5009(G5009,G3723,G4119);
  nand GNAME5010(G5010,G3719,G4121);
  nand GNAME5011(G5011,G8953,G4117);
  nand GNAME5012(G5012,G4488,G4115);
  nand GNAME5013(G5013,G4112,G22939);
  nand GNAME5014(G5014,G9379,G4114);
  nand GNAME5015(G5015,G3725,G4119);
  nand GNAME5016(G5016,G3721,G4121);
  nand GNAME5017(G5017,G9008,G4117);
  nand GNAME5018(G5018,G4661,G4115);
  nand GNAME5019(G5019,G4112,G22938);
  nand GNAME5020(G5020,G9380,G4114);
  nand GNAME5021(G5021,G3727,G4119);
  nand GNAME5022(G5022,G3723,G4121);
  nand GNAME5023(G5023,G9011,G4117);
  nand GNAME5024(G5024,G4549,G4115);
  nand GNAME5025(G5025,G4112,G22937);
  nand GNAME5026(G5026,G9378,G4114);
  nand GNAME5027(G5027,G3729,G4119);
  nand GNAME5028(G5028,G3725,G4121);
  nand GNAME5029(G5029,G8992,G4117);
  nand GNAME5030(G5030,G4410,G4115);
  nand GNAME5031(G5031,G4112,G22936);
  nand GNAME5032(G5032,G9384,G4114);
  nand GNAME5033(G5033,G3731,G4119);
  nand GNAME5034(G5034,G3727,G4121);
  nand GNAME5035(G5035,G8955,G4117);
  nand GNAME5036(G5036,G4744,G4115);
  nand GNAME5037(G5037,G4112,G22935);
  nand GNAME5038(G5038,G9374,G4114);
  nand GNAME5039(G5039,G3733,G4119);
  nand GNAME5040(G5040,G3729,G4121);
  nand GNAME5041(G5041,G9015,G4117);
  nand GNAME5042(G5042,G4603,G4115);
  nand GNAME5043(G5043,G4112,G22934);
  nand GNAME5044(G5044,G9388,G4114);
  nand GNAME5045(G5045,G3735,G4119);
  nand GNAME5046(G5046,G3731,G4121);
  nand GNAME5047(G5047,G9018,G4117);
  nand GNAME5048(G5048,G4648,G4115);
  nand GNAME5049(G5049,G4112,G22933);
  nand GNAME5050(G5050,G9396,G4114);
  nand GNAME5051(G5051,G3737,G4119);
  nand GNAME5052(G5052,G3733,G4121);
  nand GNAME5053(G5053,G8993,G4117);
  nand GNAME5054(G5054,G4506,G4115);
  nand GNAME5055(G5055,G4112,G22932);
  nand GNAME5056(G5056,G9392,G4114);
  nand GNAME5057(G5057,G3739,G4119);
  nand GNAME5058(G5058,G3735,G4121);
  nand GNAME5059(G5059,G8954,G4117);
  nand GNAME5060(G5060,G4728,G4115);
  nand GNAME5061(G5061,G4112,G22931);
  nand GNAME5062(G5062,G23018,G4114);
  nand GNAME5063(G5063,G3741,G4119);
  nand GNAME5064(G5064,G3737,G4121);
  nand GNAME5065(G5065,G4170,G4077);
  or GNAME5066(G5066,G5938,G4081);
  nand GNAME5067(G5067,G4171,G4176);
  nand GNAME5068(G5068,G5067,G4083,G5066,G4082,G5065);
  nand GNAME5069(G5069,G4562,G4115);
  nand GNAME5070(G5070,G23033,G4114);
  nand GNAME5071(G5071,G3743,G4119);
  nand GNAME5072(G5072,G3739,G4121);
  nand GNAME5073(G5073,G8991,G4117);
  nand GNAME5074(G5074,G4674,G4115);
  nand GNAME5075(G5075,G4112,G22929);
  nand GNAME5076(G5076,G23023,G4114);
  nand GNAME5077(G5077,G3741,G4121);
  nand GNAME5078(G5078,G4170,G4176);
  nand GNAME5079(G5079,G5078,G4367,G4359);
  nand GNAME5080(G5080,G4080,G5079);
  not GNAME5081(G5081,G4122);
  nand GNAME5082(G5082,G4122,G22928);
  nand GNAME5083(G5083,G4101,G4123);
  nand GNAME5084(G5084,G4122,G22927);
  nand GNAME5085(G5085,G4103,G4123);
  nand GNAME5086(G5086,G4390,G4176);
  nand GNAME5087(G5087,G4083,G4081,G5086);
  nand GNAME5088(G5088,G9042,G4124);
  nand GNAME5089(G5089,G3687,G4125);
  nand GNAME5090(G5090,G4102,G4123);
  nand GNAME5091(G5091,G9045,G4124);
  nand GNAME5092(G5092,G4122,G22925);
  nand GNAME5093(G5093,G3689,G4125);
  nand GNAME5094(G5094,G4094,G4123);
  nand GNAME5095(G5095,G3685,G4126);
  nand GNAME5096(G5096,G9048,G4124);
  nand GNAME5097(G5097,G4122,G22924);
  nand GNAME5098(G5098,G3691,G4125);
  nand GNAME5099(G5099,G4092,G4123);
  nand GNAME5100(G5100,G3687,G4126);
  nand GNAME5101(G5101,G9051,G4124);
  nand GNAME5102(G5102,G4122,G22923);
  nand GNAME5103(G5103,G3693,G4125);
  nand GNAME5104(G5104,G4100,G4123);
  nand GNAME5105(G5105,G3689,G4126);
  nand GNAME5106(G5106,G9054,G4124);
  nand GNAME5107(G5107,G4122,G22922);
  nand GNAME5108(G5108,G3695,G4125);
  nand GNAME5109(G5109,G4096,G4123);
  nand GNAME5110(G5110,G3691,G4126);
  nand GNAME5111(G5111,G9057,G4124);
  nand GNAME5112(G5112,G4122,G22921);
  nand GNAME5113(G5113,G3697,G4125);
  nand GNAME5114(G5114,G4097,G4123);
  nand GNAME5115(G5115,G3693,G4126);
  nand GNAME5116(G5116,G9060,G4124);
  nand GNAME5117(G5117,G4122,G22920);
  nand GNAME5118(G5118,G3699,G4125);
  nand GNAME5119(G5119,G4093,G4123);
  nand GNAME5120(G5120,G3695,G4126);
  nand GNAME5121(G5121,G9063,G4124);
  nand GNAME5122(G5122,G4122,G22919);
  nand GNAME5123(G5123,G3701,G4125);
  nand GNAME5124(G5124,G4099,G4123);
  nand GNAME5125(G5125,G3697,G4126);
  nand GNAME5126(G5126,G9066,G4124);
  nand GNAME5127(G5127,G4122,G22918);
  nand GNAME5128(G5128,G3703,G4125);
  nand GNAME5129(G5129,G4095,G4123);
  nand GNAME5130(G5130,G3699,G4126);
  nand GNAME5131(G5131,G9069,G4124);
  nand GNAME5132(G5132,G4122,G22917);
  nand GNAME5133(G5133,G3705,G4125);
  nand GNAME5134(G5134,G4098,G4123);
  nand GNAME5135(G5135,G3701,G4126);
  nand GNAME5136(G5136,G9075,G4124);
  nand GNAME5137(G5137,G4523,G4123);
  nand GNAME5138(G5138,G4122,G22916);
  nand GNAME5139(G5139,G3707,G4125);
  nand GNAME5140(G5140,G3703,G4126);
  nand GNAME5141(G5141,G9078,G4124);
  nand GNAME5142(G5142,G4736,G4123);
  nand GNAME5143(G5143,G4122,G22915);
  nand GNAME5144(G5144,G3709,G4125);
  nand GNAME5145(G5145,G3705,G4126);
  nand GNAME5146(G5146,G9081,G4124);
  nand GNAME5147(G5147,G4616,G4123);
  nand GNAME5148(G5148,G4122,G22914);
  nand GNAME5149(G5149,G3711,G4125);
  nand GNAME5150(G5150,G3707,G4126);
  nand GNAME5151(G5151,G9084,G4124);
  nand GNAME5152(G5152,G4595,G4123);
  nand GNAME5153(G5153,G4122,G22913);
  nand GNAME5154(G5154,G3713,G4125);
  nand GNAME5155(G5155,G3709,G4126);
  nand GNAME5156(G5156,G9087,G4124);
  nand GNAME5157(G5157,G4758,G4123);
  nand GNAME5158(G5158,G4122,G22912);
  nand GNAME5159(G5159,G3715,G4125);
  nand GNAME5160(G5160,G3711,G4126);
  nand GNAME5161(G5161,G8996,G4124);
  nand GNAME5162(G5162,G4456,G4123);
  nand GNAME5163(G5163,G4122,G22911);
  nand GNAME5164(G5164,G3717,G4125);
  nand GNAME5165(G5165,G3713,G4126);
  nand GNAME5166(G5166,G9091,G4124);
  nand GNAME5167(G5167,G4706,G4123);
  nand GNAME5168(G5168,G4122,G22910);
  nand GNAME5169(G5169,G3719,G4125);
  nand GNAME5170(G5170,G3715,G4126);
  nand GNAME5171(G5171,G9094,G4124);
  nand GNAME5172(G5172,G4576,G4123);
  nand GNAME5173(G5173,G4122,G22909);
  nand GNAME5174(G5174,G3721,G4125);
  nand GNAME5175(G5175,G3717,G4126);
  nand GNAME5176(G5176,G8997,G4124);
  nand GNAME5177(G5177,G4720,G4123);
  nand GNAME5178(G5178,G4122,G22908);
  nand GNAME5179(G5179,G3723,G4125);
  nand GNAME5180(G5180,G3719,G4126);
  nand GNAME5181(G5181,G8953,G4124);
  nand GNAME5182(G5182,G4488,G4123);
  nand GNAME5183(G5183,G4122,G22907);
  nand GNAME5184(G5184,G3725,G4125);
  nand GNAME5185(G5185,G3721,G4126);
  nand GNAME5186(G5186,G9008,G4124);
  nand GNAME5187(G5187,G4661,G4123);
  nand GNAME5188(G5188,G4122,G22906);
  nand GNAME5189(G5189,G3727,G4125);
  nand GNAME5190(G5190,G3723,G4126);
  nand GNAME5191(G5191,G9011,G4124);
  nand GNAME5192(G5192,G4549,G4123);
  nand GNAME5193(G5193,G4122,G22905);
  nand GNAME5194(G5194,G3729,G4125);
  nand GNAME5195(G5195,G3725,G4126);
  nand GNAME5196(G5196,G8992,G4124);
  nand GNAME5197(G5197,G4410,G4123);
  nand GNAME5198(G5198,G4122,G22904);
  nand GNAME5199(G5199,G3731,G4125);
  nand GNAME5200(G5200,G3727,G4126);
  nand GNAME5201(G5201,G8955,G4124);
  nand GNAME5202(G5202,G4744,G4123);
  nand GNAME5203(G5203,G4122,G22903);
  nand GNAME5204(G5204,G3733,G4125);
  nand GNAME5205(G5205,G3729,G4126);
  nand GNAME5206(G5206,G9015,G4124);
  nand GNAME5207(G5207,G4603,G4123);
  nand GNAME5208(G5208,G4122,G22902);
  nand GNAME5209(G5209,G3735,G4125);
  nand GNAME5210(G5210,G3731,G4126);
  nand GNAME5211(G5211,G9018,G4124);
  nand GNAME5212(G5212,G4648,G4123);
  nand GNAME5213(G5213,G4122,G22901);
  nand GNAME5214(G5214,G3737,G4125);
  nand GNAME5215(G5215,G3733,G4126);
  nand GNAME5216(G5216,G8993,G4124);
  nand GNAME5217(G5217,G4506,G4123);
  nand GNAME5218(G5218,G4122,G22900);
  nand GNAME5219(G5219,G3739,G4125);
  nand GNAME5220(G5220,G3735,G4126);
  nand GNAME5221(G5221,G8954,G4124);
  nand GNAME5222(G5222,G4728,G4123);
  nand GNAME5223(G5223,G4122,G22899);
  nand GNAME5224(G5224,G3741,G4125);
  nand GNAME5225(G5225,G3737,G4126);
  nand GNAME5226(G5226,G9072,G4124);
  nand GNAME5227(G5227,G4562,G4123);
  nand GNAME5228(G5228,G4122,G22898);
  nand GNAME5229(G5229,G3743,G4125);
  nand GNAME5230(G5230,G3739,G4126);
  nand GNAME5231(G5231,G8991,G4124);
  nand GNAME5232(G5232,G4674,G4123);
  nand GNAME5233(G5233,G4122,G22897);
  nand GNAME5234(G5234,G3741,G4126);
  nand GNAME5235(G5235,G4375,G6225);
  nand GNAME5236(G5236,G4086,G4411);
  nand GNAME5237(G5237,G5236,G4087);
  nand GNAME5238(G5238,G5235,G4400);
  nand GNAME5239(G5239,G5237,G5238);
  not GNAME5240(G5240,G4127);
  nand GNAME5241(G5241,G4127,G22896);
  nand GNAME5242(G5242,G4101,G4128);
  nand GNAME5243(G5243,G4127,G22895);
  nand GNAME5244(G5244,G4103,G4128);
  nand GNAME5245(G5245,G9042,G4129);
  nand GNAME5246(G5246,G3687,G4130);
  nand GNAME5247(G5247,G4102,G4128);
  nand GNAME5248(G5248,G9045,G4129);
  nand GNAME5249(G5249,G4127,G22893);
  nand GNAME5250(G5250,G3689,G4130);
  nand GNAME5251(G5251,G4094,G4128);
  nand GNAME5252(G5252,G3685,G4131);
  nand GNAME5253(G5253,G9048,G4129);
  nand GNAME5254(G5254,G4127,G22892);
  nand GNAME5255(G5255,G3691,G4130);
  nand GNAME5256(G5256,G4092,G4128);
  nand GNAME5257(G5257,G3687,G4131);
  nand GNAME5258(G5258,G9051,G4129);
  nand GNAME5259(G5259,G4127,G22891);
  nand GNAME5260(G5260,G3693,G4130);
  nand GNAME5261(G5261,G4100,G4128);
  nand GNAME5262(G5262,G3689,G4131);
  nand GNAME5263(G5263,G9054,G4129);
  nand GNAME5264(G5264,G4127,G22890);
  nand GNAME5265(G5265,G3695,G4130);
  nand GNAME5266(G5266,G4096,G4128);
  nand GNAME5267(G5267,G3691,G4131);
  nand GNAME5268(G5268,G9057,G4129);
  nand GNAME5269(G5269,G4127,G22889);
  nand GNAME5270(G5270,G3697,G4130);
  nand GNAME5271(G5271,G4097,G4128);
  nand GNAME5272(G5272,G3693,G4131);
  nand GNAME5273(G5273,G9060,G4129);
  nand GNAME5274(G5274,G4127,G22888);
  nand GNAME5275(G5275,G3699,G4130);
  nand GNAME5276(G5276,G4093,G4128);
  nand GNAME5277(G5277,G3695,G4131);
  nand GNAME5278(G5278,G9063,G4129);
  nand GNAME5279(G5279,G4127,G22887);
  nand GNAME5280(G5280,G3701,G4130);
  nand GNAME5281(G5281,G4099,G4128);
  nand GNAME5282(G5282,G3697,G4131);
  nand GNAME5283(G5283,G9066,G4129);
  nand GNAME5284(G5284,G4127,G22886);
  nand GNAME5285(G5285,G3703,G4130);
  nand GNAME5286(G5286,G4095,G4128);
  nand GNAME5287(G5287,G3699,G4131);
  nand GNAME5288(G5288,G9069,G4129);
  nand GNAME5289(G5289,G4127,G22885);
  nand GNAME5290(G5290,G3705,G4130);
  nand GNAME5291(G5291,G4098,G4128);
  nand GNAME5292(G5292,G3701,G4131);
  nand GNAME5293(G5293,G9075,G4129);
  nand GNAME5294(G5294,G4523,G4128);
  nand GNAME5295(G5295,G4127,G22884);
  nand GNAME5296(G5296,G3707,G4130);
  nand GNAME5297(G5297,G3703,G4131);
  nand GNAME5298(G5298,G9078,G4129);
  nand GNAME5299(G5299,G4736,G4128);
  nand GNAME5300(G5300,G4127,G22883);
  nand GNAME5301(G5301,G3709,G4130);
  nand GNAME5302(G5302,G3705,G4131);
  nand GNAME5303(G5303,G9081,G4129);
  nand GNAME5304(G5304,G4616,G4128);
  nand GNAME5305(G5305,G4127,G22882);
  nand GNAME5306(G5306,G3711,G4130);
  nand GNAME5307(G5307,G3707,G4131);
  nand GNAME5308(G5308,G9084,G4129);
  nand GNAME5309(G5309,G4595,G4128);
  nand GNAME5310(G5310,G4127,G22881);
  nand GNAME5311(G5311,G3713,G4130);
  nand GNAME5312(G5312,G3709,G4131);
  nand GNAME5313(G5313,G9087,G4129);
  nand GNAME5314(G5314,G4758,G4128);
  nand GNAME5315(G5315,G4127,G22880);
  nand GNAME5316(G5316,G3715,G4130);
  nand GNAME5317(G5317,G3711,G4131);
  nand GNAME5318(G5318,G8996,G4129);
  nand GNAME5319(G5319,G4456,G4128);
  nand GNAME5320(G5320,G4127,G22879);
  nand GNAME5321(G5321,G3717,G4130);
  nand GNAME5322(G5322,G3713,G4131);
  nand GNAME5323(G5323,G9091,G4129);
  nand GNAME5324(G5324,G4706,G4128);
  nand GNAME5325(G5325,G4127,G22878);
  nand GNAME5326(G5326,G3719,G4130);
  nand GNAME5327(G5327,G3715,G4131);
  nand GNAME5328(G5328,G9094,G4129);
  nand GNAME5329(G5329,G4576,G4128);
  nand GNAME5330(G5330,G4127,G22877);
  nand GNAME5331(G5331,G3721,G4130);
  nand GNAME5332(G5332,G3717,G4131);
  nand GNAME5333(G5333,G8997,G4129);
  nand GNAME5334(G5334,G4720,G4128);
  nand GNAME5335(G5335,G4127,G22876);
  nand GNAME5336(G5336,G3723,G4130);
  nand GNAME5337(G5337,G3719,G4131);
  nand GNAME5338(G5338,G8953,G4129);
  nand GNAME5339(G5339,G4488,G4128);
  nand GNAME5340(G5340,G4127,G22875);
  nand GNAME5341(G5341,G3725,G4130);
  nand GNAME5342(G5342,G3721,G4131);
  nand GNAME5343(G5343,G9008,G4129);
  nand GNAME5344(G5344,G4661,G4128);
  nand GNAME5345(G5345,G4127,G22874);
  nand GNAME5346(G5346,G3727,G4130);
  nand GNAME5347(G5347,G3723,G4131);
  nand GNAME5348(G5348,G9011,G4129);
  nand GNAME5349(G5349,G4549,G4128);
  nand GNAME5350(G5350,G4127,G22873);
  nand GNAME5351(G5351,G3729,G4130);
  nand GNAME5352(G5352,G3725,G4131);
  nand GNAME5353(G5353,G8992,G4129);
  nand GNAME5354(G5354,G4410,G4128);
  nand GNAME5355(G5355,G4127,G22872);
  nand GNAME5356(G5356,G3731,G4130);
  nand GNAME5357(G5357,G3727,G4131);
  nand GNAME5358(G5358,G8955,G4129);
  nand GNAME5359(G5359,G4744,G4128);
  nand GNAME5360(G5360,G4127,G22871);
  nand GNAME5361(G5361,G3733,G4130);
  nand GNAME5362(G5362,G3729,G4131);
  nand GNAME5363(G5363,G9015,G4129);
  nand GNAME5364(G5364,G4603,G4128);
  nand GNAME5365(G5365,G4127,G22870);
  nand GNAME5366(G5366,G3735,G4130);
  nand GNAME5367(G5367,G3731,G4131);
  nand GNAME5368(G5368,G9018,G4129);
  nand GNAME5369(G5369,G4648,G4128);
  nand GNAME5370(G5370,G4127,G22869);
  nand GNAME5371(G5371,G3737,G4130);
  nand GNAME5372(G5372,G3733,G4131);
  nand GNAME5373(G5373,G8993,G4129);
  nand GNAME5374(G5374,G4506,G4128);
  nand GNAME5375(G5375,G4127,G22868);
  nand GNAME5376(G5376,G3739,G4130);
  nand GNAME5377(G5377,G3735,G4131);
  nand GNAME5378(G5378,G8954,G4129);
  nand GNAME5379(G5379,G4728,G4128);
  nand GNAME5380(G5380,G4127,G22867);
  nand GNAME5381(G5381,G3741,G4130);
  nand GNAME5382(G5382,G3737,G4131);
  nand GNAME5383(G5383,G9072,G4129);
  nand GNAME5384(G5384,G4562,G4128);
  nand GNAME5385(G5385,G4127,G22866);
  nand GNAME5386(G5386,G3743,G4130);
  nand GNAME5387(G5387,G3739,G4131);
  nand GNAME5388(G5388,G8991,G4129);
  nand GNAME5389(G5389,G4674,G4128);
  nand GNAME5390(G5390,G4127,G22865);
  nand GNAME5391(G5391,G3741,G4131);
  not GNAME5392(G5392,G4364);
  nand GNAME5393(G5393,G22832,G4132);
  nand GNAME5394(G5394,G8892,G4133);
  nand GNAME5395(G5395,G3841,G554);
  nand GNAME5396(G5396,G8893,G4133);
  nand GNAME5397(G5397,G22831,G4132);
  nand GNAME5398(G5398,G3841,G555);
  nand GNAME5399(G5399,G22830,G4132);
  nand GNAME5400(G5400,G8861,G4133);
  nand GNAME5401(G5401,G3841,G557);
  nand GNAME5402(G5402,G22829,G4132);
  nand GNAME5403(G5403,G8866,G4133);
  nand GNAME5404(G5404,G3841,G558);
  nand GNAME5405(G5405,G22828,G4132);
  nand GNAME5406(G5406,G8894,G4133);
  nand GNAME5407(G5407,G3841,G559);
  nand GNAME5408(G5408,G22827,G4132);
  nand GNAME5409(G5409,G8860,G4133);
  nand GNAME5410(G5410,G3841,G560);
  nand GNAME5411(G5411,G4132,G22826);
  nand GNAME5412(G5412,G4133,G8895);
  nand GNAME5413(G5413,G3841,G561);
  nand GNAME5414(G5414,G22825,G4132);
  nand GNAME5415(G5415,G8867,G4133);
  nand GNAME5416(G5416,G3841,G562);
  nand GNAME5417(G5417,G22824,G4132);
  nand GNAME5418(G5418,G8896,G4133);
  nand GNAME5419(G5419,G3841,G563);
  nand GNAME5420(G5420,G22823,G4132);
  nand GNAME5421(G5421,G8859,G4133);
  nand GNAME5422(G5422,G3841,G564);
  nand GNAME5423(G5423,G22822,G4132);
  nand GNAME5424(G5424,G8897,G4133);
  nand GNAME5425(G5425,G3841,G565);
  nand GNAME5426(G5426,G22821,G4132);
  nand GNAME5427(G5427,G8868,G4133);
  nand GNAME5428(G5428,G3841,G566);
  nand GNAME5429(G5429,G22820,G4132);
  nand GNAME5430(G5430,G8899,G4133);
  nand GNAME5431(G5431,G3841,G568);
  nand GNAME5432(G5432,G22819,G4132);
  nand GNAME5433(G5433,G8858,G4133);
  nand GNAME5434(G5434,G3841,G569);
  nand GNAME5435(G5435,G22818,G4132);
  nand GNAME5436(G5436,G8900,G4133);
  nand GNAME5437(G5437,G3841,G570);
  nand GNAME5438(G5438,G22817,G4132);
  nand GNAME5439(G5439,G8869,G4133);
  nand GNAME5440(G5440,G3841,G571);
  nand GNAME5441(G5441,G22816,G4132);
  nand GNAME5442(G5442,G8901,G4133);
  nand GNAME5443(G5443,G3841,G572);
  nand GNAME5444(G5444,G22815,G4132);
  nand GNAME5445(G5445,G8857,G4133);
  nand GNAME5446(G5446,G3841,G573);
  nand GNAME5447(G5447,G22814,G4132);
  nand GNAME5448(G5448,G8902,G4133);
  nand GNAME5449(G5449,G3841,G574);
  nand GNAME5450(G5450,G22813,G4132);
  nand GNAME5451(G5451,G8870,G4133);
  nand GNAME5452(G5452,G3841,G575);
  nand GNAME5453(G5453,G22812,G4132);
  nand GNAME5454(G5454,G8903,G4133);
  nand GNAME5455(G5455,G3841,G576);
  nand GNAME5456(G5456,G22811,G4132);
  nand GNAME5457(G5457,G8856,G4133);
  nand GNAME5458(G5458,G3841,G577);
  nand GNAME5459(G5459,G22810,G4132);
  nand GNAME5460(G5460,G8888,G4133);
  nand GNAME5461(G5461,G3841,G547);
  nand GNAME5462(G5462,G22809,G4132);
  nand GNAME5463(G5463,G8864,G4133);
  nand GNAME5464(G5464,G3841,G548);
  nand GNAME5465(G5465,G22808,G4132);
  nand GNAME5466(G5466,G8889,G4133);
  nand GNAME5467(G5467,G3841,G549);
  nand GNAME5468(G5468,G22807,G4132);
  nand GNAME5469(G5469,G8863,G4133);
  nand GNAME5470(G5470,G3841,G550);
  nand GNAME5471(G5471,G22806,G4132);
  nand GNAME5472(G5472,G8890,G4133);
  nand GNAME5473(G5473,G3841,G551);
  nand GNAME5474(G5474,G22805,G4132);
  nand GNAME5475(G5475,G8865,G4133);
  nand GNAME5476(G5476,G3841,G552);
  nand GNAME5477(G5477,G22804,G4132);
  nand GNAME5478(G5478,G8891,G4133);
  nand GNAME5479(G5479,G3841,G553);
  nand GNAME5480(G5480,G22803,G4132);
  nand GNAME5481(G5481,G8862,G4133);
  nand GNAME5482(G5482,G3841,G556);
  nand GNAME5483(G5483,G22802,G4132);
  nand GNAME5484(G5484,G8886,G4133);
  nand GNAME5485(G5485,G3841,G567);
  nand GNAME5486(G5486,G22801,G4132);
  nand GNAME5487(G5487,G22801,G4133);
  nand GNAME5488(G5488,G3841,G578);
  or GNAME5489(G5489,G4059,G4368,G4079);
  not GNAME5490(G5490,G4135);
  nand GNAME5491(G5491,G5891,G5490);
  nand GNAME5492(G5492,G5891,G4171,G4176);
  nand GNAME5493(G5493,G5492,G4359);
  nand GNAME5494(G5494,G5971,G5974,G4077,G5941);
  nand GNAME5495(G5495,G5493,G4075);
  nand GNAME5496(G5496,G5494,G5495);
  nand GNAME5497(G5497,G5971,G5974);
  nand GNAME5498(G5498,G4053,G5497,G4077,G5941);
  nand GNAME5499(G5499,G5493,G4053,G4399);
  or GNAME5500(G5500,G4140,G4134);
  nand GNAME5501(G5501,G5500,G4190);
  nand GNAME5502(G5502,G3725,G5491);
  nand GNAME5503(G5503,G22906,G4136);
  nand GNAME5504(G5504,G22938,G4137);
  nand GNAME5505(G5505,G5500,G4183);
  nand GNAME5506(G5506,G3727,G5491);
  nand GNAME5507(G5507,G22905,G4136);
  nand GNAME5508(G5508,G22937,G4137);
  nand GNAME5509(G5509,G5500,G4178);
  nand GNAME5510(G5510,G3729,G5491);
  nand GNAME5511(G5511,G22904,G4136);
  nand GNAME5512(G5512,G22936,G4137);
  nand GNAME5513(G5513,G5500,G4196);
  nand GNAME5514(G5514,G3731,G5491);
  nand GNAME5515(G5515,G22903,G4136);
  nand GNAME5516(G5516,G22935,G4137);
  nand GNAME5517(G5517,G5500,G4187);
  nand GNAME5518(G5518,G3733,G5491);
  nand GNAME5519(G5519,G22902,G4136);
  nand GNAME5520(G5520,G22934,G4137);
  nand GNAME5521(G5521,G5500,G4189);
  nand GNAME5522(G5522,G3735,G5491);
  nand GNAME5523(G5523,G22901,G4136);
  nand GNAME5524(G5524,G22933,G4137);
  nand GNAME5525(G5525,G22916,G4136);
  nand GNAME5526(G5526,G22948,G4137);
  nand GNAME5527(G5527,G3687,G4138);
  nand GNAME5528(G5528,G3685,G4139);
  nand GNAME5529(G5529,G4134,G4102);
  nand GNAME5530(G5530,G4094,G4140);
  nand GNAME5531(G5531,G3681,G4147);
  nand GNAME5532(G5532,G3683,G4147);
  nand GNAME5533(G5533,G5500,G4181);
  nand GNAME5534(G5534,G3737,G5491);
  nand GNAME5535(G5535,G22900,G4136);
  nand GNAME5536(G5536,G22932,G4137);
  nand GNAME5537(G5537,G3685,G4147);
  nand GNAME5538(G5538,G5500,G4094);
  nand GNAME5539(G5539,G3687,G5491);
  nand GNAME5540(G5540,G5500,G4092);
  nand GNAME5541(G5541,G3689,G5491);
  nand GNAME5542(G5542,G5500,G4100);
  nand GNAME5543(G5543,G3691,G5491);
  nand GNAME5544(G5544,G5500,G4096);
  nand GNAME5545(G5545,G3693,G5491);
  nand GNAME5546(G5546,G5500,G4097);
  nand GNAME5547(G5547,G3695,G5491);
  nand GNAME5548(G5548,G5500,G4093);
  nand GNAME5549(G5549,G3697,G5491);
  nand GNAME5550(G5550,G5500,G4099);
  nand GNAME5551(G5551,G3699,G5491);
  nand GNAME5552(G5552,G5500,G4095);
  nand GNAME5553(G5553,G3701,G5491);
  nand GNAME5554(G5554,G5500,G4098);
  nand GNAME5555(G5555,G3703,G5491);
  nand GNAME5556(G5556,G5500,G4194);
  nand GNAME5557(G5557,G3739,G5491);
  nand GNAME5558(G5558,G22899,G4136);
  nand GNAME5559(G5559,G22931,G4137);
  nand GNAME5560(G5560,G5500,G4182);
  nand GNAME5561(G5561,G3705,G5491);
  nand GNAME5562(G5562,G5500,G4195);
  nand GNAME5563(G5563,G3707,G5491);
  nand GNAME5564(G5564,G22915,G4136);
  nand GNAME5565(G5565,G22947,G4137);
  nand GNAME5566(G5566,G5500,G4188);
  nand GNAME5567(G5567,G3709,G5491);
  nand GNAME5568(G5568,G22914,G4136);
  nand GNAME5569(G5569,G22946,G4137);
  nand GNAME5570(G5570,G5500,G4186);
  nand GNAME5571(G5571,G3711,G5491);
  nand GNAME5572(G5572,G22913,G4136);
  nand GNAME5573(G5573,G22945,G4137);
  nand GNAME5574(G5574,G5500,G4197);
  nand GNAME5575(G5575,G3713,G5491);
  nand GNAME5576(G5576,G22912,G4136);
  nand GNAME5577(G5577,G22944,G4137);
  nand GNAME5578(G5578,G5500,G4179);
  nand GNAME5579(G5579,G3715,G5491);
  nand GNAME5580(G5580,G22911,G4136);
  nand GNAME5581(G5581,G22943,G4137);
  nand GNAME5582(G5582,G5500,G4192);
  nand GNAME5583(G5583,G3717,G5491);
  nand GNAME5584(G5584,G22910,G4136);
  nand GNAME5585(G5585,G22942,G4137);
  nand GNAME5586(G5586,G5500,G4185);
  nand GNAME5587(G5587,G3719,G5491);
  nand GNAME5588(G5588,G22909,G4136);
  nand GNAME5589(G5589,G22941,G4137);
  nand GNAME5590(G5590,G5500,G4193);
  nand GNAME5591(G5591,G3721,G5491);
  nand GNAME5592(G5592,G22908,G4136);
  nand GNAME5593(G5593,G22940,G4137);
  nand GNAME5594(G5594,G5500,G4180);
  nand GNAME5595(G5595,G3723,G5491);
  nand GNAME5596(G5596,G22907,G4136);
  nand GNAME5597(G5597,G22939,G4137);
  nand GNAME5598(G5598,G5500,G4184);
  nand GNAME5599(G5599,G3741,G5491);
  nand GNAME5600(G5600,G22898,G4136);
  nand GNAME5601(G5601,G22930,G4137);
  nand GNAME5602(G5602,G5500,G4191);
  nand GNAME5603(G5603,G3743,G5491);
  nand GNAME5604(G5604,G22897,G4136);
  nand GNAME5605(G5605,G22929,G4137);
  or GNAME5606(G5606,G4136,G4137);
  nand GNAME5607(G5607,G3725,G5500);
  nand GNAME5608(G5608,G4135,G4190);
  nand GNAME5609(G5609,G5606,G4151);
  nand GNAME5610(G5610,G3727,G5500);
  nand GNAME5611(G5611,G4135,G4183);
  nand GNAME5612(G5612,G5606,G4152);
  nand GNAME5613(G5613,G3729,G5500);
  nand GNAME5614(G5614,G4135,G4178);
  nand GNAME5615(G5615,G5606,G4153);
  nand GNAME5616(G5616,G3731,G5500);
  nand GNAME5617(G5617,G4135,G4196);
  nand GNAME5618(G5618,G5606,G4154);
  nand GNAME5619(G5619,G3733,G5500);
  nand GNAME5620(G5620,G4135,G4187);
  nand GNAME5621(G5621,G5606,G4155);
  nand GNAME5622(G5622,G3735,G5500);
  nand GNAME5623(G5623,G4135,G4189);
  nand GNAME5624(G5624,G5606,G4156);
  nand GNAME5625(G5625,G5606,G4175);
  nand GNAME5626(G5626,G4102,G4139);
  nand GNAME5627(G5627,G4094,G4138);
  nand GNAME5628(G5628,G3685,G4134);
  nand GNAME5629(G5629,G3687,G4140);
  nand GNAME5630(G5630,G3737,G5500);
  nand GNAME5631(G5631,G4135,G4181);
  nand GNAME5632(G5632,G5606,G4157);
  nand GNAME5633(G5633,G3687,G5500);
  nand GNAME5634(G5634,G4135,G4094);
  nand GNAME5635(G5635,G3689,G5500);
  nand GNAME5636(G5636,G4135,G4092);
  nand GNAME5637(G5637,G3691,G5500);
  nand GNAME5638(G5638,G4135,G4100);
  nand GNAME5639(G5639,G3693,G5500);
  nand GNAME5640(G5640,G4135,G4096);
  nand GNAME5641(G5641,G3695,G5500);
  nand GNAME5642(G5642,G4135,G4097);
  nand GNAME5643(G5643,G3697,G5500);
  nand GNAME5644(G5644,G4135,G4093);
  nand GNAME5645(G5645,G3699,G5500);
  nand GNAME5646(G5646,G4135,G4099);
  nand GNAME5647(G5647,G3701,G5500);
  nand GNAME5648(G5648,G4135,G4095);
  nand GNAME5649(G5649,G3703,G5500);
  nand GNAME5650(G5650,G4135,G4098);
  nand GNAME5651(G5651,G3739,G5500);
  nand GNAME5652(G5652,G4135,G4194);
  nand GNAME5653(G5653,G5606,G4158);
  nand GNAME5654(G5654,G3705,G5500);
  nand GNAME5655(G5655,G4135,G4182);
  nand GNAME5656(G5656,G3707,G5500);
  nand GNAME5657(G5657,G4135,G4195);
  nand GNAME5658(G5658,G5606,G4160);
  nand GNAME5659(G5659,G3709,G5500);
  nand GNAME5660(G5660,G4135,G4188);
  nand GNAME5661(G5661,G5606,G4161);
  nand GNAME5662(G5662,G3711,G5500);
  nand GNAME5663(G5663,G4135,G4186);
  nand GNAME5664(G5664,G5606,G4162);
  nand GNAME5665(G5665,G3713,G5500);
  nand GNAME5666(G5666,G4135,G4197);
  nand GNAME5667(G5667,G5606,G4163);
  nand GNAME5668(G5668,G3715,G5500);
  nand GNAME5669(G5669,G4135,G4179);
  nand GNAME5670(G5670,G5606,G4164);
  nand GNAME5671(G5671,G3717,G5500);
  nand GNAME5672(G5672,G4135,G4192);
  nand GNAME5673(G5673,G5606,G4165);
  nand GNAME5674(G5674,G3719,G5500);
  nand GNAME5675(G5675,G4135,G4185);
  nand GNAME5676(G5676,G5606,G4166);
  nand GNAME5677(G5677,G3721,G5500);
  nand GNAME5678(G5678,G4135,G4193);
  nand GNAME5679(G5679,G5606,G4167);
  nand GNAME5680(G5680,G3723,G5500);
  nand GNAME5681(G5681,G4135,G4180);
  nand GNAME5682(G5682,G5606,G4168);
  nand GNAME5683(G5683,G3741,G5500);
  nand GNAME5684(G5684,G4135,G4184);
  nand GNAME5685(G5685,G5606,G4159);
  nand GNAME5686(G5686,G3743,G5500);
  nand GNAME5687(G5687,G4135,G4191);
  nand GNAME5688(G5688,G5606,G4169);
  nand GNAME5689(G5689,G4171,G5962);
  nand GNAME5690(G5690,G4369,G4144);
  nand GNAME5691(G5691,G4147,G4061);
  not GNAME5692(G5692,G4143);
  nand GNAME5693(G5693,G5692,G4051,G5065);
  nand GNAME5694(G5694,G3725,G5693);
  nand GNAME5695(G5695,G5690,G4190);
  nand GNAME5696(G5696,G3727,G5891);
  nand GNAME5697(G5697,G3727,G5693);
  nand GNAME5698(G5698,G5690,G4183);
  nand GNAME5699(G5699,G3729,G5891);
  nand GNAME5700(G5700,G3729,G5693);
  nand GNAME5701(G5701,G5690,G4178);
  nand GNAME5702(G5702,G3731,G5891);
  nand GNAME5703(G5703,G3731,G5693);
  nand GNAME5704(G5704,G5690,G4196);
  nand GNAME5705(G5705,G3733,G5891);
  nand GNAME5706(G5706,G3733,G5693);
  nand GNAME5707(G5707,G5690,G4187);
  nand GNAME5708(G5708,G3735,G5891);
  nand GNAME5709(G5709,G3735,G5693);
  nand GNAME5710(G5710,G5690,G4189);
  nand GNAME5711(G5711,G3737,G5891);
  nand GNAME5712(G5712,G3681,G5693);
  nand GNAME5713(G5713,G5690,G4101);
  nand GNAME5714(G5714,G3683,G5693);
  nand GNAME5715(G5715,G5690,G4103);
  nand GNAME5716(G5716,G3737,G5693);
  nand GNAME5717(G5717,G5690,G4181);
  nand GNAME5718(G5718,G3739,G5891);
  nand GNAME5719(G5719,G3685,G5693);
  nand GNAME5720(G5720,G5690,G4102);
  nand GNAME5721(G5721,G3687,G5891);
  nand GNAME5722(G5722,G3687,G5693);
  nand GNAME5723(G5723,G5690,G4094);
  nand GNAME5724(G5724,G3689,G5891);
  nand GNAME5725(G5725,G3689,G5693);
  nand GNAME5726(G5726,G5690,G4092);
  nand GNAME5727(G5727,G3691,G5891);
  nand GNAME5728(G5728,G3691,G5693);
  nand GNAME5729(G5729,G5690,G4100);
  nand GNAME5730(G5730,G3693,G5891);
  nand GNAME5731(G5731,G3693,G5693);
  nand GNAME5732(G5732,G5690,G4096);
  nand GNAME5733(G5733,G3695,G5891);
  nand GNAME5734(G5734,G3695,G5693);
  nand GNAME5735(G5735,G5690,G4097);
  nand GNAME5736(G5736,G3697,G5891);
  nand GNAME5737(G5737,G3697,G5693);
  nand GNAME5738(G5738,G5690,G4093);
  nand GNAME5739(G5739,G3699,G5891);
  nand GNAME5740(G5740,G3699,G5693);
  nand GNAME5741(G5741,G5690,G4099);
  nand GNAME5742(G5742,G3701,G5891);
  nand GNAME5743(G5743,G3701,G5693);
  nand GNAME5744(G5744,G5690,G4095);
  nand GNAME5745(G5745,G3703,G5891);
  nand GNAME5746(G5746,G3703,G5693);
  nand GNAME5747(G5747,G5690,G4098);
  nand GNAME5748(G5748,G3705,G5891);
  nand GNAME5749(G5749,G3739,G5693);
  nand GNAME5750(G5750,G5690,G4194);
  nand GNAME5751(G5751,G3741,G5891);
  nand GNAME5752(G5752,G3705,G5693);
  nand GNAME5753(G5753,G5690,G4182);
  nand GNAME5754(G5754,G3707,G5891);
  nand GNAME5755(G5755,G3707,G5693);
  nand GNAME5756(G5756,G5690,G4195);
  nand GNAME5757(G5757,G3709,G5891);
  nand GNAME5758(G5758,G3709,G5693);
  nand GNAME5759(G5759,G5690,G4188);
  nand GNAME5760(G5760,G3711,G5891);
  nand GNAME5761(G5761,G3711,G5693);
  nand GNAME5762(G5762,G5690,G4186);
  nand GNAME5763(G5763,G3713,G5891);
  nand GNAME5764(G5764,G3713,G5693);
  nand GNAME5765(G5765,G5690,G4197);
  nand GNAME5766(G5766,G3715,G5891);
  nand GNAME5767(G5767,G3715,G5693);
  nand GNAME5768(G5768,G5690,G4179);
  nand GNAME5769(G5769,G3717,G5891);
  nand GNAME5770(G5770,G3717,G5693);
  nand GNAME5771(G5771,G5690,G4192);
  nand GNAME5772(G5772,G3719,G5891);
  nand GNAME5773(G5773,G3719,G5693);
  nand GNAME5774(G5774,G5690,G4185);
  nand GNAME5775(G5775,G3721,G5891);
  nand GNAME5776(G5776,G3721,G5693);
  nand GNAME5777(G5777,G5690,G4193);
  nand GNAME5778(G5778,G3723,G5891);
  nand GNAME5779(G5779,G3723,G5693);
  nand GNAME5780(G5780,G5690,G4180);
  nand GNAME5781(G5781,G3725,G5891);
  nand GNAME5782(G5782,G3741,G5693);
  nand GNAME5783(G5783,G5690,G4184);
  nand GNAME5784(G5784,G3743,G5891);
  nand GNAME5785(G5785,G3743,G5693);
  nand GNAME5786(G5786,G5690,G4191);
  or GNAME5787(G5787,G546,G4369);
  nand GNAME5788(G5788,G5787,G4144);
  nand GNAME5789(G5789,G3725,G4145);
  nand GNAME5790(G5790,G3725,G5788);
  nand GNAME5791(G5791,G4143,G4190);
  nand GNAME5792(G5792,G4145,G3727);
  nand GNAME5793(G5793,G3727,G5788);
  nand GNAME5794(G5794,G4143,G4183);
  nand GNAME5795(G5795,G4145,G3729);
  nand GNAME5796(G5796,G3729,G5788);
  nand GNAME5797(G5797,G4143,G4178);
  nand GNAME5798(G5798,G4145,G3731);
  nand GNAME5799(G5799,G3731,G5788);
  nand GNAME5800(G5800,G4143,G4196);
  nand GNAME5801(G5801,G4145,G3733);
  nand GNAME5802(G5802,G3733,G5788);
  nand GNAME5803(G5803,G4143,G4187);
  nand GNAME5804(G5804,G4145,G3735);
  nand GNAME5805(G5805,G3735,G5788);
  nand GNAME5806(G5806,G4143,G4189);
  nand GNAME5807(G5807,G4145,G9369);
  nand GNAME5808(G5808,G3681,G5788);
  nand GNAME5809(G5809,G4143,G4101);
  nand GNAME5810(G5810,G4145,G9368);
  nand GNAME5811(G5811,G3683,G5788);
  nand GNAME5812(G5812,G4143,G4103);
  nand GNAME5813(G5813,G4145,G3737);
  nand GNAME5814(G5814,G3737,G5788);
  nand GNAME5815(G5815,G4143,G4181);
  nand GNAME5816(G5816,G4145,G3685);
  nand GNAME5817(G5817,G3685,G5788);
  nand GNAME5818(G5818,G4143,G4102);
  nand GNAME5819(G5819,G4145,G3687);
  nand GNAME5820(G5820,G3687,G5788);
  nand GNAME5821(G5821,G4143,G4094);
  nand GNAME5822(G5822,G4145,G3689);
  nand GNAME5823(G5823,G3689,G5788);
  nand GNAME5824(G5824,G4143,G4092);
  nand GNAME5825(G5825,G4145,G3691);
  nand GNAME5826(G5826,G3691,G5788);
  nand GNAME5827(G5827,G4143,G4100);
  nand GNAME5828(G5828,G4145,G3693);
  nand GNAME5829(G5829,G3693,G5788);
  nand GNAME5830(G5830,G4143,G4096);
  nand GNAME5831(G5831,G4145,G3695);
  nand GNAME5832(G5832,G3695,G5788);
  nand GNAME5833(G5833,G4143,G4097);
  nand GNAME5834(G5834,G4145,G3697);
  nand GNAME5835(G5835,G3697,G5788);
  nand GNAME5836(G5836,G4143,G4093);
  nand GNAME5837(G5837,G4145,G3699);
  nand GNAME5838(G5838,G3699,G5788);
  nand GNAME5839(G5839,G4143,G4099);
  nand GNAME5840(G5840,G4145,G3701);
  nand GNAME5841(G5841,G3701,G5788);
  nand GNAME5842(G5842,G4143,G4095);
  nand GNAME5843(G5843,G4145,G3703);
  nand GNAME5844(G5844,G3703,G5788);
  nand GNAME5845(G5845,G4143,G4098);
  nand GNAME5846(G5846,G4145,G3739);
  nand GNAME5847(G5847,G3739,G5788);
  nand GNAME5848(G5848,G4143,G4194);
  nand GNAME5849(G5849,G4145,G3705);
  nand GNAME5850(G5850,G3705,G5788);
  nand GNAME5851(G5851,G4143,G4182);
  nand GNAME5852(G5852,G4145,G3707);
  nand GNAME5853(G5853,G3707,G5788);
  nand GNAME5854(G5854,G4143,G4195);
  nand GNAME5855(G5855,G4145,G3709);
  nand GNAME5856(G5856,G3709,G5788);
  nand GNAME5857(G5857,G4143,G4188);
  nand GNAME5858(G5858,G4145,G3711);
  nand GNAME5859(G5859,G3711,G5788);
  nand GNAME5860(G5860,G4143,G4186);
  nand GNAME5861(G5861,G4145,G3713);
  nand GNAME5862(G5862,G3713,G5788);
  nand GNAME5863(G5863,G4143,G4197);
  nand GNAME5864(G5864,G4145,G3715);
  nand GNAME5865(G5865,G3715,G5788);
  nand GNAME5866(G5866,G4143,G4179);
  nand GNAME5867(G5867,G4145,G3717);
  nand GNAME5868(G5868,G3717,G5788);
  nand GNAME5869(G5869,G4143,G4192);
  nand GNAME5870(G5870,G4145,G3719);
  nand GNAME5871(G5871,G3719,G5788);
  nand GNAME5872(G5872,G4143,G4185);
  nand GNAME5873(G5873,G4145,G3721);
  nand GNAME5874(G5874,G3721,G5788);
  nand GNAME5875(G5875,G4143,G4193);
  nand GNAME5876(G5876,G4145,G3723);
  nand GNAME5877(G5877,G3723,G5788);
  nand GNAME5878(G5878,G4143,G4180);
  nand GNAME5879(G5879,G4145,G3741);
  nand GNAME5880(G5880,G3741,G5788);
  nand GNAME5881(G5881,G4143,G4184);
  nand GNAME5882(G5882,G4145,G3743);
  nand GNAME5883(G5883,G3743,G5788);
  nand GNAME5884(G5884,G4143,G4191);
  nand GNAME5885(G5885,G4886,G5974);
  nand GNAME5886(G5886,G4884,G4174);
  nand GNAME5887(G5887,G4064,G5080,G4173);
  nand GNAME5888(G5888,G4064,G4886,G5971);
  nand GNAME5889(G5889,G4052,G22824);
  nand GNAME5890(G5890,G22832,G8896);
  not GNAME5891(G5891,G4147);
  or GNAME5892(G5892,G8895,G4052);
  or GNAME5893(G5893,G22826,G22832);
  nand GNAME5894(G5894,G4052,G22827);
  nand GNAME5895(G5895,G8860,G22832);
  nand GNAME5896(G5896,G4052,G22825);
  nand GNAME5897(G5897,G22832,G8867);
  nand GNAME5898(G5898,G4052,G22810);
  nand GNAME5899(G5899,G22832,G8888);
  nand GNAME5900(G5900,G4052,G22809);
  nand GNAME5901(G5901,G22832,G8864);
  nand GNAME5902(G5902,G4052,G22808);
  nand GNAME5903(G5903,G22832,G8889);
  nand GNAME5904(G5904,G4052,G22807);
  nand GNAME5905(G5905,G22832,G8863);
  nand GNAME5906(G5906,G4052,G22806);
  nand GNAME5907(G5907,G22832,G8890);
  nand GNAME5908(G5908,G4052,G22805);
  nand GNAME5909(G5909,G22832,G8865);
  nand GNAME5910(G5910,G4052,G22804);
  nand GNAME5911(G5911,G22832,G8891);
  nand GNAME5912(G5912,G4052,G22803);
  nand GNAME5913(G5913,G22832,G8862);
  nand GNAME5914(G5914,G4052,G22802);
  nand GNAME5915(G5915,G22832,G8886);
  nand GNAME5916(G5916,G4052,G22819);
  nand GNAME5917(G5917,G22832,G8858);
  nand GNAME5918(G5918,G4052,G22818);
  nand GNAME5919(G5919,G22832,G8900);
  nand GNAME5920(G5920,G4052,G22817);
  nand GNAME5921(G5921,G22832,G8869);
  nand GNAME5922(G5922,G4052,G22816);
  nand GNAME5923(G5923,G22832,G8901);
  nand GNAME5924(G5924,G4052,G22815);
  nand GNAME5925(G5925,G22832,G8857);
  nand GNAME5926(G5926,G4052,G22814);
  nand GNAME5927(G5927,G22832,G8902);
  nand GNAME5928(G5928,G4052,G22813);
  nand GNAME5929(G5929,G22832,G8870);
  nand GNAME5930(G5930,G4052,G22812);
  nand GNAME5931(G5931,G22832,G8903);
  nand GNAME5932(G5932,G4052,G22811);
  nand GNAME5933(G5933,G22832,G8856);
  nand GNAME5934(G5934,G4052,G22801);
  nand GNAME5935(G5935,G22832,G22801);
  nand GNAME5936(G5936,G4052,G22823);
  nand GNAME5937(G5937,G22832,G8859);
  not GNAME5938(G5938,G4170);
  nand GNAME5939(G5939,G4052,G22822);
  nand GNAME5940(G5940,G22832,G8897);
  not GNAME5941(G5941,G4171);
  nand GNAME5942(G5942,G4052,G22828);
  nand GNAME5943(G5943,G22832,G8894);
  not GNAME5944(G5944,G4172);
  or GNAME5945(G5945,G22832,G22831,G4070);
  nand GNAME5946(G5946,G22832,G4071,G8861);
  nand GNAME5947(G5947,G5945,G5946);
  nand GNAME5948(G5948,G4052,G4070,G22831);
  nand GNAME5949(G5949,G22832,G4069,G8893);
  nand GNAME5950(G5950,G5948,G5949);
  nand GNAME5951(G5951,G4052,G22830,G22831);
  nand GNAME5952(G5952,G22832,G8861,G8893);
  nand GNAME5953(G5953,G5951,G5952);
  or GNAME5954(G5954,G22832,G22830,G22831);
  nand GNAME5955(G5955,G22832,G4069,G4071);
  nand GNAME5956(G5956,G5954,G5955);
  nand GNAME5957(G5957,G4052,G22820);
  nand GNAME5958(G5958,G22832,G8899);
  not GNAME5959(G5959,G4175);
  nand GNAME5960(G5960,G4052,G22821);
  nand GNAME5961(G5961,G22832,G8868);
  not GNAME5962(G5962,G4176);
  nand GNAME5963(G5963,G4056,G4065);
  or GNAME5964(G5964,G4056,G22832,G22829);
  nand GNAME5965(G5965,G4055,G4066);
  or GNAME5966(G5966,G4055,G8866,G4052);
  nand GNAME5967(G5967,G6336,G4149);
  or GNAME5968(G5968,G6336,G4149,G4150);
  nand GNAME5969(G5969,G4393,G22833);
  nand GNAME5970(G5970,G4063,G4397);
  not GNAME5971(G5971,G4173);
  nand GNAME5972(G5972,G4393,G22834);
  nand GNAME5973(G5973,G4063,G4398);
  not GNAME5974(G5974,G4174);
  or GNAME5975(G5975,G22832,G22828,G22829);
  or GNAME5976(G5976,G4052,G8866,G8894);
  not GNAME5977(G5977,G4177);
  nand GNAME5978(G5978,G4370,G549);
  nand GNAME5979(G5979,G4153,G4356);
  not GNAME5980(G5980,G4178);
  nand GNAME5981(G5981,G4370,G573);
  nand GNAME5982(G5982,G4164,G4356);
  not GNAME5983(G5983,G4179);
  nand GNAME5984(G5984,G4370,G577);
  nand GNAME5985(G5985,G4168,G4356);
  not GNAME5986(G5986,G4180);
  nand GNAME5987(G5987,G4370,G553);
  nand GNAME5988(G5988,G4157,G4356);
  not GNAME5989(G5989,G4181);
  nand GNAME5990(G5990,G4370,G568);
  nand GNAME5991(G5991,G4175,G4356);
  not GNAME5992(G5992,G4182);
  nand GNAME5993(G5993,G4370,G548);
  nand GNAME5994(G5994,G4152,G4356);
  not GNAME5995(G5995,G4183);
  nand GNAME5996(G5996,G4370,G567);
  nand GNAME5997(G5997,G4159,G4356);
  not GNAME5998(G5998,G4184);
  nand GNAME5999(G5999,G4370,G575);
  nand GNAME6000(G6000,G4166,G4356);
  not GNAME6001(G6001,G4185);
  nand GNAME6002(G6002,G4370,G571);
  nand GNAME6003(G6003,G4162,G4356);
  not GNAME6004(G6004,G4186);
  nand GNAME6005(G6005,G4370,G551);
  nand GNAME6006(G6006,G4155,G4356);
  not GNAME6007(G6007,G4187);
  nand GNAME6008(G6008,G4370,G570);
  nand GNAME6009(G6009,G4161,G4356);
  not GNAME6010(G6010,G4188);
  nand GNAME6011(G6011,G4370,G552);
  nand GNAME6012(G6012,G4156,G4356);
  not GNAME6013(G6013,G4189);
  nand GNAME6014(G6014,G4370,G547);
  nand GNAME6015(G6015,G4151,G4356);
  not GNAME6016(G6016,G4190);
  nand GNAME6017(G6017,G4370,G578);
  nand GNAME6018(G6018,G4169,G4356);
  not GNAME6019(G6019,G4191);
  nand GNAME6020(G6020,G4370,G574);
  nand GNAME6021(G6021,G4165,G4356);
  not GNAME6022(G6022,G4192);
  nand GNAME6023(G6023,G4370,G576);
  nand GNAME6024(G6024,G4167,G4356);
  not GNAME6025(G6025,G4193);
  nand GNAME6026(G6026,G4370,G556);
  nand GNAME6027(G6027,G4158,G4356);
  not GNAME6028(G6028,G4194);
  nand GNAME6029(G6029,G4370,G569);
  nand GNAME6030(G6030,G4160,G4356);
  not GNAME6031(G6031,G4195);
  nand GNAME6032(G6032,G4370,G550);
  nand GNAME6033(G6033,G4154,G4356);
  not GNAME6034(G6034,G4196);
  nand GNAME6035(G6035,G4370,G572);
  nand GNAME6036(G6036,G4163,G4356);
  not GNAME6037(G6037,G4197);
  nand GNAME6038(G6038,G4357,G4765,G23013);
  or GNAME6039(G6039,G4104,G4357);
  nand GNAME6040(G6040,G4486,G6016);
  nand GNAME6041(G6041,G3725,G4190);
  nand GNAME6042(G6042,G6040,G6041);
  nand GNAME6043(G6043,G4659,G5986);
  nand GNAME6044(G6044,G3723,G4180);
  nand GNAME6045(G6045,G6043,G6044);
  nand GNAME6046(G6046,G4641,G6007);
  nand GNAME6047(G6047,G3733,G4187);
  nand GNAME6048(G6048,G6046,G6047);
  nand GNAME6049(G6049,G4547,G5980);
  nand GNAME6050(G6050,G3729,G4178);
  nand GNAME6051(G6051,G6049,G6050);
  nand GNAME6052(G6052,G4389,G6034);
  nand GNAME6053(G6053,G3731,G4196);
  nand GNAME6054(G6054,G6052,G6053);
  nand GNAME6055(G6055,G4504,G6028);
  nand GNAME6056(G6056,G3739,G4194);
  nand GNAME6057(G6057,G6055,G6056);
  nand GNAME6058(G6058,G4499,G6013);
  nand GNAME6059(G6059,G3735,G4189);
  nand GNAME6060(G6060,G6058,G6059);
  nand GNAME6061(G6061,G4672,G5998);
  nand GNAME6062(G6062,G3741,G4184);
  nand GNAME6063(G6063,G6061,G6062);
  nand GNAME6064(G6064,G4384,G5995);
  nand GNAME6065(G6065,G3727,G4183);
  nand GNAME6066(G6066,G6064,G6065);
  nand GNAME6067(G6067,G4646,G5989);
  nand GNAME6068(G6068,G3737,G4181);
  nand GNAME6069(G6069,G6067,G6068);
  nand GNAME6070(G6070,G4521,G6031);
  nand GNAME6071(G6071,G3707,G4195);
  nand GNAME6072(G6072,G6070,G6071);
  nand GNAME6073(G6073,G4688,G5992);
  nand GNAME6074(G6074,G3705,G4182);
  nand GNAME6075(G6075,G6073,G6074);
  nand GNAME6076(G6076,G4593,G6010);
  nand GNAME6077(G6077,G3709,G4188);
  nand GNAME6078(G6078,G6076,G6077);
  nand GNAME6079(G6079,G4704,G6001);
  nand GNAME6080(G6080,G3719,G4185);
  nand GNAME6081(G6081,G6079,G6080);
  nand GNAME6082(G6082,G4614,G6004);
  nand GNAME6083(G6083,G3711,G4186);
  nand GNAME6084(G6084,G6082,G6083);
  nand GNAME6085(G6085,G4454,G6022);
  nand GNAME6086(G6086,G3717,G4192);
  nand GNAME6087(G6087,G6085,G6086);
  nand GNAME6088(G6088,G4699,G5983);
  nand GNAME6089(G6089,G3715,G4179);
  nand GNAME6090(G6090,G6088,G6089);
  nand GNAME6091(G6091,G4481,G6025);
  nand GNAME6092(G6092,G3721,G4193);
  nand GNAME6093(G6093,G6091,G6092);
  nand GNAME6094(G6094,G4449,G6037);
  nand GNAME6095(G6095,G3713,G4197);
  nand GNAME6096(G6096,G6094,G6095);
  nand GNAME6097(G6097,G4560,G6019);
  nand GNAME6098(G6098,G3743,G4191);
  nand GNAME6099(G6099,G6097,G6098);
  nand GNAME6100(G6100,G3691,G4100);
  or GNAME6101(G6101,G3691,G4100);
  nand GNAME6102(G6102,G6100,G6101);
  nand GNAME6103(G6103,G3687,G4094);
  or GNAME6104(G6104,G3687,G4094);
  nand GNAME6105(G6105,G6103,G6104);
  nand GNAME6106(G6106,G3681,G4101);
  or GNAME6107(G6107,G3681,G4101);
  nand GNAME6108(G6108,G6106,G6107);
  nand GNAME6109(G6109,G3689,G4092);
  or GNAME6110(G6110,G3689,G4092);
  nand GNAME6111(G6111,G6109,G6110);
  nand GNAME6112(G6112,G3699,G4099);
  or GNAME6113(G6113,G3699,G4099);
  nand GNAME6114(G6114,G6112,G6113);
  nand GNAME6115(G6115,G3703,G4098);
  or GNAME6116(G6116,G3703,G4098);
  nand GNAME6117(G6117,G6115,G6116);
  nand GNAME6118(G6118,G3697,G4093);
  or GNAME6119(G6119,G3697,G4093);
  nand GNAME6120(G6120,G6118,G6119);
  nand GNAME6121(G6121,G3693,G4096);
  or GNAME6122(G6122,G3693,G4096);
  nand GNAME6123(G6123,G6121,G6122);
  nand GNAME6124(G6124,G3685,G4102);
  or GNAME6125(G6125,G3685,G4102);
  nand GNAME6126(G6126,G6124,G6125);
  nand GNAME6127(G6127,G3701,G4095);
  or GNAME6128(G6128,G3701,G4095);
  nand GNAME6129(G6129,G6127,G6128);
  nand GNAME6130(G6130,G3683,G4103);
  or GNAME6131(G6131,G3683,G4103);
  nand GNAME6132(G6132,G6130,G6131);
  nand GNAME6133(G6133,G3695,G4097);
  or GNAME6134(G6134,G3695,G4097);
  nand GNAME6135(G6135,G6133,G6134);
  nand GNAME6136(G6136,G5941,G4358,G4078);
  nand GNAME6137(G6137,G4171,G6337,G4077);
  nand GNAME6138(G6138,G8728,G5941);
  nand GNAME6139(G6139,G4104,G4171);
  nand GNAME6140(G6140,G5941,G4772);
  nand GNAME6141(G6141,G4171,G5938,G6370);
  nand GNAME6142(G6142,G5962,G6138,G6139);
  nand GNAME6143(G6143,G4176,G4773,G6140,G6141);
  or GNAME6144(G6144,G8728,G4359);
  nand GNAME6145(G6145,G4368,G8728);
  nand GNAME6146(G6146,G4106,G23012);
  nand GNAME6147(G6147,G3681,G4365);
  nand GNAME6148(G6148,G4106,G23011);
  nand GNAME6149(G6149,G3683,G4365);
  nand GNAME6150(G6150,G4106,G23010);
  nand GNAME6151(G6151,G3685,G4365);
  nand GNAME6152(G6152,G4106,G23009);
  nand GNAME6153(G6153,G3687,G4365);
  nand GNAME6154(G6154,G4106,G23008);
  nand GNAME6155(G6155,G3689,G4365);
  nand GNAME6156(G6156,G4106,G23007);
  nand GNAME6157(G6157,G3691,G4365);
  nand GNAME6158(G6158,G4106,G23006);
  nand GNAME6159(G6159,G3693,G4365);
  nand GNAME6160(G6160,G4106,G23005);
  nand GNAME6161(G6161,G3695,G4365);
  nand GNAME6162(G6162,G4106,G23004);
  nand GNAME6163(G6163,G3697,G4365);
  nand GNAME6164(G6164,G4106,G23003);
  nand GNAME6165(G6165,G3699,G4365);
  nand GNAME6166(G6166,G4106,G23002);
  nand GNAME6167(G6167,G3701,G4365);
  nand GNAME6168(G6168,G4106,G23001);
  nand GNAME6169(G6169,G3703,G4365);
  nand GNAME6170(G6170,G4106,G23000);
  nand GNAME6171(G6171,G3705,G4365);
  nand GNAME6172(G6172,G4106,G22999);
  nand GNAME6173(G6173,G3707,G4365);
  nand GNAME6174(G6174,G4106,G22998);
  nand GNAME6175(G6175,G3709,G4365);
  nand GNAME6176(G6176,G4106,G22997);
  nand GNAME6177(G6177,G3711,G4365);
  nand GNAME6178(G6178,G4106,G22996);
  nand GNAME6179(G6179,G3713,G4365);
  nand GNAME6180(G6180,G4106,G22995);
  nand GNAME6181(G6181,G3715,G4365);
  nand GNAME6182(G6182,G4106,G22994);
  nand GNAME6183(G6183,G3717,G4365);
  nand GNAME6184(G6184,G4106,G22993);
  nand GNAME6185(G6185,G3719,G4365);
  nand GNAME6186(G6186,G4106,G22992);
  nand GNAME6187(G6187,G3721,G4365);
  nand GNAME6188(G6188,G4106,G22991);
  nand GNAME6189(G6189,G3723,G4365);
  nand GNAME6190(G6190,G4106,G22990);
  nand GNAME6191(G6191,G3725,G4365);
  nand GNAME6192(G6192,G4106,G22989);
  nand GNAME6193(G6193,G3727,G4365);
  nand GNAME6194(G6194,G4106,G22988);
  nand GNAME6195(G6195,G3729,G4365);
  nand GNAME6196(G6196,G4106,G22987);
  nand GNAME6197(G6197,G3731,G4365);
  nand GNAME6198(G6198,G4106,G22986);
  nand GNAME6199(G6199,G3733,G4365);
  nand GNAME6200(G6200,G4106,G22985);
  nand GNAME6201(G6201,G3735,G4365);
  nand GNAME6202(G6202,G4106,G22984);
  nand GNAME6203(G6203,G3737,G4365);
  nand GNAME6204(G6204,G4106,G22983);
  nand GNAME6205(G6205,G3739,G4365);
  nand GNAME6206(G6206,G4106,G22982);
  nand GNAME6207(G6207,G3741,G4365);
  nand GNAME6208(G6208,G4106,G22981);
  nand GNAME6209(G6209,G3743,G4365);
  nand GNAME6210(G6210,G4057,G4365);
  or GNAME6211(G6211,G4057,G4107,G4781);
  nand GNAME6212(G6212,G6210,G6211);
  nand GNAME6213(G6213,G5885,G4173);
  nand GNAME6214(G6214,G5886,G5971);
  nand GNAME6215(G6215,G4112,G22958);
  nand GNAME6216(G6216,G4889,G4360);
  nand GNAME6217(G6217,G4112,G22930);
  nand GNAME6218(G6218,G4889,G5068,G9072);
  nand GNAME6219(G6219,G5888,G4174);
  nand GNAME6220(G6220,G5887,G5974);
  nand GNAME6221(G6221,G4122,G22926);
  nand GNAME6222(G6222,G5081,G4360);
  nand GNAME6223(G6223,G5938,G4363);
  or GNAME6224(G6224,G4363,G5938);
  nand GNAME6225(G6225,G6223,G6224);
  nand GNAME6226(G6226,G4127,G22894);
  nand GNAME6227(G6227,G5240,G4360);
  nand GNAME6228(G6228,G4398,G4364);
  nand GNAME6229(G6229,G5392,G22834);
  nand GNAME6230(G6230,G4397,G4364);
  nand GNAME6231(G6231,G5392,G22833);
  nand GNAME6232(G6232,G9008,G8728);
  nand GNAME6233(G6233,G4104,G3725);
  nand GNAME6234(G6234,G9011,G8728);
  nand GNAME6235(G6235,G4104,G3727);
  nand GNAME6236(G6236,G8992,G8728);
  nand GNAME6237(G6237,G4104,G3729);
  nand GNAME6238(G6238,G8955,G8728);
  nand GNAME6239(G6239,G4104,G3731);
  nand GNAME6240(G6240,G9015,G8728);
  nand GNAME6241(G6241,G4104,G3733);
  nand GNAME6242(G6242,G9018,G8728);
  nand GNAME6243(G6243,G4104,G3735);
  nand GNAME6244(G6244,G8728,G8994);
  nand GNAME6245(G6245,G4104,G3681);
  nand GNAME6246(G6246,G8728,G8995);
  nand GNAME6247(G6247,G4104,G3683);
  nand GNAME6248(G6248,G8993,G8728);
  nand GNAME6249(G6249,G4104,G3737);
  nand GNAME6250(G6250,G8728,G9042);
  nand GNAME6251(G6251,G4104,G3685);
  nand GNAME6252(G6252,G9045,G8728);
  nand GNAME6253(G6253,G4104,G3687);
  nand GNAME6254(G6254,G9048,G8728);
  nand GNAME6255(G6255,G4104,G3689);
  nand GNAME6256(G6256,G9051,G8728);
  nand GNAME6257(G6257,G4104,G3691);
  nand GNAME6258(G6258,G9054,G8728);
  nand GNAME6259(G6259,G4104,G3693);
  nand GNAME6260(G6260,G9057,G8728);
  nand GNAME6261(G6261,G4104,G3695);
  nand GNAME6262(G6262,G9060,G8728);
  nand GNAME6263(G6263,G4104,G3697);
  nand GNAME6264(G6264,G9063,G8728);
  nand GNAME6265(G6265,G4104,G3699);
  nand GNAME6266(G6266,G9066,G8728);
  nand GNAME6267(G6267,G4104,G3701);
  nand GNAME6268(G6268,G9069,G8728);
  nand GNAME6269(G6269,G4104,G3703);
  nand GNAME6270(G6270,G8954,G8728);
  nand GNAME6271(G6271,G4104,G3739);
  nand GNAME6272(G6272,G9075,G8728);
  nand GNAME6273(G6273,G4104,G3705);
  nand GNAME6274(G6274,G9078,G8728);
  nand GNAME6275(G6275,G4104,G3707);
  nand GNAME6276(G6276,G9081,G8728);
  nand GNAME6277(G6277,G4104,G3709);
  nand GNAME6278(G6278,G9084,G8728);
  nand GNAME6279(G6279,G4104,G3711);
  nand GNAME6280(G6280,G9087,G8728);
  nand GNAME6281(G6281,G4104,G3713);
  nand GNAME6282(G6282,G8996,G8728);
  nand GNAME6283(G6283,G4104,G3715);
  nand GNAME6284(G6284,G9091,G8728);
  nand GNAME6285(G6285,G4104,G3717);
  nand GNAME6286(G6286,G9094,G8728);
  nand GNAME6287(G6287,G4104,G3719);
  nand GNAME6288(G6288,G8997,G8728);
  nand GNAME6289(G6289,G4104,G3721);
  nand GNAME6290(G6290,G8953,G8728);
  nand GNAME6291(G6291,G4104,G3723);
  nand GNAME6292(G6292,G9072,G8728);
  nand GNAME6293(G6293,G4104,G3741);
  nand GNAME6294(G6294,G8991,G8728);
  nand GNAME6295(G6295,G4104,G3743);
  nand GNAME6296(G6296,G22906,G5944);
  nand GNAME6297(G6297,G22938,G4172);
  nand GNAME6298(G6298,G22905,G5944);
  nand GNAME6299(G6299,G22937,G4172);
  nand GNAME6300(G6300,G22904,G5944);
  nand GNAME6301(G6301,G22936,G4172);
  nand GNAME6302(G6302,G22903,G5944);
  nand GNAME6303(G6303,G22935,G4172);
  nand GNAME6304(G6304,G22902,G5944);
  nand GNAME6305(G6305,G22934,G4172);
  nand GNAME6306(G6306,G22901,G5944);
  nand GNAME6307(G6307,G22933,G4172);
  nand GNAME6308(G6308,G22900,G5944);
  nand GNAME6309(G6309,G22932,G4172);
  nand GNAME6310(G6310,G22899,G5944);
  nand GNAME6311(G6311,G22931,G4172);
  nand GNAME6312(G6312,G22916,G5944);
  nand GNAME6313(G6313,G22948,G4172);
  nand GNAME6314(G6314,G22915,G5944);
  nand GNAME6315(G6315,G22947,G4172);
  nand GNAME6316(G6316,G22914,G5944);
  nand GNAME6317(G6317,G22946,G4172);
  nand GNAME6318(G6318,G22913,G5944);
  nand GNAME6319(G6319,G22945,G4172);
  nand GNAME6320(G6320,G22912,G5944);
  nand GNAME6321(G6321,G22944,G4172);
  nand GNAME6322(G6322,G22911,G5944);
  nand GNAME6323(G6323,G22943,G4172);
  nand GNAME6324(G6324,G22910,G5944);
  nand GNAME6325(G6325,G22942,G4172);
  nand GNAME6326(G6326,G22909,G5944);
  nand GNAME6327(G6327,G22941,G4172);
  nand GNAME6328(G6328,G22908,G5944);
  nand GNAME6329(G6329,G22940,G4172);
  nand GNAME6330(G6330,G22907,G5944);
  nand GNAME6331(G6331,G22939,G4172);
  nand GNAME6332(G6332,G22898,G5944);
  nand GNAME6333(G6333,G22930,G4172);
  nand GNAME6334(G6334,G22897,G5944);
  nand GNAME6335(G6335,G22929,G4172);
  not GNAME6336(G6336,G23013);
  not GNAME6337(G6337,G6370);
  not GNAME6338(G6338,G4263);
  not GNAME6339(G6339,G4101);
  not GNAME6340(G6340,G4103);
  not GNAME6341(G6341,G4241);
  not GNAME6342(G6342,G4094);
  not GNAME6343(G6343,G4243);
  not GNAME6344(G6344,G4100);
  not GNAME6345(G6345,G4245);
  not GNAME6346(G6346,G4097);
  not GNAME6347(G6347,G4247);
  not GNAME6348(G6348,G4099);
  not GNAME6349(G6349,G4249);
  not GNAME6350(G6350,G4098);
  not GNAME6351(G6351,G4252);
  not GNAME6352(G6352,G4195);
  not GNAME6353(G6353,G4254);
  not GNAME6354(G6354,G4186);
  not GNAME6355(G6355,G4256);
  not GNAME6356(G6356,G4179);
  not GNAME6357(G6357,G4258);
  not GNAME6358(G6358,G4185);
  not GNAME6359(G6359,G4260);
  not GNAME6360(G6360,G4180);
  not GNAME6361(G6361,G4232);
  not GNAME6362(G6362,G4183);
  not GNAME6363(G6363,G4234);
  not GNAME6364(G6364,G4196);
  not GNAME6365(G6365,G4236);
  not GNAME6366(G6366,G4189);
  not GNAME6367(G6367,G4240);
  not GNAME6368(G6368,G4194);
  not GNAME6369(G6369,G4262);
  nand GNAME6370(G6370,G848,G849);
  nand GNAME6371(G6371,G9403,G23038);
  nand GNAME6372(G6372,G9404,G23019);
  nand GNAME6373(G6373,G9405,G23031);
  nand GNAME6374(G6374,G9406,G23021);
  nand GNAME6375(G6375,G9407,G23040);
  nand GNAME6376(G6376,G9408,G23014);
  nand GNAME6377(G6377,G9409,G23029);
  nand GNAME6378(G6378,G9410,G23027);
  nand GNAME6379(G6379,G9411,G23017);
  nand GNAME6380(G6380,G9412,G23036);
  nand GNAME6381(G6381,G9413,G23022);
  nand GNAME6382(G6382,G9414,G23032);
  nand GNAME6383(G6383,G9415,G23020);
  nand GNAME6384(G6384,G9416,G23039);
  nand GNAME6385(G6385,G9417,G23026);
  nand GNAME6386(G6386,G9418,G23030);
  nand GNAME6387(G6387,G9419,G23015);
  nand GNAME6388(G6388,G6398,G23041);
  and GNAME6389(G6389,G6397,G23035);
  nand GNAME6390(G6390,G23037,G23025);
  nand GNAME6391(G6391,G9398,G23028);
  nand GNAME6392(G6392,G9399,G23016);
  nand GNAME6393(G6393,G9400,G23042);
  nand GNAME6394(G6394,G9401,G23034);
  nand GNAME6395(G6395,G9402,G23024);
  nor GNAME6396(G6396,G23035,G6397);
  or GNAME6397(G6397,G23041,G6398);
  or GNAME6398(G6398,G23015,G9419);
  and GNAME6399(G6399,G6623,G6624);
  and GNAME6400(G6400,G6619,G6621);
  and GNAME6401(G6401,G6617,G6618);
  and GNAME6402(G6402,G6613,G6615);
  and GNAME6403(G6403,G6611,G6612);
  and GNAME6404(G6404,G6606,G6608);
  nand GNAME6405(G6405,G6628,G6716,G6717);
  not GNAME6406(G6406,G642);
  nand GNAME6407(G6407,G32,G642);
  not GNAME6408(G6408,G31);
  not GNAME6409(G6409,G630);
  not GNAME6410(G6410,G30);
  not GNAME6411(G6411,G619);
  not GNAME6412(G6412,G29);
  not GNAME6413(G6413,G613);
  not GNAME6414(G6414,G25);
  not GNAME6415(G6415,G612);
  not GNAME6416(G6416,G24);
  not GNAME6417(G6417,G23);
  not GNAME6418(G6418,G611);
  not GNAME6419(G6419,G17);
  not GNAME6420(G6420,G21);
  not GNAME6421(G6421,G638);
  not GNAME6422(G6422,G20);
  not GNAME6423(G6423,G637);
  not GNAME6424(G6424,G19);
  not GNAME6425(G6425,G634);
  not GNAME6426(G6426,G16);
  not GNAME6427(G6427,G633);
  not GNAME6428(G6428,G15);
  not GNAME6429(G6429,G632);
  not GNAME6430(G6430,G14);
  not GNAME6431(G6431,G631);
  not GNAME6432(G6432,G13);
  not GNAME6433(G6433,G629);
  not GNAME6434(G6434,G12);
  not GNAME6435(G6435,G628);
  not GNAME6436(G6436,G11);
  not GNAME6437(G6437,G627);
  not GNAME6438(G6438,G10);
  not GNAME6439(G6439,G626);
  not GNAME6440(G6440,G9);
  not GNAME6441(G6441,G625);
  not GNAME6442(G6442,G8);
  not GNAME6443(G6443,G624);
  not GNAME6444(G6444,G7);
  not GNAME6445(G6445,G623);
  not GNAME6446(G6446,G6);
  not GNAME6447(G6447,G4);
  not GNAME6448(G6448,G621);
  nor GNAME6449(G6449,G6754,G6456);
  not GNAME6450(G6450,G3);
  not GNAME6451(G6451,G620);
  and GNAME6452(G6452,G6600,G6601);
  not GNAME6453(G6453,G2);
  not GNAME6454(G6454,G618);
  and GNAME6455(G6455,G6592,G6593);
  nor GNAME6456(G6456,G6594,G6455);
  and GNAME6457(G6457,G6558,G6559);
  and GNAME6458(G6458,G6555,G6556);
  or GNAME6459(G6459,G6557,G6458);
  and GNAME6460(G6460,G6548,G6549);
  and GNAME6461(G6461,G6545,G6546);
  or GNAME6462(G6462,G6547,G6461);
  nand GNAME6463(G6463,G6752,G6753);
  nand GNAME6464(G6464,G6632,G6633);
  nand GNAME6465(G6465,G6637,G6638);
  nand GNAME6466(G6466,G6642,G6643);
  nand GNAME6467(G6467,G6644,G6645);
  nand GNAME6468(G6468,G6646,G6647);
  nand GNAME6469(G6469,G6648,G6649);
  nand GNAME6470(G6470,G6653,G6654);
  nand GNAME6471(G6471,G6661,G6662);
  nand GNAME6472(G6472,G6666,G6667);
  nand GNAME6473(G6473,G6671,G6672);
  nand GNAME6474(G6474,G6676,G6677);
  nand GNAME6475(G6475,G6681,G6682);
  nand GNAME6476(G6476,G6686,G6687);
  nand GNAME6477(G6477,G6691,G6692);
  nand GNAME6478(G6478,G6696,G6697);
  nand GNAME6479(G6479,G6701,G6702);
  nand GNAME6480(G6480,G6706,G6707);
  nand GNAME6481(G6481,G6711,G6712);
  nand GNAME6482(G6482,G6721,G6722);
  nand GNAME6483(G6483,G6726,G6727);
  nand GNAME6484(G6484,G6731,G6732);
  nand GNAME6485(G6485,G6736,G6737);
  nand GNAME6486(G6486,G6743,G6744);
  nand GNAME6487(G6487,G6748,G6749);
  nand GNAME6488(G6488,G6537,G6538);
  nand GNAME6489(G6489,G6534,G6535);
  nand GNAME6490(G6490,G6539,G6532);
  and GNAME6491(G6491,G6529,G6527);
  and GNAME6492(G6492,G6540,G6525);
  and GNAME6493(G6493,G6521,G6522);
  nand GNAME6494(G6494,G6518,G6519);
  not GNAME6495(G6495,G1);
  not GNAME6496(G6496,G617);
  or GNAME6497(G6497,G6516,G6506);
  and GNAME6498(G6498,G6596,G6597);
  nand GNAME6499(G6499,G6589,G6590);
  nand GNAME6500(G6500,G6586,G6587);
  nand GNAME6501(G6501,G6583,G6584);
  nand GNAME6502(G6502,G6580,G6581);
  nand GNAME6503(G6503,G6577,G6578);
  nand GNAME6504(G6504,G6574,G6575);
  nand GNAME6505(G6505,G6571,G6572);
  nor GNAME6506(G6506,G6407,G6408);
  nand GNAME6507(G6507,G6568,G6569);
  nand GNAME6508(G6508,G6565,G6566);
  nand GNAME6509(G6509,G6562,G6563);
  or GNAME6510(G6510,G6560,G6457);
  nand GNAME6511(G6511,G6552,G6553);
  or GNAME6512(G6512,G6550,G6460);
  not GNAME6513(G6513,G6449);
  not GNAME6514(G6514,G6407);
  or GNAME6515(G6515,G6514,G31);
  and GNAME6516(G6516,G6515,G641);
  nand GNAME6517(G6517,G6410,G6409);
  nand GNAME6518(G6518,G6497,G6517);
  or GNAME6519(G6519,G6409,G6410);
  nand GNAME6520(G6520,G6412,G6411);
  nand GNAME6521(G6521,G6494,G6520);
  or GNAME6522(G6522,G6411,G6412);
  not GNAME6523(G6523,G6493);
  or GNAME6524(G6524,G616,G28);
  nand GNAME6525(G6525,G6523,G6524);
  not GNAME6526(G6526,G6492);
  nand GNAME6527(G6527,G615,G27);
  or GNAME6528(G6528,G27,G615);
  nand GNAME6529(G6529,G6526,G6528);
  not GNAME6530(G6530,G6491);
  or GNAME6531(G6531,G26,G614);
  nand GNAME6532(G6532,G6530,G6531);
  nand GNAME6533(G6533,G6414,G6413);
  nand GNAME6534(G6534,G6490,G6533);
  or GNAME6535(G6535,G6413,G6414);
  nand GNAME6536(G6536,G6416,G6415);
  nand GNAME6537(G6537,G6489,G6536);
  or GNAME6538(G6538,G6415,G6416);
  nand GNAME6539(G6539,G614,G26);
  nand GNAME6540(G6540,G28,G616);
  nand GNAME6541(G6541,G622,G5);
  and GNAME6542(G6542,G636,G18);
  and GNAME6543(G6543,G640,G22);
  nand GNAME6544(G6544,G6417,G6418);
  nand GNAME6545(G6545,G6488,G6544);
  or GNAME6546(G6546,G6417,G6418);
  nor GNAME6547(G6547,G22,G640);
  nand GNAME6548(G6548,G6756,G6462);
  or GNAME6549(G6549,G639,G21);
  and GNAME6550(G6550,G639,G21);
  nand GNAME6551(G6551,G6422,G6421);
  nand GNAME6552(G6552,G6512,G6551);
  or GNAME6553(G6553,G6421,G6422);
  nand GNAME6554(G6554,G6424,G6423);
  nand GNAME6555(G6555,G6511,G6554);
  or GNAME6556(G6556,G6423,G6424);
  nor GNAME6557(G6557,G18,G636);
  nand GNAME6558(G6558,G6755,G6459);
  or GNAME6559(G6559,G635,G17);
  and GNAME6560(G6560,G635,G17);
  nand GNAME6561(G6561,G6426,G6425);
  nand GNAME6562(G6562,G6510,G6561);
  or GNAME6563(G6563,G6425,G6426);
  nand GNAME6564(G6564,G6428,G6427);
  nand GNAME6565(G6565,G6509,G6564);
  or GNAME6566(G6566,G6427,G6428);
  nand GNAME6567(G6567,G6430,G6429);
  nand GNAME6568(G6568,G6508,G6567);
  or GNAME6569(G6569,G6429,G6430);
  nand GNAME6570(G6570,G6432,G6431);
  nand GNAME6571(G6571,G6507,G6570);
  or GNAME6572(G6572,G6431,G6432);
  nand GNAME6573(G6573,G6434,G6433);
  nand GNAME6574(G6574,G6505,G6573);
  or GNAME6575(G6575,G6433,G6434);
  nand GNAME6576(G6576,G6436,G6435);
  nand GNAME6577(G6577,G6504,G6576);
  or GNAME6578(G6578,G6435,G6436);
  nand GNAME6579(G6579,G6438,G6437);
  nand GNAME6580(G6580,G6503,G6579);
  or GNAME6581(G6581,G6437,G6438);
  nand GNAME6582(G6582,G6440,G6439);
  nand GNAME6583(G6583,G6502,G6582);
  or GNAME6584(G6584,G6439,G6440);
  nand GNAME6585(G6585,G6442,G6441);
  nand GNAME6586(G6586,G6501,G6585);
  or GNAME6587(G6587,G6441,G6442);
  nand GNAME6588(G6588,G6444,G6443);
  nand GNAME6589(G6589,G6500,G6588);
  or GNAME6590(G6590,G6443,G6444);
  nand GNAME6591(G6591,G6446,G6445);
  nand GNAME6592(G6592,G6499,G6591);
  or GNAME6593(G6593,G6445,G6446);
  nor GNAME6594(G6594,G622,G5);
  or GNAME6595(G6595,G6447,G6448);
  nand GNAME6596(G6596,G6595,G6449);
  nand GNAME6597(G6597,G6447,G6448);
  not GNAME6598(G6598,G6498);
  or GNAME6599(G6599,G6450,G6451);
  nand GNAME6600(G6600,G6598,G6599);
  nand GNAME6601(G6601,G6450,G6451);
  not GNAME6602(G6602,G6452);
  nand GNAME6603(G6603,G6454,G6453);
  nand GNAME6604(G6604,G6603,G6452);
  or GNAME6605(G6605,G6453,G6454);
  nand GNAME6606(G6606,G6655,G6656,G6604,G6605);
  nand GNAME6607(G6607,G6602,G6605);
  nand GNAME6608(G6608,G6657,G6607,G6603);
  or GNAME6609(G6609,G5,G622);
  nand GNAME6610(G6610,G6541,G6609);
  nand GNAME6611(G6611,G6610,G6455);
  nand GNAME6612(G6612,G6541,G6456);
  nand GNAME6613(G6613,G6738,G6739,G6755,G6459);
  nand GNAME6614(G6614,G635,G17);
  nand GNAME6615(G6615,G6614,G6457);
  or GNAME6616(G6616,G6542,G6557);
  nand GNAME6617(G6617,G6616,G6458);
  or GNAME6618(G6618,G6542,G6459);
  nand GNAME6619(G6619,G6750,G6751,G6756,G6462);
  nand GNAME6620(G6620,G639,G21);
  nand GNAME6621(G6621,G6620,G6460);
  or GNAME6622(G6622,G6543,G6547);
  nand GNAME6623(G6623,G6622,G6461);
  or GNAME6624(G6624,G6543,G6462);
  nand GNAME6625(G6625,G6531,G6539);
  nand GNAME6626(G6626,G6527,G6528);
  nand GNAME6627(G6627,G6524,G6540);
  nand GNAME6628(G6628,G6408,G6715);
  or GNAME6629(G6629,G611,G6417);
  or GNAME6630(G6630,G23,G6418);
  and GNAME6631(G6631,G6629,G6630);
  nand GNAME6632(G6632,G6488,G6629,G6630);
  or GNAME6633(G6633,G6631,G6488);
  or GNAME6634(G6634,G612,G6416);
  or GNAME6635(G6635,G24,G6415);
  and GNAME6636(G6636,G6634,G6635);
  nand GNAME6637(G6637,G6489,G6634,G6635);
  or GNAME6638(G6638,G6636,G6489);
  or GNAME6639(G6639,G613,G6414);
  or GNAME6640(G6640,G25,G6413);
  and GNAME6641(G6641,G6639,G6640);
  nand GNAME6642(G6642,G6490,G6639,G6640);
  or GNAME6643(G6643,G6641,G6490);
  nand GNAME6644(G6644,G6530,G6625);
  nand GNAME6645(G6645,G6491,G6531,G6539);
  nand GNAME6646(G6646,G6526,G6626);
  nand GNAME6647(G6647,G6492,G6527,G6528);
  nand GNAME6648(G6648,G6523,G6627);
  nand GNAME6649(G6649,G6493,G6524,G6540);
  or GNAME6650(G6650,G619,G6412);
  or GNAME6651(G6651,G29,G6411);
  and GNAME6652(G6652,G6650,G6651);
  nand GNAME6653(G6653,G6494,G6650,G6651);
  or GNAME6654(G6654,G6652,G6494);
  or GNAME6655(G6655,G617,G6495);
  or GNAME6656(G6656,G1,G6496);
  nand GNAME6657(G6657,G6655,G6656);
  or GNAME6658(G6658,G2,G6454);
  or GNAME6659(G6659,G618,G6453);
  nand GNAME6660(G6660,G6658,G6659);
  nand GNAME6661(G6661,G6602,G6660);
  nand GNAME6662(G6662,G6452,G6658,G6659);
  or GNAME6663(G6663,G630,G6410);
  or GNAME6664(G6664,G30,G6409);
  and GNAME6665(G6665,G6663,G6664);
  nand GNAME6666(G6666,G6497,G6663,G6664);
  or GNAME6667(G6667,G6665,G6497);
  or GNAME6668(G6668,G3,G6451);
  or GNAME6669(G6669,G620,G6450);
  nand GNAME6670(G6670,G6668,G6669);
  nand GNAME6671(G6671,G6598,G6670);
  nand GNAME6672(G6672,G6498,G6668,G6669);
  or GNAME6673(G6673,G4,G6448);
  or GNAME6674(G6674,G621,G6447);
  nand GNAME6675(G6675,G6673,G6674);
  nand GNAME6676(G6676,G6513,G6673,G6674);
  nand GNAME6677(G6677,G6449,G6675);
  or GNAME6678(G6678,G623,G6446);
  or GNAME6679(G6679,G6,G6445);
  and GNAME6680(G6680,G6678,G6679);
  nand GNAME6681(G6681,G6499,G6678,G6679);
  or GNAME6682(G6682,G6680,G6499);
  or GNAME6683(G6683,G624,G6444);
  or GNAME6684(G6684,G7,G6443);
  and GNAME6685(G6685,G6683,G6684);
  nand GNAME6686(G6686,G6500,G6683,G6684);
  or GNAME6687(G6687,G6685,G6500);
  or GNAME6688(G6688,G625,G6442);
  or GNAME6689(G6689,G8,G6441);
  and GNAME6690(G6690,G6688,G6689);
  nand GNAME6691(G6691,G6501,G6688,G6689);
  or GNAME6692(G6692,G6690,G6501);
  or GNAME6693(G6693,G626,G6440);
  or GNAME6694(G6694,G9,G6439);
  and GNAME6695(G6695,G6693,G6694);
  nand GNAME6696(G6696,G6502,G6693,G6694);
  or GNAME6697(G6697,G6695,G6502);
  or GNAME6698(G6698,G627,G6438);
  or GNAME6699(G6699,G10,G6437);
  and GNAME6700(G6700,G6698,G6699);
  nand GNAME6701(G6701,G6503,G6698,G6699);
  or GNAME6702(G6702,G6700,G6503);
  or GNAME6703(G6703,G628,G6436);
  or GNAME6704(G6704,G11,G6435);
  and GNAME6705(G6705,G6703,G6704);
  nand GNAME6706(G6706,G6504,G6703,G6704);
  or GNAME6707(G6707,G6705,G6504);
  or GNAME6708(G6708,G629,G6434);
  or GNAME6709(G6709,G12,G6433);
  and GNAME6710(G6710,G6708,G6709);
  nand GNAME6711(G6711,G6505,G6708,G6709);
  or GNAME6712(G6712,G6710,G6505);
  nand GNAME6713(G6713,G6407,G641);
  or GNAME6714(G6714,G641,G6407);
  nand GNAME6715(G6715,G6713,G6714);
  or GNAME6716(G6716,G641,G6514,G6408);
  nand GNAME6717(G6717,G641,G6506);
  or GNAME6718(G6718,G631,G6432);
  or GNAME6719(G6719,G13,G6431);
  and GNAME6720(G6720,G6718,G6719);
  nand GNAME6721(G6721,G6507,G6718,G6719);
  or GNAME6722(G6722,G6720,G6507);
  or GNAME6723(G6723,G632,G6430);
  or GNAME6724(G6724,G14,G6429);
  and GNAME6725(G6725,G6723,G6724);
  nand GNAME6726(G6726,G6508,G6723,G6724);
  or GNAME6727(G6727,G6725,G6508);
  or GNAME6728(G6728,G633,G6428);
  or GNAME6729(G6729,G15,G6427);
  and GNAME6730(G6730,G6728,G6729);
  nand GNAME6731(G6731,G6509,G6728,G6729);
  or GNAME6732(G6732,G6730,G6509);
  or GNAME6733(G6733,G634,G6426);
  or GNAME6734(G6734,G16,G6425);
  and GNAME6735(G6735,G6733,G6734);
  nand GNAME6736(G6736,G6510,G6733,G6734);
  or GNAME6737(G6737,G6735,G6510);
  or GNAME6738(G6738,G635,G6419);
  nand GNAME6739(G6739,G6419,G635);
  or GNAME6740(G6740,G637,G6424);
  or GNAME6741(G6741,G19,G6423);
  and GNAME6742(G6742,G6740,G6741);
  nand GNAME6743(G6743,G6511,G6740,G6741);
  or GNAME6744(G6744,G6742,G6511);
  or GNAME6745(G6745,G638,G6422);
  or GNAME6746(G6746,G20,G6421);
  and GNAME6747(G6747,G6745,G6746);
  nand GNAME6748(G6748,G6512,G6745,G6746);
  or GNAME6749(G6749,G6747,G6512);
  or GNAME6750(G6750,G639,G6420);
  nand GNAME6751(G6751,G6420,G639);
  or GNAME6752(G6752,G32,G6406);
  nand GNAME6753(G6753,G6406,G32);
  not GNAME6754(G6754,G6541);
  not GNAME6755(G6755,G6542);
  not GNAME6756(G6756,G6543);
  not GNAME6757(G6757,G22716);
  and GNAME6758(G6758,G6895,G6896);
  and GNAME6759(G6759,G6891,G6893);
  and GNAME6760(G6760,G6888,G6890);
  and GNAME6761(G6761,G6886,G6887);
  and GNAME6762(G6762,G6881,G6883);
  nand GNAME6763(G6763,G6900,G6935,G6936);
  not GNAME6764(G6764,G22735);
  nand GNAME6765(G6765,G22980,G22735);
  not GNAME6766(G6766,G22979);
  not GNAME6767(G6767,G22733);
  not GNAME6768(G6768,G22978);
  not GNAME6769(G6769,G22732);
  not GNAME6770(G6770,G22977);
  not GNAME6771(G6771,G22728);
  not GNAME6772(G6772,G22973);
  not GNAME6773(G6773,G22727);
  not GNAME6774(G6774,G22972);
  not GNAME6775(G6775,G22971);
  not GNAME6776(G6776,G22726);
  not GNAME6777(G6777,G22969);
  not GNAME6778(G6778,G22723);
  not GNAME6779(G6779,G22968);
  not GNAME6780(G6780,G22722);
  not GNAME6781(G6781,G22967);
  not GNAME6782(G6782,G22964);
  not GNAME6783(G6783,G22719);
  nor GNAME6784(G6784,G6969,G6790);
  not GNAME6785(G6785,G22963);
  not GNAME6786(G6786,G22718);
  and GNAME6787(G6787,G6875,G6876);
  not GNAME6788(G6788,G22962);
  not GNAME6789(G6789,G22717);
  and GNAME6790(G6790,G6869,G6884);
  or GNAME6791(G6791,G6868,G6792);
  and GNAME6792(G6792,G6866,G6867);
  and GNAME6793(G6793,G6859,G6860);
  and GNAME6794(G6794,G6856,G6857);
  or GNAME6795(G6795,G6858,G6794);
  nand GNAME6796(G6796,G6967,G6968);
  nand GNAME6797(G6797,G6904,G6905);
  nand GNAME6798(G6798,G6909,G6910);
  nand GNAME6799(G6799,G6914,G6915);
  nand GNAME6800(G6800,G6916,G6917);
  nand GNAME6801(G6801,G6918,G6919);
  nand GNAME6802(G6802,G6920,G6921);
  nand GNAME6803(G6803,G6925,G6926);
  nand GNAME6804(G6804,G6930,G6931);
  nand GNAME6805(G6805,G6943,G6944);
  nand GNAME6806(G6806,G6948,G6949);
  nand GNAME6807(G6807,G6953,G6954);
  nand GNAME6808(G6808,G6958,G6959);
  nand GNAME6809(G6809,G6963,G6964);
  nand GNAME6810(G6810,G6848,G6849);
  nand GNAME6811(G6811,G6845,G6846);
  nand GNAME6812(G6812,G6850,G6843);
  and GNAME6813(G6813,G6840,G6838);
  and GNAME6814(G6814,G6851,G6836);
  and GNAME6815(G6815,G6832,G6833);
  nand GNAME6816(G6816,G6829,G6830);
  or GNAME6817(G6817,G6827,G6818);
  nor GNAME6818(G6818,G6765,G6766);
  not GNAME6819(G6819,G22961);
  not GNAME6820(G6820,G22716);
  and GNAME6821(G6821,G6871,G6872);
  nand GNAME6822(G6822,G6863,G6864);
  or GNAME6823(G6823,G6861,G6793);
  not GNAME6824(G6824,G6784);
  not GNAME6825(G6825,G6765);
  or GNAME6826(G6826,G6825,G22979);
  and GNAME6827(G6827,G6826,G22734);
  nand GNAME6828(G6828,G6768,G6767);
  nand GNAME6829(G6829,G6817,G6828);
  or GNAME6830(G6830,G6767,G6768);
  nand GNAME6831(G6831,G6770,G6769);
  nand GNAME6832(G6832,G6816,G6831);
  or GNAME6833(G6833,G6769,G6770);
  not GNAME6834(G6834,G6815);
  or GNAME6835(G6835,G22731,G22976);
  nand GNAME6836(G6836,G6834,G6835);
  not GNAME6837(G6837,G6814);
  nand GNAME6838(G6838,G22730,G22975);
  or GNAME6839(G6839,G22975,G22730);
  nand GNAME6840(G6840,G6837,G6839);
  not GNAME6841(G6841,G6813);
  or GNAME6842(G6842,G22974,G22729);
  nand GNAME6843(G6843,G6841,G6842);
  nand GNAME6844(G6844,G6772,G6771);
  nand GNAME6845(G6845,G6812,G6844);
  or GNAME6846(G6846,G6771,G6772);
  nand GNAME6847(G6847,G6774,G6773);
  nand GNAME6848(G6848,G6811,G6847);
  or GNAME6849(G6849,G6773,G6774);
  nand GNAME6850(G6850,G22729,G22974);
  nand GNAME6851(G6851,G22976,G22731);
  nand GNAME6852(G6852,G22720,G22965);
  and GNAME6853(G6853,G22721,G22966);
  and GNAME6854(G6854,G22725,G22970);
  nand GNAME6855(G6855,G6775,G6776);
  nand GNAME6856(G6856,G6810,G6855);
  or GNAME6857(G6857,G6775,G6776);
  nor GNAME6858(G6858,G22970,G22725);
  nand GNAME6859(G6859,G6971,G6795);
  or GNAME6860(G6860,G22724,G22969);
  and GNAME6861(G6861,G22724,G22969);
  nand GNAME6862(G6862,G6779,G6778);
  nand GNAME6863(G6863,G6823,G6862);
  or GNAME6864(G6864,G6778,G6779);
  nand GNAME6865(G6865,G6781,G6780);
  nand GNAME6866(G6866,G6822,G6865);
  or GNAME6867(G6867,G6780,G6781);
  nor GNAME6868(G6868,G22966,G22721);
  nand GNAME6869(G6869,G6970,G6791);
  or GNAME6870(G6870,G6782,G6783);
  nand GNAME6871(G6871,G6870,G6784);
  nand GNAME6872(G6872,G6782,G6783);
  not GNAME6873(G6873,G6821);
  or GNAME6874(G6874,G6785,G6786);
  nand GNAME6875(G6875,G6873,G6874);
  nand GNAME6876(G6876,G6785,G6786);
  not GNAME6877(G6877,G6787);
  nand GNAME6878(G6878,G6789,G6788);
  nand GNAME6879(G6879,G6878,G6787);
  or GNAME6880(G6880,G6788,G6789);
  nand GNAME6881(G6881,G6937,G6938,G6879,G6880);
  nand GNAME6882(G6882,G6877,G6880);
  nand GNAME6883(G6883,G6939,G6882,G6878);
  or GNAME6884(G6884,G22965,G22720);
  nand GNAME6885(G6885,G6852,G6884);
  nand GNAME6886(G6886,G6885,G6970,G6791);
  nand GNAME6887(G6887,G6852,G6790);
  or GNAME6888(G6888,G6853,G6791);
  or GNAME6889(G6889,G6853,G6868);
  nand GNAME6890(G6890,G6889,G6792);
  nand GNAME6891(G6891,G6965,G6966,G6971,G6795);
  nand GNAME6892(G6892,G22724,G22969);
  nand GNAME6893(G6893,G6892,G6793);
  or GNAME6894(G6894,G6854,G6858);
  nand GNAME6895(G6895,G6894,G6794);
  or GNAME6896(G6896,G6854,G6795);
  nand GNAME6897(G6897,G6842,G6850);
  nand GNAME6898(G6898,G6838,G6839);
  nand GNAME6899(G6899,G6835,G6851);
  nand GNAME6900(G6900,G6766,G6934);
  or GNAME6901(G6901,G22726,G6775);
  or GNAME6902(G6902,G22971,G6776);
  and GNAME6903(G6903,G6901,G6902);
  nand GNAME6904(G6904,G6810,G6901,G6902);
  or GNAME6905(G6905,G6903,G6810);
  or GNAME6906(G6906,G22727,G6774);
  or GNAME6907(G6907,G22972,G6773);
  and GNAME6908(G6908,G6906,G6907);
  nand GNAME6909(G6909,G6811,G6906,G6907);
  or GNAME6910(G6910,G6908,G6811);
  or GNAME6911(G6911,G22728,G6772);
  or GNAME6912(G6912,G22973,G6771);
  and GNAME6913(G6913,G6911,G6912);
  nand GNAME6914(G6914,G6812,G6911,G6912);
  or GNAME6915(G6915,G6913,G6812);
  nand GNAME6916(G6916,G6841,G6897);
  nand GNAME6917(G6917,G6813,G6842,G6850);
  nand GNAME6918(G6918,G6837,G6898);
  nand GNAME6919(G6919,G6814,G6838,G6839);
  nand GNAME6920(G6920,G6834,G6899);
  nand GNAME6921(G6921,G6815,G6835,G6851);
  or GNAME6922(G6922,G22732,G6770);
  or GNAME6923(G6923,G22977,G6769);
  and GNAME6924(G6924,G6922,G6923);
  nand GNAME6925(G6925,G6816,G6922,G6923);
  or GNAME6926(G6926,G6924,G6816);
  or GNAME6927(G6927,G22733,G6768);
  or GNAME6928(G6928,G22978,G6767);
  and GNAME6929(G6929,G6927,G6928);
  nand GNAME6930(G6930,G6817,G6927,G6928);
  or GNAME6931(G6931,G6929,G6817);
  nand GNAME6932(G6932,G6765,G22734);
  or GNAME6933(G6933,G22734,G6765);
  nand GNAME6934(G6934,G6932,G6933);
  or GNAME6935(G6935,G22734,G6825,G6766);
  nand GNAME6936(G6936,G22734,G6818);
  or GNAME6937(G6937,G22716,G6819);
  or GNAME6938(G6938,G22961,G6820);
  nand GNAME6939(G6939,G6937,G6938);
  or GNAME6940(G6940,G22962,G6789);
  or GNAME6941(G6941,G22717,G6788);
  nand GNAME6942(G6942,G6940,G6941);
  nand GNAME6943(G6943,G6877,G6942);
  nand GNAME6944(G6944,G6787,G6940,G6941);
  or GNAME6945(G6945,G22963,G6786);
  or GNAME6946(G6946,G22718,G6785);
  nand GNAME6947(G6947,G6945,G6946);
  nand GNAME6948(G6948,G6873,G6947);
  nand GNAME6949(G6949,G6821,G6945,G6946);
  or GNAME6950(G6950,G22964,G6783);
  or GNAME6951(G6951,G22719,G6782);
  nand GNAME6952(G6952,G6950,G6951);
  nand GNAME6953(G6953,G6824,G6950,G6951);
  nand GNAME6954(G6954,G6784,G6952);
  or GNAME6955(G6955,G22722,G6781);
  or GNAME6956(G6956,G22967,G6780);
  and GNAME6957(G6957,G6955,G6956);
  nand GNAME6958(G6958,G6822,G6955,G6956);
  or GNAME6959(G6959,G6957,G6822);
  or GNAME6960(G6960,G22723,G6779);
  or GNAME6961(G6961,G22968,G6778);
  and GNAME6962(G6962,G6960,G6961);
  nand GNAME6963(G6963,G6823,G6960,G6961);
  or GNAME6964(G6964,G6962,G6823);
  or GNAME6965(G6965,G22724,G6777);
  nand GNAME6966(G6966,G6777,G22724);
  or GNAME6967(G6967,G22980,G6764);
  nand GNAME6968(G6968,G6764,G22980);
  not GNAME6969(G6969,G6852);
  not GNAME6970(G6970,G6853);
  not GNAME6971(G6971,G6854);
  not GNAME6972(G6972,G22961);
  and GNAME6973(G6973,G7238,G7239);
  and GNAME6974(G6974,G7234,G7235);
  and GNAME6975(G6975,G7159,G7160);
  not GNAME6976(G6976,G869);
  not GNAME6977(G6977,G928);
  not GNAME6978(G6978,G929);
  not GNAME6979(G6979,G932);
  not GNAME6980(G6980,G933);
  not GNAME6981(G6981,G934);
  not GNAME6982(G6982,G931);
  not GNAME6983(G6983,G930);
  not GNAME6984(G6984,G927);
  not GNAME6985(G6985,G926);
  not GNAME6986(G6986,G925);
  and GNAME6987(G6987,G7147,G7117);
  not GNAME6988(G6988,G924);
  not GNAME6989(G6989,G923);
  not GNAME6990(G6990,G922);
  not GNAME6991(G6991,G921);
  not GNAME6992(G6992,G920);
  not GNAME6993(G6993,G919);
  not GNAME6994(G6994,G918);
  not GNAME6995(G6995,G917);
  not GNAME6996(G6996,G916);
  not GNAME6997(G6997,G915);
  not GNAME6998(G6998,G914);
  not GNAME6999(G6999,G913);
  not GNAME7000(G7000,G912);
  not GNAME7001(G7001,G911);
  not GNAME7002(G7002,G910);
  not GNAME7003(G7003,G909);
  not GNAME7004(G7004,G908);
  not GNAME7005(G7005,G907);
  not GNAME7006(G7006,G906);
  not GNAME7007(G7007,G903);
  and GNAME7008(G7008,G7139,G7119);
  and GNAME7009(G7009,G7188,G7121);
  and GNAME7010(G7010,G7333,G7334);
  nand GNAME7011(G7011,G7383,G7384);
  nand GNAME7012(G7012,G7274,G7275);
  nand GNAME7013(G7013,G7280,G7281);
  nand GNAME7014(G7014,G7339,G7340);
  nand GNAME7015(G7015,G7341,G7342);
  nand GNAME7016(G7016,G7375,G7376);
  nand GNAME7017(G7017,G7381,G7382);
  not GNAME7018(G7018,G893);
  not GNAME7019(G7019,G895);
  not GNAME7020(G7020,G897);
  not GNAME7021(G7021,G899);
  not GNAME7022(G7022,G900);
  not GNAME7023(G7023,G896);
  not GNAME7024(G7024,G892);
  not GNAME7025(G7025,G891);
  nand GNAME7026(G7026,G7154,G7152);
  and GNAME7027(G7027,G7156,G7155);
  and GNAME7028(G7028,G7270,G7271);
  nand GNAME7029(G7029,G7151,G7124);
  and GNAME7030(G7030,G7153,G7152);
  and GNAME7031(G7031,G7272,G7273);
  nor GNAME7032(G7032,G7386,G6987);
  nand GNAME7033(G7033,G7145,G7129);
  and GNAME7034(G7034,G7146,G7126);
  and GNAME7035(G7035,G7276,G7277);
  nand GNAME7036(G7036,G7143,G7130);
  and GNAME7037(G7037,G7144,G7129);
  and GNAME7038(G7038,G7278,G7279);
  nor GNAME7039(G7039,G7385,G7008);
  not GNAME7040(G7040,G889);
  not GNAME7041(G7041,G888);
  not GNAME7042(G7042,G887);
  not GNAME7043(G7043,G885);
  not GNAME7044(G7044,G884);
  not GNAME7045(G7045,G883);
  not GNAME7046(G7046,G882);
  not GNAME7047(G7047,G881);
  not GNAME7048(G7048,G880);
  not GNAME7049(G7049,G879);
  not GNAME7050(G7050,G878);
  not GNAME7051(G7051,G877);
  not GNAME7052(G7052,G876);
  not GNAME7053(G7053,G875);
  not GNAME7054(G7054,G874);
  not GNAME7055(G7055,G873);
  not GNAME7056(G7056,G872);
  not GNAME7057(G7057,G901);
  and GNAME7058(G7058,G7230,G7123);
  and GNAME7059(G7059,G7228,G7164);
  nand GNAME7060(G7060,G7226,G7165);
  and GNAME7061(G7061,G7227,G7164);
  and GNAME7062(G7062,G7343,G7344);
  nand GNAME7063(G7063,G7224,G7166);
  and GNAME7064(G7064,G7225,G7165);
  and GNAME7065(G7065,G7345,G7346);
  nand GNAME7066(G7066,G7222,G7167);
  and GNAME7067(G7067,G7223,G7166);
  and GNAME7068(G7068,G7347,G7348);
  nand GNAME7069(G7069,G7220,G7168);
  and GNAME7070(G7070,G7221,G7167);
  and GNAME7071(G7071,G7349,G7350);
  nand GNAME7072(G7072,G7218,G7169);
  and GNAME7073(G7073,G7219,G7168);
  and GNAME7074(G7074,G7351,G7352);
  nand GNAME7075(G7075,G7216,G7170);
  and GNAME7076(G7076,G7217,G7169);
  and GNAME7077(G7077,G7353,G7354);
  nand GNAME7078(G7078,G7214,G7171);
  and GNAME7079(G7079,G7215,G7170);
  and GNAME7080(G7080,G7355,G7356);
  nand GNAME7081(G7081,G7212,G7172);
  and GNAME7082(G7082,G7213,G7171);
  and GNAME7083(G7083,G7357,G7358);
  nand GNAME7084(G7084,G7210,G7173);
  and GNAME7085(G7085,G7211,G7172);
  and GNAME7086(G7086,G7359,G7360);
  nand GNAME7087(G7087,G7208,G7174);
  and GNAME7088(G7088,G7209,G7173);
  and GNAME7089(G7089,G7361,G7362);
  nand GNAME7090(G7090,G7137,G7135);
  and GNAME7091(G7091,G7138,G7132);
  and GNAME7092(G7092,G7363,G7364);
  nand GNAME7093(G7093,G7206,G7175);
  and GNAME7094(G7094,G7207,G7174);
  and GNAME7095(G7095,G7365,G7366);
  nand GNAME7096(G7096,G7204,G7176);
  and GNAME7097(G7097,G7205,G7175);
  and GNAME7098(G7098,G7367,G7368);
  nand GNAME7099(G7099,G7202,G7177);
  and GNAME7100(G7100,G7203,G7176);
  and GNAME7101(G7101,G7369,G7370);
  nand GNAME7102(G7102,G7200,G7178);
  and GNAME7103(G7103,G7201,G7177);
  and GNAME7104(G7104,G7371,G7372);
  nand GNAME7105(G7105,G7198,G7122);
  and GNAME7106(G7106,G7199,G7178);
  and GNAME7107(G7107,G7373,G7374);
  and GNAME7108(G7108,G7196,G7182);
  nand GNAME7109(G7109,G7194,G7183);
  and GNAME7110(G7110,G7195,G7182);
  and GNAME7111(G7111,G7377,G7378);
  nand GNAME7112(G7112,G7192,G7184);
  and GNAME7113(G7113,G7193,G7183);
  and GNAME7114(G7114,G7379,G7380);
  nor GNAME7115(G7115,G7387,G7009);
  and GNAME7116(G7116,G7136,G7135);
  nand GNAME7117(G7117,G7128,G6977,G7127);
  nand GNAME7118(G7118,G7162,G7007,G7161);
  nand GNAME7119(G7119,G7134,G6979,G7133);
  nand GNAME7120(G7120,G7180,G6992,G7179);
  nand GNAME7121(G7121,G7187,G6988,G7186);
  nand GNAME7122(G7122,G7181,G920);
  nand GNAME7123(G7123,G7163,G903);
  nand GNAME7124(G7124,G7263,G927);
  nand GNAME7125(G7125,G6984,G7246,G7247);
  nand GNAME7126(G7126,G7250,G929);
  or GNAME7127(G7127,G894,G6976);
  nand GNAME7128(G7128,G6976,G894);
  nand GNAME7129(G7129,G7262,G930);
  nand GNAME7130(G7130,G7259,G931);
  nand GNAME7131(G7131,G6982,G7251,G7252);
  nand GNAME7132(G7132,G7255,G933);
  or GNAME7133(G7133,G898,G6976);
  nand GNAME7134(G7134,G6976,G898);
  nand GNAME7135(G7135,G7258,G934);
  nand GNAME7136(G7136,G6981,G7256,G7257);
  nand GNAME7137(G7137,G7136,G869);
  nand GNAME7138(G7138,G6980,G7253,G7254);
  nand GNAME7139(G7139,G7132,G7232);
  nand GNAME7140(G7140,G7133,G7134);
  nand GNAME7141(G7141,G7140,G932);
  not GNAME7142(G7142,G7039);
  nand GNAME7143(G7143,G7131,G7142);
  nand GNAME7144(G7144,G6983,G7260,G7261);
  nand GNAME7145(G7145,G7036,G7144);
  nand GNAME7146(G7146,G6978,G7248,G7249);
  nand GNAME7147(G7147,G7126,G7157);
  nand GNAME7148(G7148,G7127,G7128);
  nand GNAME7149(G7149,G7148,G928);
  not GNAME7150(G7150,G7032);
  nand GNAME7151(G7151,G7125,G7150);
  nand GNAME7152(G7152,G7266,G926);
  nand GNAME7153(G7153,G6985,G7264,G7265);
  nand GNAME7154(G7154,G7029,G7153);
  nand GNAME7155(G7155,G7269,G925);
  nand GNAME7156(G7156,G6986,G7267,G7268);
  nand GNAME7157(G7157,G7033,G7146);
  nand GNAME7158(G7158,G7117,G7149);
  nand GNAME7159(G7159,G7158,G7126,G7157);
  nand GNAME7160(G7160,G7149,G6987);
  or GNAME7161(G7161,G870,G6976);
  nand GNAME7162(G7162,G6976,G870);
  nand GNAME7163(G7163,G7162,G7161);
  nand GNAME7164(G7164,G7335,G905);
  nand GNAME7165(G7165,G7332,G906);
  nand GNAME7166(G7166,G7329,G907);
  nand GNAME7167(G7167,G7326,G908);
  nand GNAME7168(G7168,G7323,G909);
  nand GNAME7169(G7169,G7320,G910);
  nand GNAME7170(G7170,G7317,G911);
  nand GNAME7171(G7171,G7314,G912);
  nand GNAME7172(G7172,G7311,G913);
  nand GNAME7173(G7173,G7308,G914);
  nand GNAME7174(G7174,G7305,G915);
  nand GNAME7175(G7175,G7302,G916);
  nand GNAME7176(G7176,G7299,G917);
  nand GNAME7177(G7177,G7296,G918);
  nand GNAME7178(G7178,G7293,G919);
  or GNAME7179(G7179,G886,G6976);
  nand GNAME7180(G7180,G6976,G886);
  nand GNAME7181(G7181,G7180,G7179);
  nand GNAME7182(G7182,G7290,G921);
  nand GNAME7183(G7183,G7287,G922);
  nand GNAME7184(G7184,G7284,G923);
  nand GNAME7185(G7185,G6989,G7282,G7283);
  or GNAME7186(G7186,G890,G6976);
  nand GNAME7187(G7187,G6976,G890);
  nand GNAME7188(G7188,G7155,G7237);
  nand GNAME7189(G7189,G7186,G7187);
  nand GNAME7190(G7190,G7189,G924);
  not GNAME7191(G7191,G7115);
  nand GNAME7192(G7192,G7185,G7191);
  nand GNAME7193(G7193,G6990,G7285,G7286);
  nand GNAME7194(G7194,G7112,G7193);
  nand GNAME7195(G7195,G6991,G7288,G7289);
  nand GNAME7196(G7196,G7109,G7195);
  not GNAME7197(G7197,G7108);
  nand GNAME7198(G7198,G7120,G7197);
  nand GNAME7199(G7199,G6993,G7291,G7292);
  nand GNAME7200(G7200,G7105,G7199);
  nand GNAME7201(G7201,G6994,G7294,G7295);
  nand GNAME7202(G7202,G7102,G7201);
  nand GNAME7203(G7203,G6995,G7297,G7298);
  nand GNAME7204(G7204,G7099,G7203);
  nand GNAME7205(G7205,G6996,G7300,G7301);
  nand GNAME7206(G7206,G7096,G7205);
  nand GNAME7207(G7207,G6997,G7303,G7304);
  nand GNAME7208(G7208,G7093,G7207);
  nand GNAME7209(G7209,G6998,G7306,G7307);
  nand GNAME7210(G7210,G7087,G7209);
  nand GNAME7211(G7211,G6999,G7309,G7310);
  nand GNAME7212(G7212,G7084,G7211);
  nand GNAME7213(G7213,G7000,G7312,G7313);
  nand GNAME7214(G7214,G7081,G7213);
  nand GNAME7215(G7215,G7001,G7315,G7316);
  nand GNAME7216(G7216,G7078,G7215);
  nand GNAME7217(G7217,G7002,G7318,G7319);
  nand GNAME7218(G7218,G7075,G7217);
  nand GNAME7219(G7219,G7003,G7321,G7322);
  nand GNAME7220(G7220,G7072,G7219);
  nand GNAME7221(G7221,G7004,G7324,G7325);
  nand GNAME7222(G7222,G7069,G7221);
  nand GNAME7223(G7223,G7005,G7327,G7328);
  nand GNAME7224(G7224,G7066,G7223);
  nand GNAME7225(G7225,G7006,G7330,G7331);
  nand GNAME7226(G7226,G7063,G7225);
  or GNAME7227(G7227,G905,G7335);
  nand GNAME7228(G7228,G7060,G7227);
  not GNAME7229(G7229,G7059);
  nand GNAME7230(G7230,G7118,G7229);
  not GNAME7231(G7231,G7058);
  nand GNAME7232(G7232,G7090,G7138);
  nand GNAME7233(G7233,G7119,G7141);
  nand GNAME7234(G7234,G7233,G7132,G7232);
  nand GNAME7235(G7235,G7141,G7008);
  nand GNAME7236(G7236,G7121,G7190);
  nand GNAME7237(G7237,G7026,G7156);
  nand GNAME7238(G7238,G7237,G7155,G7236);
  nand GNAME7239(G7239,G7190,G7009);
  not GNAME7240(G7240,G7116);
  nand GNAME7241(G7241,G7124,G7125);
  nand GNAME7242(G7242,G7130,G7131);
  nand GNAME7243(G7243,G7118,G7123);
  nand GNAME7244(G7244,G7120,G7122);
  nand GNAME7245(G7245,G7184,G7185);
  or GNAME7246(G7246,G893,G6976);
  or GNAME7247(G7247,G869,G7018);
  or GNAME7248(G7248,G895,G6976);
  or GNAME7249(G7249,G869,G7019);
  nand GNAME7250(G7250,G7248,G7249);
  or GNAME7251(G7251,G897,G6976);
  or GNAME7252(G7252,G869,G7020);
  or GNAME7253(G7253,G899,G6976);
  or GNAME7254(G7254,G869,G7021);
  nand GNAME7255(G7255,G7253,G7254);
  or GNAME7256(G7256,G900,G6976);
  or GNAME7257(G7257,G869,G7022);
  nand GNAME7258(G7258,G7256,G7257);
  nand GNAME7259(G7259,G7251,G7252);
  or GNAME7260(G7260,G896,G6976);
  or GNAME7261(G7261,G869,G7023);
  nand GNAME7262(G7262,G7260,G7261);
  nand GNAME7263(G7263,G7246,G7247);
  or GNAME7264(G7264,G892,G6976);
  or GNAME7265(G7265,G869,G7024);
  nand GNAME7266(G7266,G7264,G7265);
  or GNAME7267(G7267,G891,G6976);
  or GNAME7268(G7268,G869,G7025);
  nand GNAME7269(G7269,G7267,G7268);
  or GNAME7270(G7270,G7027,G7026);
  nand GNAME7271(G7271,G7026,G7027);
  or GNAME7272(G7272,G7030,G7029);
  nand GNAME7273(G7273,G7029,G7030);
  nand GNAME7274(G7274,G7150,G7241);
  nand GNAME7275(G7275,G7032,G7124,G7125);
  or GNAME7276(G7276,G7034,G7033);
  nand GNAME7277(G7277,G7033,G7034);
  or GNAME7278(G7278,G7037,G7036);
  nand GNAME7279(G7279,G7036,G7037);
  nand GNAME7280(G7280,G7142,G7242);
  nand GNAME7281(G7281,G7039,G7130,G7131);
  or GNAME7282(G7282,G889,G6976);
  or GNAME7283(G7283,G869,G7040);
  nand GNAME7284(G7284,G7282,G7283);
  or GNAME7285(G7285,G888,G6976);
  or GNAME7286(G7286,G869,G7041);
  nand GNAME7287(G7287,G7285,G7286);
  or GNAME7288(G7288,G887,G6976);
  or GNAME7289(G7289,G869,G7042);
  nand GNAME7290(G7290,G7288,G7289);
  or GNAME7291(G7291,G885,G6976);
  or GNAME7292(G7292,G869,G7043);
  nand GNAME7293(G7293,G7291,G7292);
  or GNAME7294(G7294,G884,G6976);
  or GNAME7295(G7295,G869,G7044);
  nand GNAME7296(G7296,G7294,G7295);
  or GNAME7297(G7297,G883,G6976);
  or GNAME7298(G7298,G869,G7045);
  nand GNAME7299(G7299,G7297,G7298);
  or GNAME7300(G7300,G882,G6976);
  or GNAME7301(G7301,G869,G7046);
  nand GNAME7302(G7302,G7300,G7301);
  or GNAME7303(G7303,G881,G6976);
  or GNAME7304(G7304,G869,G7047);
  nand GNAME7305(G7305,G7303,G7304);
  or GNAME7306(G7306,G880,G6976);
  or GNAME7307(G7307,G869,G7048);
  nand GNAME7308(G7308,G7306,G7307);
  or GNAME7309(G7309,G879,G6976);
  or GNAME7310(G7310,G869,G7049);
  nand GNAME7311(G7311,G7309,G7310);
  or GNAME7312(G7312,G878,G6976);
  or GNAME7313(G7313,G869,G7050);
  nand GNAME7314(G7314,G7312,G7313);
  or GNAME7315(G7315,G877,G6976);
  or GNAME7316(G7316,G869,G7051);
  nand GNAME7317(G7317,G7315,G7316);
  or GNAME7318(G7318,G876,G6976);
  or GNAME7319(G7319,G869,G7052);
  nand GNAME7320(G7320,G7318,G7319);
  or GNAME7321(G7321,G875,G6976);
  or GNAME7322(G7322,G869,G7053);
  nand GNAME7323(G7323,G7321,G7322);
  or GNAME7324(G7324,G874,G6976);
  or GNAME7325(G7325,G869,G7054);
  nand GNAME7326(G7326,G7324,G7325);
  or GNAME7327(G7327,G873,G6976);
  or GNAME7328(G7328,G869,G7055);
  nand GNAME7329(G7329,G7327,G7328);
  or GNAME7330(G7330,G872,G6976);
  or GNAME7331(G7331,G869,G7056);
  nand GNAME7332(G7332,G7330,G7331);
  or GNAME7333(G7333,G871,G6976);
  nand GNAME7334(G7334,G6976,G871);
  not GNAME7335(G7335,G7010);
  or GNAME7336(G7336,G7058,G7057);
  or GNAME7337(G7337,G901,G7231);
  nand GNAME7338(G7338,G7336,G7337);
  nand GNAME7339(G7339,G7010,G7336,G7337);
  nand GNAME7340(G7340,G7335,G7338);
  nand GNAME7341(G7341,G7229,G7243);
  nand GNAME7342(G7342,G7059,G7118,G7123);
  or GNAME7343(G7343,G7061,G7060);
  nand GNAME7344(G7344,G7060,G7061);
  or GNAME7345(G7345,G7064,G7063);
  nand GNAME7346(G7346,G7063,G7064);
  or GNAME7347(G7347,G7067,G7066);
  nand GNAME7348(G7348,G7066,G7067);
  or GNAME7349(G7349,G7070,G7069);
  nand GNAME7350(G7350,G7069,G7070);
  or GNAME7351(G7351,G7073,G7072);
  nand GNAME7352(G7352,G7072,G7073);
  or GNAME7353(G7353,G7076,G7075);
  nand GNAME7354(G7354,G7075,G7076);
  or GNAME7355(G7355,G7079,G7078);
  nand GNAME7356(G7356,G7078,G7079);
  or GNAME7357(G7357,G7082,G7081);
  nand GNAME7358(G7358,G7081,G7082);
  or GNAME7359(G7359,G7085,G7084);
  nand GNAME7360(G7360,G7084,G7085);
  or GNAME7361(G7361,G7088,G7087);
  nand GNAME7362(G7362,G7087,G7088);
  or GNAME7363(G7363,G7091,G7090);
  nand GNAME7364(G7364,G7090,G7091);
  or GNAME7365(G7365,G7094,G7093);
  nand GNAME7366(G7366,G7093,G7094);
  or GNAME7367(G7367,G7097,G7096);
  nand GNAME7368(G7368,G7096,G7097);
  or GNAME7369(G7369,G7100,G7099);
  nand GNAME7370(G7370,G7099,G7100);
  or GNAME7371(G7371,G7103,G7102);
  nand GNAME7372(G7372,G7102,G7103);
  or GNAME7373(G7373,G7106,G7105);
  nand GNAME7374(G7374,G7105,G7106);
  nand GNAME7375(G7375,G7197,G7244);
  nand GNAME7376(G7376,G7108,G7120,G7122);
  or GNAME7377(G7377,G7110,G7109);
  nand GNAME7378(G7378,G7109,G7110);
  or GNAME7379(G7379,G7113,G7112);
  nand GNAME7380(G7380,G7112,G7113);
  nand GNAME7381(G7381,G7191,G7245);
  nand GNAME7382(G7382,G7115,G7184,G7185);
  or GNAME7383(G7383,G7116,G6976);
  or GNAME7384(G7384,G869,G7240);
  not GNAME7385(G7385,G7141);
  not GNAME7386(G7386,G7149);
  not GNAME7387(G7387,G7190);
  and GNAME7388(G7388,G7531,G7533);
  and GNAME7389(G7389,G7525,G7527);
  and GNAME7390(G7390,G7520,G7521);
  and GNAME7391(G7391,G7513,G7516);
  not GNAME7392(G7392,G1364);
  and GNAME7393(G7393,G1544,G1364);
  not GNAME7394(G7394,G1543);
  and GNAME7395(G7395,G7465,G7466);
  not GNAME7396(G7396,G1532);
  not GNAME7397(G7397,G1531);
  nand GNAME7398(G7398,G7468,G7469);
  and GNAME7399(G7399,G7472,G7473);
  not GNAME7400(G7400,G1529);
  and GNAME7401(G7401,G7463,G7475);
  and GNAME7402(G7402,G7477,G7478);
  not GNAME7403(G7403,G1349);
  and GNAME7404(G7404,G7480,G7481);
  not GNAME7405(G7405,G1527);
  and GNAME7406(G7406,G7483,G7484);
  not GNAME7407(G7407,G1526);
  not GNAME7408(G7408,G1525);
  not GNAME7409(G7409,G1346);
  nand GNAME7410(G7410,G7486,G7487);
  not GNAME7411(G7411,G1542);
  or GNAME7412(G7412,G7492,G7429);
  not GNAME7413(G7413,G1541);
  not GNAME7414(G7414,G1362);
  and GNAME7415(G7415,G7495,G7496);
  not GNAME7416(G7416,G1540);
  not GNAME7417(G7417,G1539);
  nand GNAME7418(G7418,G7498,G7499);
  not GNAME7419(G7419,G1538);
  and GNAME7420(G7420,G7489,G7426);
  not GNAME7421(G7421,G1357);
  and GNAME7422(G7422,G7505,G7506);
  not GNAME7423(G7423,G1356);
  not GNAME7424(G7424,G1534);
  and GNAME7425(G7425,G7508,G7509);
  nand GNAME7426(G7426,G7503,G7517);
  not GNAME7427(G7427,G1360);
  nand GNAME7428(G7428,G7522,G7501,G7502);
  and GNAME7429(G7429,G7528,G7490,G7491);
  nand GNAME7430(G7430,G7548,G7549);
  nand GNAME7431(G7431,G7554,G7555);
  nand GNAME7432(G7432,G7566,G7567);
  nand GNAME7433(G7433,G7600,G7601);
  nand GNAME7434(G7434,G7596,G7597);
  and GNAME7435(G7435,G7534,G7535);
  and GNAME7436(G7436,G7538,G7539);
  and GNAME7437(G7437,G7542,G7543);
  and GNAME7438(G7438,G7546,G7547);
  and GNAME7439(G7439,G7550,G7551);
  and GNAME7440(G7440,G7556,G7557);
  and GNAME7441(G7441,G7560,G7561);
  and GNAME7442(G7442,G7564,G7565);
  and GNAME7443(G7443,G7571,G7572);
  and GNAME7444(G7444,G7575,G7576);
  and GNAME7445(G7445,G7579,G7580);
  and GNAME7446(G7446,G7585,G7586);
  and GNAME7447(G7447,G7589,G7590);
  and GNAME7448(G7448,G7536,G7537);
  and GNAME7449(G7449,G7540,G7541);
  and GNAME7450(G7450,G7544,G7545);
  and GNAME7451(G7451,G7552,G7553);
  nand GNAME7452(G7452,G7474,G7463);
  not GNAME7453(G7453,G1352);
  and GNAME7454(G7454,G7558,G7559);
  and GNAME7455(G7455,G7562,G7563);
  not GNAME7456(G7456,G1533);
  not GNAME7457(G7457,G3200);
  and GNAME7458(G7458,G7573,G7574);
  and GNAME7459(G7459,G7577,G7578);
  and GNAME7460(G7460,G7581,G7582);
  and GNAME7461(G7461,G7587,G7588);
  and GNAME7462(G7462,G7591,G7592);
  nand GNAME7463(G7463,G1351,G1530);
  or GNAME7464(G7464,G1543,G1354);
  nand GNAME7465(G7465,G7464,G7393);
  nand GNAME7466(G7466,G1354,G1543);
  nand GNAME7467(G7467,G7396,G7395);
  nand GNAME7468(G7468,G7467,G1353);
  or GNAME7469(G7469,G7395,G7396);
  not GNAME7470(G7470,G7398);
  nand GNAME7471(G7471,G7398,G1531);
  nand GNAME7472(G7472,G7453,G7471);
  nand GNAME7473(G7473,G7397,G7470);
  or GNAME7474(G7474,G1530,G1351);
  nand GNAME7475(G7475,G7474,G7399);
  nand GNAME7476(G7476,G1350,G1529);
  nand GNAME7477(G7477,G7476,G7401);
  or GNAME7478(G7478,G1350,G1529);
  or GNAME7479(G7479,G1349,G1528);
  nand GNAME7480(G7480,G7479,G7402);
  nand GNAME7481(G7481,G1528,G1349);
  nand GNAME7482(G7482,G7405,G7404);
  nand GNAME7483(G7483,G7482,G1348);
  or GNAME7484(G7484,G7404,G7405);
  nand GNAME7485(G7485,G7407,G7406);
  nand GNAME7486(G7486,G7485,G1347);
  or GNAME7487(G7487,G7406,G7407);
  not GNAME7488(G7488,G7410);
  nand GNAME7489(G7489,G1358,G1537);
  nand GNAME7490(G7490,G7408,G7530);
  or GNAME7491(G7491,G1363,G1542);
  and GNAME7492(G7492,G1363,G1542);
  not GNAME7493(G7493,G7412);
  nand GNAME7494(G7494,G7414,G7493);
  nand GNAME7495(G7495,G7494,G1541);
  nand GNAME7496(G7496,G7412,G1362);
  nand GNAME7497(G7497,G7416,G7415);
  nand GNAME7498(G7498,G7497,G1361);
  or GNAME7499(G7499,G7415,G7416);
  not GNAME7500(G7500,G7418);
  nand GNAME7501(G7501,G7427,G7524);
  or GNAME7502(G7502,G1359,G1538);
  nand GNAME7503(G7503,G7428,G7519);
  nand GNAME7504(G7504,G7421,G7420);
  nand GNAME7505(G7505,G7504,G1536);
  or GNAME7506(G7506,G7420,G7421);
  nand GNAME7507(G7507,G7423,G7422);
  nand GNAME7508(G7508,G7507,G1535);
  or GNAME7509(G7509,G7422,G7423);
  nor GNAME7510(G7510,G1534,G1355);
  or GNAME7511(G7511,G7425,G7510);
  nand GNAME7512(G7512,G1355,G1534);
  nand GNAME7513(G7513,G7568,G7569,G7511,G7512);
  nand GNAME7514(G7514,G7512,G7425);
  or GNAME7515(G7515,G1355,G1534);
  nand GNAME7516(G7516,G7570,G7514,G7515);
  or GNAME7517(G7517,G1537,G1358);
  nand GNAME7518(G7518,G7489,G7517);
  nand GNAME7519(G7519,G1359,G1538);
  nand GNAME7520(G7520,G7519,G7428,G7518);
  nand GNAME7521(G7521,G7489,G7602);
  nand GNAME7522(G7522,G7417,G7500);
  nand GNAME7523(G7523,G7522,G1360);
  nand GNAME7524(G7524,G7418,G1539);
  nand GNAME7525(G7525,G7583,G7584,G7523,G7524);
  and GNAME7526(G7526,G1359,G1538);
  or GNAME7527(G7527,G7526,G7428);
  nand GNAME7528(G7528,G7409,G7488);
  nand GNAME7529(G7529,G7528,G1525);
  nand GNAME7530(G7530,G7410,G1346);
  nand GNAME7531(G7531,G7598,G7599,G7529,G7530);
  nand GNAME7532(G7532,G1363,G1542);
  nand GNAME7533(G7533,G7532,G7429);
  nand GNAME7534(G7534,G7409,G1525);
  nand GNAME7535(G7535,G7408,G1346);
  nand GNAME7536(G7536,G7488,G7435);
  or GNAME7537(G7537,G7488,G7435);
  nand GNAME7538(G7538,G7407,G1347);
  or GNAME7539(G7539,G1347,G7407);
  nand GNAME7540(G7540,G7406,G7436);
  or GNAME7541(G7541,G7406,G7436);
  nand GNAME7542(G7542,G7405,G1348);
  or GNAME7543(G7543,G1348,G7405);
  nand GNAME7544(G7544,G7404,G7437);
  or GNAME7545(G7545,G7404,G7437);
  or GNAME7546(G7546,G1528,G7403);
  nand GNAME7547(G7547,G7403,G1528);
  nand GNAME7548(G7548,G7402,G7438);
  or GNAME7549(G7549,G7402,G7438);
  nand GNAME7550(G7550,G7400,G7401);
  or GNAME7551(G7551,G7401,G7400);
  nand GNAME7552(G7552,G1350,G7439);
  or GNAME7553(G7553,G1350,G7439);
  nand GNAME7554(G7554,G7452,G7399);
  or GNAME7555(G7555,G7399,G7452);
  nand GNAME7556(G7556,G7397,G1352);
  nand GNAME7557(G7557,G7453,G1531);
  nand GNAME7558(G7558,G7470,G7440);
  or GNAME7559(G7559,G7470,G7440);
  nand GNAME7560(G7560,G7396,G1353);
  or GNAME7561(G7561,G1353,G7396);
  nand GNAME7562(G7562,G7395,G7441);
  or GNAME7563(G7563,G7395,G7441);
  or GNAME7564(G7564,G1354,G7394);
  nand GNAME7565(G7565,G7394,G1354);
  nand GNAME7566(G7566,G7393,G7442);
  or GNAME7567(G7567,G7393,G7442);
  nand GNAME7568(G7568,G7457,G1533);
  nand GNAME7569(G7569,G7456,G3200);
  nand GNAME7570(G7570,G7568,G7569);
  or GNAME7571(G7571,G1355,G7424);
  nand GNAME7572(G7572,G7424,G1355);
  nand GNAME7573(G7573,G7425,G7443);
  or GNAME7574(G7574,G7425,G7443);
  nand GNAME7575(G7575,G7423,G1535);
  or GNAME7576(G7576,G1535,G7423);
  nand GNAME7577(G7577,G7422,G7444);
  or GNAME7578(G7578,G7422,G7444);
  nand GNAME7579(G7579,G7421,G1536);
  or GNAME7580(G7580,G1536,G7421);
  nand GNAME7581(G7581,G7420,G7445);
  or GNAME7582(G7582,G7420,G7445);
  or GNAME7583(G7583,G1359,G7419);
  nand GNAME7584(G7584,G7419,G1359);
  nand GNAME7585(G7585,G7417,G1360);
  nand GNAME7586(G7586,G7427,G1539);
  nand GNAME7587(G7587,G7500,G7446);
  or GNAME7588(G7588,G7500,G7446);
  nand GNAME7589(G7589,G7416,G1361);
  or GNAME7590(G7590,G1361,G7416);
  nand GNAME7591(G7591,G7415,G7447);
  or GNAME7592(G7592,G7415,G7447);
  nand GNAME7593(G7593,G7414,G1541);
  nand GNAME7594(G7594,G7413,G1362);
  nand GNAME7595(G7595,G7593,G7594);
  nand GNAME7596(G7596,G7412,G7593,G7594);
  nand GNAME7597(G7597,G7493,G7595);
  or GNAME7598(G7598,G1363,G7411);
  nand GNAME7599(G7599,G7411,G1363);
  or GNAME7600(G7600,G1544,G7392);
  nand GNAME7601(G7601,G7392,G1544);
  not GNAME7602(G7602,G7426);
  nand GNAME7603(G7603,G7728,G7727);
  not GNAME7604(G7604,G1389);
  not GNAME7605(G7605,G1421);
  not GNAME7606(G7606,G1375);
  not GNAME7607(G7607,G1416);
  not GNAME7608(G7608,G1373);
  not GNAME7609(G7609,G1423);
  not GNAME7610(G7610,G1371);
  not GNAME7611(G7611,G1410);
  not GNAME7612(G7612,G1369);
  not GNAME7613(G7613,G1407);
  not GNAME7614(G7614,G1398);
  not GNAME7615(G7615,G1412);
  not GNAME7616(G7616,G1396);
  not GNAME7617(G7617,G1406);
  not GNAME7618(G7618,G1394);
  not GNAME7619(G7619,G1413);
  not GNAME7620(G7620,G1392);
  not GNAME7621(G7621,G1422);
  not GNAME7622(G7622,G1390);
  not GNAME7623(G7623,G1249);
  not GNAME7624(G7624,G1387);
  not GNAME7625(G7625,G1250);
  not GNAME7626(G7626,G1385);
  not GNAME7627(G7627,G1248);
  not GNAME7628(G7628,G1383);
  not GNAME7629(G7629,G1251);
  not GNAME7630(G7630,G1381);
  not GNAME7631(G7631,G1245);
  not GNAME7632(G7632,G1379);
  not GNAME7633(G7633,G1256);
  not GNAME7634(G7634,G1255);
  not GNAME7635(G7635,G1400);
  or GNAME7636(G7636,G1411,G7604);
  nand GNAME7637(G7637,G1418,G7635,G7636);
  or GNAME7638(G7638,G1378,G7605);
  nand GNAME7639(G7639,G7604,G1411);
  nand GNAME7640(G7640,G7639,G7637,G7638);
  or GNAME7641(G7641,G1408,G7606);
  nand GNAME7642(G7642,G7605,G1378);
  nand GNAME7643(G7643,G7642,G7640,G7641);
  or GNAME7644(G7644,G1374,G7607);
  nand GNAME7645(G7645,G7606,G1408);
  nand GNAME7646(G7646,G7645,G7643,G7644);
  or GNAME7647(G7647,G1414,G7608);
  nand GNAME7648(G7648,G7607,G1374);
  nand GNAME7649(G7649,G7648,G7646,G7647);
  or GNAME7650(G7650,G1372,G7609);
  nand GNAME7651(G7651,G7608,G1414);
  nand GNAME7652(G7652,G7651,G7649,G7650);
  or GNAME7653(G7653,G1405,G7610);
  nand GNAME7654(G7654,G7609,G1372);
  nand GNAME7655(G7655,G7654,G7652,G7653);
  or GNAME7656(G7656,G1370,G7611);
  nand GNAME7657(G7657,G7610,G1405);
  nand GNAME7658(G7658,G7657,G7655,G7656);
  or GNAME7659(G7659,G1417,G7612);
  nand GNAME7660(G7660,G7611,G1370);
  nand GNAME7661(G7661,G7660,G7658,G7659);
  or GNAME7662(G7662,G1399,G7613);
  nand GNAME7663(G7663,G7612,G1417);
  nand GNAME7664(G7664,G7663,G7661,G7662);
  or GNAME7665(G7665,G1420,G7614);
  nand GNAME7666(G7666,G7613,G1399);
  nand GNAME7667(G7667,G7666,G7664,G7665);
  or GNAME7668(G7668,G1397,G7615);
  nand GNAME7669(G7669,G7614,G1420);
  nand GNAME7670(G7670,G7669,G7667,G7668);
  or GNAME7671(G7671,G1419,G7616);
  nand GNAME7672(G7672,G7615,G1397);
  nand GNAME7673(G7673,G7672,G7670,G7671);
  or GNAME7674(G7674,G1395,G7617);
  nand GNAME7675(G7675,G7616,G1419);
  nand GNAME7676(G7676,G7675,G7673,G7674);
  or GNAME7677(G7677,G1424,G7618);
  nand GNAME7678(G7678,G7617,G1395);
  nand GNAME7679(G7679,G7678,G7676,G7677);
  or GNAME7680(G7680,G1393,G7619);
  nand GNAME7681(G7681,G7618,G1424);
  nand GNAME7682(G7682,G7681,G7679,G7680);
  or GNAME7683(G7683,G1415,G7620);
  nand GNAME7684(G7684,G7619,G1393);
  nand GNAME7685(G7685,G7684,G7682,G7683);
  or GNAME7686(G7686,G1391,G7621);
  nand GNAME7687(G7687,G7620,G1415);
  nand GNAME7688(G7688,G7687,G7685,G7686);
  or GNAME7689(G7689,G1409,G7622);
  nand GNAME7690(G7690,G7621,G1391);
  nand GNAME7691(G7691,G7690,G7688,G7689);
  or GNAME7692(G7692,G1388,G7623);
  nand GNAME7693(G7693,G7622,G1409);
  nand GNAME7694(G7694,G7693,G7691,G7692);
  or GNAME7695(G7695,G1246,G7624);
  nand GNAME7696(G7696,G7623,G1388);
  nand GNAME7697(G7697,G7696,G7694,G7695);
  or GNAME7698(G7698,G1386,G7625);
  nand GNAME7699(G7699,G7624,G1246);
  nand GNAME7700(G7700,G7699,G7697,G7698);
  or GNAME7701(G7701,G1244,G7626);
  nand GNAME7702(G7702,G7625,G1386);
  nand GNAME7703(G7703,G7702,G7700,G7701);
  or GNAME7704(G7704,G1384,G7627);
  nand GNAME7705(G7705,G7626,G1244);
  nand GNAME7706(G7706,G7705,G7703,G7704);
  or GNAME7707(G7707,G1247,G7628);
  nand GNAME7708(G7708,G7627,G1384);
  nand GNAME7709(G7709,G7708,G7706,G7707);
  or GNAME7710(G7710,G1382,G7629);
  nand GNAME7711(G7711,G7628,G1247);
  nand GNAME7712(G7712,G7711,G7709,G7710);
  or GNAME7713(G7713,G1243,G7630);
  nand GNAME7714(G7714,G7629,G1382);
  nand GNAME7715(G7715,G7714,G7712,G7713);
  or GNAME7716(G7716,G1380,G7631);
  nand GNAME7717(G7717,G7630,G1243);
  nand GNAME7718(G7718,G7717,G7715,G7716);
  or GNAME7719(G7719,G1253,G7632);
  nand GNAME7720(G7720,G7631,G1380);
  nand GNAME7721(G7721,G7720,G7718,G7719);
  or GNAME7722(G7722,G1377,G7633);
  nand GNAME7723(G7723,G7632,G1253);
  nand GNAME7724(G7724,G7723,G7721,G7722);
  or GNAME7725(G7725,G1376,G7634);
  nand GNAME7726(G7726,G7633,G1377);
  nand GNAME7727(G7727,G7726,G7724,G7725);
  nand GNAME7728(G7728,G7634,G1376);
  nand GNAME7729(G7729,G7855,G7858,G7859);
  nor GNAME7730(G7730,G1000,G7731);
  not GNAME7731(G7731,G936);
  not GNAME7732(G7732,G999);
  not GNAME7733(G7733,G966);
  not GNAME7734(G7734,G997);
  not GNAME7735(G7735,G964);
  not GNAME7736(G7736,G995);
  not GNAME7737(G7737,G962);
  not GNAME7738(G7738,G993);
  not GNAME7739(G7739,G960);
  not GNAME7740(G7740,G991);
  not GNAME7741(G7741,G958);
  not GNAME7742(G7742,G989);
  not GNAME7743(G7743,G956);
  not GNAME7744(G7744,G987);
  not GNAME7745(G7745,G954);
  not GNAME7746(G7746,G985);
  not GNAME7747(G7747,G952);
  not GNAME7748(G7748,G983);
  not GNAME7749(G7749,G950);
  not GNAME7750(G7750,G981);
  not GNAME7751(G7751,G948);
  not GNAME7752(G7752,G979);
  not GNAME7753(G7753,G946);
  not GNAME7754(G7754,G977);
  not GNAME7755(G7755,G944);
  not GNAME7756(G7756,G975);
  not GNAME7757(G7757,G942);
  not GNAME7758(G7758,G973);
  not GNAME7759(G7759,G940);
  not GNAME7760(G7760,G971);
  not GNAME7761(G7761,G970);
  not GNAME7762(G7762,G937);
  or GNAME7763(G7763,G7730,G968);
  or GNAME7764(G7764,G967,G7732);
  nand GNAME7765(G7765,G7731,G1000);
  nand GNAME7766(G7766,G7765,G7763,G7764);
  or GNAME7767(G7767,G998,G7733);
  nand GNAME7768(G7768,G7732,G967);
  nand GNAME7769(G7769,G7768,G7766,G7767);
  or GNAME7770(G7770,G965,G7734);
  nand GNAME7771(G7771,G7733,G998);
  nand GNAME7772(G7772,G7771,G7769,G7770);
  or GNAME7773(G7773,G996,G7735);
  nand GNAME7774(G7774,G7734,G965);
  nand GNAME7775(G7775,G7774,G7772,G7773);
  or GNAME7776(G7776,G963,G7736);
  nand GNAME7777(G7777,G7735,G996);
  nand GNAME7778(G7778,G7777,G7775,G7776);
  or GNAME7779(G7779,G994,G7737);
  nand GNAME7780(G7780,G7736,G963);
  nand GNAME7781(G7781,G7780,G7778,G7779);
  or GNAME7782(G7782,G961,G7738);
  nand GNAME7783(G7783,G7737,G994);
  nand GNAME7784(G7784,G7783,G7781,G7782);
  or GNAME7785(G7785,G992,G7739);
  nand GNAME7786(G7786,G7738,G961);
  nand GNAME7787(G7787,G7786,G7784,G7785);
  or GNAME7788(G7788,G959,G7740);
  nand GNAME7789(G7789,G7739,G992);
  nand GNAME7790(G7790,G7789,G7787,G7788);
  or GNAME7791(G7791,G990,G7741);
  nand GNAME7792(G7792,G7740,G959);
  nand GNAME7793(G7793,G7792,G7790,G7791);
  or GNAME7794(G7794,G957,G7742);
  nand GNAME7795(G7795,G7741,G990);
  nand GNAME7796(G7796,G7795,G7793,G7794);
  or GNAME7797(G7797,G988,G7743);
  nand GNAME7798(G7798,G7742,G957);
  nand GNAME7799(G7799,G7798,G7796,G7797);
  or GNAME7800(G7800,G955,G7744);
  nand GNAME7801(G7801,G7743,G988);
  nand GNAME7802(G7802,G7801,G7799,G7800);
  or GNAME7803(G7803,G986,G7745);
  nand GNAME7804(G7804,G7744,G955);
  nand GNAME7805(G7805,G7804,G7802,G7803);
  or GNAME7806(G7806,G953,G7746);
  nand GNAME7807(G7807,G7745,G986);
  nand GNAME7808(G7808,G7807,G7805,G7806);
  or GNAME7809(G7809,G984,G7747);
  nand GNAME7810(G7810,G7746,G953);
  nand GNAME7811(G7811,G7810,G7808,G7809);
  or GNAME7812(G7812,G951,G7748);
  nand GNAME7813(G7813,G7747,G984);
  nand GNAME7814(G7814,G7813,G7811,G7812);
  or GNAME7815(G7815,G982,G7749);
  nand GNAME7816(G7816,G7748,G951);
  nand GNAME7817(G7817,G7816,G7814,G7815);
  or GNAME7818(G7818,G949,G7750);
  nand GNAME7819(G7819,G7749,G982);
  nand GNAME7820(G7820,G7819,G7817,G7818);
  or GNAME7821(G7821,G980,G7751);
  nand GNAME7822(G7822,G7750,G949);
  nand GNAME7823(G7823,G7822,G7820,G7821);
  or GNAME7824(G7824,G947,G7752);
  nand GNAME7825(G7825,G7751,G980);
  nand GNAME7826(G7826,G7825,G7823,G7824);
  or GNAME7827(G7827,G978,G7753);
  nand GNAME7828(G7828,G7752,G947);
  nand GNAME7829(G7829,G7828,G7826,G7827);
  or GNAME7830(G7830,G945,G7754);
  nand GNAME7831(G7831,G7753,G978);
  nand GNAME7832(G7832,G7831,G7829,G7830);
  or GNAME7833(G7833,G976,G7755);
  nand GNAME7834(G7834,G7754,G945);
  nand GNAME7835(G7835,G7834,G7832,G7833);
  or GNAME7836(G7836,G943,G7756);
  nand GNAME7837(G7837,G7755,G976);
  nand GNAME7838(G7838,G7837,G7835,G7836);
  or GNAME7839(G7839,G974,G7757);
  nand GNAME7840(G7840,G7756,G943);
  nand GNAME7841(G7841,G7840,G7838,G7839);
  or GNAME7842(G7842,G941,G7758);
  nand GNAME7843(G7843,G7757,G974);
  nand GNAME7844(G7844,G7843,G7841,G7842);
  or GNAME7845(G7845,G972,G7759);
  nand GNAME7846(G7846,G7758,G941);
  nand GNAME7847(G7847,G7846,G7844,G7845);
  or GNAME7848(G7848,G939,G7760);
  nand GNAME7849(G7849,G7759,G972);
  nand GNAME7850(G7850,G7849,G7847,G7848);
  nand GNAME7851(G7851,G7761,G938);
  nand GNAME7852(G7852,G7760,G939);
  nand GNAME7853(G7853,G7852,G7850,G7851);
  or GNAME7854(G7854,G938,G7761);
  nand GNAME7855(G7855,G7856,G7857,G7853,G7854);
  or GNAME7856(G7856,G969,G7762);
  nand GNAME7857(G7857,G7762,G969);
  or GNAME7858(G7858,G969,G935,G7762);
  nand GNAME7859(G7859,G969,G7762,G935);
  and GNAME7860(G7860,G7879,G7925);
  and GNAME7861(G7861,G7881,G7922);
  and GNAME7862(G7862,G7883,G7920);
  and GNAME7863(G7863,G7885,G7918);
  and GNAME7864(G7864,G7887,G7916);
  and GNAME7865(G7865,G7889,G7914);
  and GNAME7866(G7866,G7875,G7913);
  and GNAME7867(G7867,G7877,G7910);
  and GNAME7868(G7868,G7878,G7909);
  and GNAME7869(G7869,G7876,G7911);
  and GNAME7870(G7870,G7888,G7915);
  and GNAME7871(G7871,G7886,G7917);
  and GNAME7872(G7872,G7884,G7919);
  and GNAME7873(G7873,G7882,G7921);
  and GNAME7874(G7874,G7880,G7923);
  or GNAME7875(G7875,G22557,G22558,G22556);
  or GNAME7876(G7876,G7875,G22559,G22560);
  or GNAME7877(G7877,G7876,G22562,G22561);
  or GNAME7878(G7878,G7877,G22563,G22564);
  or GNAME7879(G7879,G7878,G22565,G22566);
  or GNAME7880(G7880,G7879,G22567,G22568);
  or GNAME7881(G7881,G7880,G22570,G22569);
  or GNAME7882(G7882,G7881,G22571,G22572);
  or GNAME7883(G7883,G7882,G22574,G22573);
  or GNAME7884(G7884,G7883,G22575,G22576);
  or GNAME7885(G7885,G7884,G22578,G22577);
  or GNAME7886(G7886,G7885,G22579,G22580);
  or GNAME7887(G7887,G7886,G22582,G22581);
  or GNAME7888(G7888,G7887,G22583,G22584);
  or GNAME7889(G7889,G22585,G7888);
  nand GNAME7890(G7890,G7945,G7946);
  not GNAME7891(G7891,G22565);
  and GNAME7892(G7892,G7926,G7924);
  and GNAME7893(G7893,G7927,G7928);
  and GNAME7894(G7894,G7929,G7930);
  and GNAME7895(G7895,G7931,G7932);
  and GNAME7896(G7896,G7933,G7934);
  and GNAME7897(G7897,G7935,G7936);
  and GNAME7898(G7898,G7937,G7938);
  and GNAME7899(G7899,G7939,G7940);
  and GNAME7900(G7900,G7941,G7942);
  and GNAME7901(G7901,G7943,G7944);
  not GNAME7902(G7902,G22556);
  and GNAME7903(G7903,G7947,G7948);
  and GNAME7904(G7904,G7949,G7950);
  and GNAME7905(G7905,G7951,G7952);
  and GNAME7906(G7906,G7953,G7954);
  and GNAME7907(G7907,G7955,G7956);
  not GNAME7908(G7908,G7878);
  nand GNAME7909(G7909,G7928,G22564);
  nand GNAME7910(G7910,G7930,G22562);
  nand GNAME7911(G7911,G7932,G22560);
  or GNAME7912(G7912,G22557,G22556);
  nand GNAME7913(G7913,G7912,G22558);
  nand GNAME7914(G7914,G7888,G22585);
  nand GNAME7915(G7915,G7938,G22584);
  nand GNAME7916(G7916,G7940,G22582);
  nand GNAME7917(G7917,G7942,G22580);
  nand GNAME7918(G7918,G7944,G22578);
  nand GNAME7919(G7919,G7948,G22576);
  nand GNAME7920(G7920,G7950,G22574);
  nand GNAME7921(G7921,G7952,G22572);
  nand GNAME7922(G7922,G7954,G22570);
  nand GNAME7923(G7923,G7956,G22568);
  nand GNAME7924(G7924,G7891,G7908);
  nand GNAME7925(G7925,G7924,G22566);
  nand GNAME7926(G7926,G7878,G22565);
  nand GNAME7927(G7927,G7877,G22563);
  or GNAME7928(G7928,G22563,G7877);
  nand GNAME7929(G7929,G7876,G22561);
  or GNAME7930(G7930,G22561,G7876);
  nand GNAME7931(G7931,G7875,G22559);
  or GNAME7932(G7932,G22559,G7875);
  nand GNAME7933(G7933,G7936,G22587);
  or GNAME7934(G7934,G22587,G7936);
  nand GNAME7935(G7935,G7889,G22586);
  or GNAME7936(G7936,G22586,G7889);
  nand GNAME7937(G7937,G7887,G22583);
  or GNAME7938(G7938,G22583,G7887);
  nand GNAME7939(G7939,G7886,G22581);
  or GNAME7940(G7940,G22581,G7886);
  nand GNAME7941(G7941,G7885,G22579);
  or GNAME7942(G7942,G22579,G7885);
  nand GNAME7943(G7943,G7884,G22577);
  or GNAME7944(G7944,G22577,G7884);
  or GNAME7945(G7945,G22557,G7902);
  nand GNAME7946(G7946,G7902,G22557);
  nand GNAME7947(G7947,G7883,G22575);
  or GNAME7948(G7948,G22575,G7883);
  nand GNAME7949(G7949,G7882,G22573);
  or GNAME7950(G7950,G22573,G7882);
  nand GNAME7951(G7951,G7881,G22571);
  or GNAME7952(G7952,G22571,G7881);
  nand GNAME7953(G7953,G7880,G22569);
  or GNAME7954(G7954,G22569,G7880);
  nand GNAME7955(G7955,G7879,G22567);
  or GNAME7956(G7956,G22567,G7879);
  and GNAME7957(G7957,G7958,G904);
  not GNAME7958(G7958,G902);
  not GNAME7959(G7959,G22792);
  and GNAME7960(G7960,G22796,G22790,G7988);
  not GNAME7961(G7961,G22783);
  nand GNAME7962(G7962,G22783,G22792,G22780);
  and GNAME7963(G7963,G22771,G8081);
  not GNAME7964(G7964,G22797);
  and GNAME7965(G7965,G7963,G22797);
  not GNAME7966(G7966,G22789);
  nand GNAME7967(G7967,G7965,G22789);
  and GNAME7968(G7968,G22779,G8082);
  not GNAME7969(G7969,G22793);
  not GNAME7970(G7970,G22774);
  nand GNAME7971(G7971,G22774,G7968,G22793);
  not GNAME7972(G7972,G22776);
  nand GNAME7973(G7973,G22776,G22786,G8025);
  not GNAME7974(G7974,G22769);
  nand GNAME7975(G7975,G22769,G22795,G8026);
  not GNAME7976(G7976,G22782);
  nand GNAME7977(G7977,G22782,G22784,G8027);
  not GNAME7978(G7978,G22791);
  nand GNAME7979(G7979,G22791,G22772,G8028);
  not GNAME7980(G7980,G22787);
  nand GNAME7981(G7981,G22787,G22777,G8029);
  not GNAME7982(G7982,G22794);
  nand GNAME7983(G7983,G22794,G22775,G8030);
  and GNAME7984(G7984,G22781,G8083);
  not GNAME7985(G7985,G22770);
  not GNAME7986(G7986,G22785);
  not GNAME7987(G7987,G22790);
  and GNAME7988(G7988,G22785,G7984,G22770);
  not GNAME7989(G7989,G22796);
  nand GNAME7990(G7990,G8031,G8032);
  nand GNAME7991(G7991,G8033,G8034);
  nand GNAME7992(G7992,G8035,G8036);
  nand GNAME7993(G7993,G8037,G8038);
  nand GNAME7994(G7994,G8039,G8040);
  nand GNAME7995(G7995,G8041,G8042);
  nand GNAME7996(G7996,G8043,G8044);
  nand GNAME7997(G7997,G8045,G8046);
  nand GNAME7998(G7998,G8047,G8048);
  nand GNAME7999(G7999,G8049,G8050);
  nand GNAME8000(G8000,G8051,G8052);
  nand GNAME8001(G8001,G8053,G8054);
  nand GNAME8002(G8002,G8055,G8056);
  nand GNAME8003(G8003,G8057,G8058);
  nand GNAME8004(G8004,G8059,G8060);
  nand GNAME8005(G8005,G8061,G8062);
  nand GNAME8006(G8006,G8063,G8064);
  nand GNAME8007(G8007,G8065,G8066);
  nand GNAME8008(G8008,G8067,G8068);
  nand GNAME8009(G8009,G8069,G8070);
  nand GNAME8010(G8010,G8071,G8072);
  nand GNAME8011(G8011,G8073,G8074);
  nand GNAME8012(G8012,G8075,G8076);
  nand GNAME8013(G8013,G8077,G8078);
  nand GNAME8014(G8014,G8079,G8080);
  and GNAME8015(G8015,G22792,G22780);
  and GNAME8016(G8016,G7988,G22796);
  and GNAME8017(G8017,G7984,G22785);
  and GNAME8018(G8018,G22775,G8030);
  and GNAME8019(G8019,G22777,G8029);
  and GNAME8020(G8020,G22772,G8028);
  and GNAME8021(G8021,G22784,G8027);
  and GNAME8022(G8022,G22795,G8026);
  and GNAME8023(G8023,G22786,G8025);
  and GNAME8024(G8024,G7968,G22793);
  not GNAME8025(G8025,G7971);
  not GNAME8026(G8026,G7973);
  not GNAME8027(G8027,G7975);
  not GNAME8028(G8028,G7977);
  not GNAME8029(G8029,G7979);
  not GNAME8030(G8030,G7981);
  nand GNAME8031(G8031,G7967,G22779);
  or GNAME8032(G8032,G22779,G7967);
  or GNAME8033(G8033,G7965,G7966);
  nand GNAME8034(G8034,G7966,G7965);
  or GNAME8035(G8035,G7963,G7964);
  nand GNAME8036(G8036,G7964,G7963);
  or GNAME8037(G8037,G22771,G7962);
  nand GNAME8038(G8038,G7962,G22771);
  or GNAME8039(G8039,G8015,G7961);
  nand GNAME8040(G8040,G7961,G8015);
  or GNAME8041(G8041,G7959,G22780);
  nand GNAME8042(G8042,G7959,G22780);
  or GNAME8043(G8043,G8016,G7987);
  nand GNAME8044(G8044,G7987,G8016);
  or GNAME8045(G8045,G7988,G7989);
  nand GNAME8046(G8046,G7989,G7988);
  or GNAME8047(G8047,G8017,G7985);
  nand GNAME8048(G8048,G7985,G8017);
  or GNAME8049(G8049,G7984,G7986);
  nand GNAME8050(G8050,G7986,G7984);
  or GNAME8051(G8051,G22781,G7983);
  nand GNAME8052(G8052,G7983,G22781);
  or GNAME8053(G8053,G8018,G7982);
  nand GNAME8054(G8054,G7982,G8018);
  or GNAME8055(G8055,G22775,G7981);
  nand GNAME8056(G8056,G7981,G22775);
  or GNAME8057(G8057,G8019,G7980);
  nand GNAME8058(G8058,G7980,G8019);
  or GNAME8059(G8059,G22777,G7979);
  nand GNAME8060(G8060,G7979,G22777);
  or GNAME8061(G8061,G8020,G7978);
  nand GNAME8062(G8062,G7978,G8020);
  or GNAME8063(G8063,G22772,G7977);
  nand GNAME8064(G8064,G7977,G22772);
  or GNAME8065(G8065,G8021,G7976);
  nand GNAME8066(G8066,G7976,G8021);
  or GNAME8067(G8067,G22784,G7975);
  nand GNAME8068(G8068,G7975,G22784);
  or GNAME8069(G8069,G8022,G7974);
  nand GNAME8070(G8070,G7974,G8022);
  or GNAME8071(G8071,G22795,G7973);
  nand GNAME8072(G8072,G7973,G22795);
  or GNAME8073(G8073,G8023,G7972);
  nand GNAME8074(G8074,G7972,G8023);
  or GNAME8075(G8075,G22786,G7971);
  nand GNAME8076(G8076,G7971,G22786);
  or GNAME8077(G8077,G8024,G7970);
  nand GNAME8078(G8078,G7970,G8024);
  or GNAME8079(G8079,G7968,G7969);
  nand GNAME8080(G8080,G7969,G7968);
  not GNAME8081(G8081,G7962);
  not GNAME8082(G8082,G7967);
  not GNAME8083(G8083,G7983);
  nand GNAME8084(G8084,G8330,G8326);
  nand GNAME8085(G8085,G8331,G8208);
  not GNAME8086(G8086,G1033);
  not GNAME8087(G8087,G1032);
  nand GNAME8088(G8088,G8210,G8211);
  not GNAME8089(G8089,G1031);
  not GNAME8090(G8090,G1063);
  nand GNAME8091(G8091,G8214,G8215);
  not GNAME8092(G8092,G1030);
  not GNAME8093(G8093,G1062);
  nand GNAME8094(G8094,G8218,G8219);
  not GNAME8095(G8095,G1029);
  not GNAME8096(G8096,G1061);
  nand GNAME8097(G8097,G8222,G8223);
  not GNAME8098(G8098,G1028);
  not GNAME8099(G8099,G1060);
  nand GNAME8100(G8100,G8226,G8227);
  not GNAME8101(G8101,G1027);
  not GNAME8102(G8102,G1059);
  nand GNAME8103(G8103,G8230,G8231);
  not GNAME8104(G8104,G1026);
  not GNAME8105(G8105,G1058);
  nand GNAME8106(G8106,G8234,G8235);
  not GNAME8107(G8107,G1025);
  not GNAME8108(G8108,G1057);
  not GNAME8109(G8109,G1056);
  not GNAME8110(G8110,G1024);
  nand GNAME8111(G8111,G8238,G8239);
  nand GNAME8112(G8112,G8242,G8243);
  not GNAME8113(G8113,G1023);
  not GNAME8114(G8114,G1055);
  nand GNAME8115(G8115,G8246,G8247);
  not GNAME8116(G8116,G1022);
  not GNAME8117(G8117,G1054);
  nand GNAME8118(G8118,G8250,G8251);
  not GNAME8119(G8119,G1021);
  not GNAME8120(G8120,G1053);
  nand GNAME8121(G8121,G8254,G8255);
  not GNAME8122(G8122,G1020);
  not GNAME8123(G8123,G1052);
  nand GNAME8124(G8124,G8258,G8259);
  not GNAME8125(G8125,G1019);
  not GNAME8126(G8126,G1051);
  nand GNAME8127(G8127,G8262,G8263);
  not GNAME8128(G8128,G1018);
  not GNAME8129(G8129,G1050);
  nand GNAME8130(G8130,G8266,G8267);
  not GNAME8131(G8131,G1017);
  not GNAME8132(G8132,G1049);
  nand GNAME8133(G8133,G8270,G8271);
  not GNAME8134(G8134,G1016);
  not GNAME8135(G8135,G1048);
  nand GNAME8136(G8136,G8274,G8275);
  not GNAME8137(G8137,G1015);
  not GNAME8138(G8138,G1047);
  nand GNAME8139(G8139,G8278,G8279);
  not GNAME8140(G8140,G1014);
  not GNAME8141(G8141,G1046);
  nand GNAME8142(G8142,G8282,G8283);
  not GNAME8143(G8143,G1013);
  not GNAME8144(G8144,G1045);
  nand GNAME8145(G8145,G8286,G8287);
  not GNAME8146(G8146,G1012);
  not GNAME8147(G8147,G1044);
  nand GNAME8148(G8148,G8290,G8291);
  not GNAME8149(G8149,G1011);
  not GNAME8150(G8150,G1043);
  nand GNAME8151(G8151,G8294,G8295);
  not GNAME8152(G8152,G1010);
  not GNAME8153(G8153,G1042);
  nand GNAME8154(G8154,G8298,G8299);
  not GNAME8155(G8155,G1009);
  not GNAME8156(G8156,G1041);
  nand GNAME8157(G8157,G8302,G8303);
  not GNAME8158(G8158,G1008);
  not GNAME8159(G8159,G1040);
  nand GNAME8160(G8160,G8306,G8307);
  not GNAME8161(G8161,G1007);
  not GNAME8162(G8162,G1039);
  nand GNAME8163(G8163,G8310,G8311);
  not GNAME8164(G8164,G1006);
  not GNAME8165(G8165,G1038);
  nand GNAME8166(G8166,G8314,G8315);
  not GNAME8167(G8167,G1005);
  not GNAME8168(G8168,G1037);
  nand GNAME8169(G8169,G8318,G8319);
  not GNAME8170(G8170,G1004);
  not GNAME8171(G8171,G1036);
  nand GNAME8172(G8172,G8322,G8323);
  not GNAME8173(G8173,G1035);
  not GNAME8174(G8174,G1003);
  nand GNAME8175(G8175,G8432,G8433);
  nand GNAME8176(G8176,G8335,G8336);
  nand GNAME8177(G8177,G8340,G8341);
  nand GNAME8178(G8178,G8345,G8346);
  nand GNAME8179(G8179,G8350,G8351);
  nand GNAME8180(G8180,G8355,G8356);
  nand GNAME8181(G8181,G8360,G8361);
  nand GNAME8182(G8182,G8365,G8366);
  nand GNAME8183(G8183,G8373,G8374);
  nand GNAME8184(G8184,G8378,G8379);
  nand GNAME8185(G8185,G8383,G8384);
  nand GNAME8186(G8186,G8388,G8389);
  nand GNAME8187(G8187,G8393,G8394);
  nand GNAME8188(G8188,G8398,G8399);
  nand GNAME8189(G8189,G8403,G8404);
  nand GNAME8190(G8190,G8408,G8409);
  nand GNAME8191(G8191,G8413,G8414);
  nand GNAME8192(G8192,G8418,G8419);
  nand GNAME8193(G8193,G8423,G8424);
  nand GNAME8194(G8194,G8428,G8429);
  nand GNAME8195(G8195,G8437,G8438);
  nand GNAME8196(G8196,G8442,G8443);
  nand GNAME8197(G8197,G8447,G8448);
  nand GNAME8198(G8198,G8452,G8453);
  nand GNAME8199(G8199,G8457,G8458);
  nand GNAME8200(G8200,G8462,G8463);
  nand GNAME8201(G8201,G8467,G8468);
  nand GNAME8202(G8202,G8472,G8473);
  nand GNAME8203(G8203,G8477,G8478);
  nand GNAME8204(G8204,G8482,G8483);
  and GNAME8205(G8205,G8430,G8431);
  not GNAME8206(G8206,G1034);
  not GNAME8207(G8207,G1002);
  or GNAME8208(G8208,G1065,G8086);
  or GNAME8209(G8209,G1064,G8087);
  nand GNAME8210(G8210,G8208,G8209);
  nand GNAME8211(G8211,G8087,G1064);
  not GNAME8212(G8212,G8088);
  nand GNAME8213(G8213,G8212,G1031);
  nand GNAME8214(G8214,G8213,G1063);
  nand GNAME8215(G8215,G8089,G8088);
  not GNAME8216(G8216,G8091);
  nand GNAME8217(G8217,G8216,G1030);
  nand GNAME8218(G8218,G8217,G1062);
  nand GNAME8219(G8219,G8092,G8091);
  not GNAME8220(G8220,G8094);
  nand GNAME8221(G8221,G8220,G1029);
  nand GNAME8222(G8222,G8221,G1061);
  nand GNAME8223(G8223,G8095,G8094);
  not GNAME8224(G8224,G8097);
  nand GNAME8225(G8225,G8224,G1028);
  nand GNAME8226(G8226,G8225,G1060);
  nand GNAME8227(G8227,G8098,G8097);
  not GNAME8228(G8228,G8100);
  nand GNAME8229(G8229,G8228,G1027);
  nand GNAME8230(G8230,G8229,G1059);
  nand GNAME8231(G8231,G8101,G8100);
  not GNAME8232(G8232,G8103);
  nand GNAME8233(G8233,G8232,G1026);
  nand GNAME8234(G8234,G8233,G1058);
  nand GNAME8235(G8235,G8104,G8103);
  not GNAME8236(G8236,G8106);
  nand GNAME8237(G8237,G8236,G1025);
  nand GNAME8238(G8238,G8237,G1057);
  nand GNAME8239(G8239,G8107,G8106);
  not GNAME8240(G8240,G8111);
  nand GNAME8241(G8241,G1024,G8240);
  nand GNAME8242(G8242,G8241,G1056);
  nand GNAME8243(G8243,G8110,G8111);
  not GNAME8244(G8244,G8112);
  nand GNAME8245(G8245,G8244,G1023);
  nand GNAME8246(G8246,G8245,G1055);
  nand GNAME8247(G8247,G8113,G8112);
  not GNAME8248(G8248,G8115);
  nand GNAME8249(G8249,G8248,G1022);
  nand GNAME8250(G8250,G8249,G1054);
  nand GNAME8251(G8251,G8116,G8115);
  not GNAME8252(G8252,G8118);
  nand GNAME8253(G8253,G8252,G1021);
  nand GNAME8254(G8254,G8253,G1053);
  nand GNAME8255(G8255,G8119,G8118);
  not GNAME8256(G8256,G8121);
  nand GNAME8257(G8257,G8256,G1020);
  nand GNAME8258(G8258,G8257,G1052);
  nand GNAME8259(G8259,G8122,G8121);
  not GNAME8260(G8260,G8124);
  nand GNAME8261(G8261,G8260,G1019);
  nand GNAME8262(G8262,G8261,G1051);
  nand GNAME8263(G8263,G8125,G8124);
  not GNAME8264(G8264,G8127);
  nand GNAME8265(G8265,G8264,G1018);
  nand GNAME8266(G8266,G8265,G1050);
  nand GNAME8267(G8267,G8128,G8127);
  not GNAME8268(G8268,G8130);
  nand GNAME8269(G8269,G8268,G1017);
  nand GNAME8270(G8270,G8269,G1049);
  nand GNAME8271(G8271,G8131,G8130);
  not GNAME8272(G8272,G8133);
  nand GNAME8273(G8273,G8272,G1016);
  nand GNAME8274(G8274,G8273,G1048);
  nand GNAME8275(G8275,G8134,G8133);
  not GNAME8276(G8276,G8136);
  nand GNAME8277(G8277,G8276,G1015);
  nand GNAME8278(G8278,G8277,G1047);
  nand GNAME8279(G8279,G8137,G8136);
  not GNAME8280(G8280,G8139);
  nand GNAME8281(G8281,G8280,G1014);
  nand GNAME8282(G8282,G8281,G1046);
  nand GNAME8283(G8283,G8140,G8139);
  not GNAME8284(G8284,G8142);
  nand GNAME8285(G8285,G8284,G1013);
  nand GNAME8286(G8286,G8285,G1045);
  nand GNAME8287(G8287,G8143,G8142);
  not GNAME8288(G8288,G8145);
  nand GNAME8289(G8289,G8288,G1012);
  nand GNAME8290(G8290,G8289,G1044);
  nand GNAME8291(G8291,G8146,G8145);
  not GNAME8292(G8292,G8148);
  nand GNAME8293(G8293,G8292,G1011);
  nand GNAME8294(G8294,G8293,G1043);
  nand GNAME8295(G8295,G8149,G8148);
  not GNAME8296(G8296,G8151);
  nand GNAME8297(G8297,G8296,G1010);
  nand GNAME8298(G8298,G8297,G1042);
  nand GNAME8299(G8299,G8152,G8151);
  not GNAME8300(G8300,G8154);
  nand GNAME8301(G8301,G8300,G1009);
  nand GNAME8302(G8302,G8301,G1041);
  nand GNAME8303(G8303,G8155,G8154);
  not GNAME8304(G8304,G8157);
  nand GNAME8305(G8305,G8304,G1008);
  nand GNAME8306(G8306,G8305,G1040);
  nand GNAME8307(G8307,G8158,G8157);
  not GNAME8308(G8308,G8160);
  nand GNAME8309(G8309,G8308,G1007);
  nand GNAME8310(G8310,G8309,G1039);
  nand GNAME8311(G8311,G8161,G8160);
  not GNAME8312(G8312,G8163);
  nand GNAME8313(G8313,G8312,G1006);
  nand GNAME8314(G8314,G8313,G1038);
  nand GNAME8315(G8315,G8164,G8163);
  not GNAME8316(G8316,G8166);
  nand GNAME8317(G8317,G8316,G1005);
  nand GNAME8318(G8318,G8317,G1037);
  nand GNAME8319(G8319,G8167,G8166);
  not GNAME8320(G8320,G8169);
  nand GNAME8321(G8321,G8320,G1004);
  nand GNAME8322(G8322,G8321,G1036);
  nand GNAME8323(G8323,G8170,G8169);
  not GNAME8324(G8324,G8172);
  nand GNAME8325(G8325,G8329,G1003);
  nand GNAME8326(G8326,G8369,G8325,G8327);
  nand GNAME8327(G8327,G8173,G8324);
  nand GNAME8328(G8328,G8174,G8327);
  nand GNAME8329(G8329,G8172,G1035);
  nand GNAME8330(G8330,G8367,G8368,G8328,G8329);
  nand GNAME8331(G8331,G8086,G1065);
  nand GNAME8332(G8332,G8110,G1056);
  nand GNAME8333(G8333,G8109,G1024);
  nand GNAME8334(G8334,G8332,G8333);
  nand GNAME8335(G8335,G8111,G8334);
  nand GNAME8336(G8336,G8240,G8332,G8333);
  nand GNAME8337(G8337,G8107,G1057);
  nand GNAME8338(G8338,G8108,G1025);
  nand GNAME8339(G8339,G8337,G8338);
  nand GNAME8340(G8340,G8106,G8339);
  nand GNAME8341(G8341,G8236,G8337,G8338);
  nand GNAME8342(G8342,G8104,G1058);
  nand GNAME8343(G8343,G8105,G1026);
  nand GNAME8344(G8344,G8342,G8343);
  nand GNAME8345(G8345,G8103,G8344);
  nand GNAME8346(G8346,G8232,G8342,G8343);
  nand GNAME8347(G8347,G8101,G1059);
  nand GNAME8348(G8348,G8102,G1027);
  nand GNAME8349(G8349,G8347,G8348);
  nand GNAME8350(G8350,G8100,G8349);
  nand GNAME8351(G8351,G8228,G8347,G8348);
  nand GNAME8352(G8352,G8098,G1060);
  nand GNAME8353(G8353,G8099,G1028);
  nand GNAME8354(G8354,G8352,G8353);
  nand GNAME8355(G8355,G8097,G8354);
  nand GNAME8356(G8356,G8224,G8352,G8353);
  nand GNAME8357(G8357,G8095,G1061);
  nand GNAME8358(G8358,G8096,G1029);
  nand GNAME8359(G8359,G8357,G8358);
  nand GNAME8360(G8360,G8094,G8359);
  nand GNAME8361(G8361,G8220,G8357,G8358);
  nand GNAME8362(G8362,G8092,G1062);
  nand GNAME8363(G8363,G8093,G1030);
  nand GNAME8364(G8364,G8362,G8363);
  nand GNAME8365(G8365,G8091,G8364);
  nand GNAME8366(G8366,G8216,G8362,G8363);
  nand GNAME8367(G8367,G8207,G1034);
  nand GNAME8368(G8368,G8206,G1002);
  nand GNAME8369(G8369,G8367,G8368);
  nand GNAME8370(G8370,G8173,G1003);
  nand GNAME8371(G8371,G8174,G1035);
  nand GNAME8372(G8372,G8370,G8371);
  nand GNAME8373(G8373,G8172,G8372);
  nand GNAME8374(G8374,G8324,G8370,G8371);
  nand GNAME8375(G8375,G8089,G1063);
  nand GNAME8376(G8376,G8090,G1031);
  nand GNAME8377(G8377,G8375,G8376);
  nand GNAME8378(G8378,G8088,G8377);
  nand GNAME8379(G8379,G8212,G8375,G8376);
  nand GNAME8380(G8380,G8170,G1036);
  nand GNAME8381(G8381,G8171,G1004);
  nand GNAME8382(G8382,G8380,G8381);
  nand GNAME8383(G8383,G8169,G8382);
  nand GNAME8384(G8384,G8320,G8380,G8381);
  nand GNAME8385(G8385,G8167,G1037);
  nand GNAME8386(G8386,G8168,G1005);
  nand GNAME8387(G8387,G8385,G8386);
  nand GNAME8388(G8388,G8166,G8387);
  nand GNAME8389(G8389,G8316,G8385,G8386);
  nand GNAME8390(G8390,G8164,G1038);
  nand GNAME8391(G8391,G8165,G1006);
  nand GNAME8392(G8392,G8390,G8391);
  nand GNAME8393(G8393,G8163,G8392);
  nand GNAME8394(G8394,G8312,G8390,G8391);
  nand GNAME8395(G8395,G8161,G1039);
  nand GNAME8396(G8396,G8162,G1007);
  nand GNAME8397(G8397,G8395,G8396);
  nand GNAME8398(G8398,G8160,G8397);
  nand GNAME8399(G8399,G8308,G8395,G8396);
  nand GNAME8400(G8400,G8158,G1040);
  nand GNAME8401(G8401,G8159,G1008);
  nand GNAME8402(G8402,G8400,G8401);
  nand GNAME8403(G8403,G8157,G8402);
  nand GNAME8404(G8404,G8304,G8400,G8401);
  nand GNAME8405(G8405,G8155,G1041);
  nand GNAME8406(G8406,G8156,G1009);
  nand GNAME8407(G8407,G8405,G8406);
  nand GNAME8408(G8408,G8154,G8407);
  nand GNAME8409(G8409,G8300,G8405,G8406);
  nand GNAME8410(G8410,G8152,G1042);
  nand GNAME8411(G8411,G8153,G1010);
  nand GNAME8412(G8412,G8410,G8411);
  nand GNAME8413(G8413,G8151,G8412);
  nand GNAME8414(G8414,G8296,G8410,G8411);
  nand GNAME8415(G8415,G8149,G1043);
  nand GNAME8416(G8416,G8150,G1011);
  nand GNAME8417(G8417,G8415,G8416);
  nand GNAME8418(G8418,G8148,G8417);
  nand GNAME8419(G8419,G8292,G8415,G8416);
  nand GNAME8420(G8420,G8146,G1044);
  nand GNAME8421(G8421,G8147,G1012);
  nand GNAME8422(G8422,G8420,G8421);
  nand GNAME8423(G8423,G8145,G8422);
  nand GNAME8424(G8424,G8288,G8420,G8421);
  nand GNAME8425(G8425,G8143,G1045);
  nand GNAME8426(G8426,G8144,G1013);
  nand GNAME8427(G8427,G8425,G8426);
  nand GNAME8428(G8428,G8142,G8427);
  nand GNAME8429(G8429,G8284,G8425,G8426);
  or GNAME8430(G8430,G1032,G8208);
  nand GNAME8431(G8431,G8208,G1032);
  nand GNAME8432(G8432,G1064,G8205);
  or GNAME8433(G8433,G1064,G8205);
  nand GNAME8434(G8434,G8140,G1046);
  nand GNAME8435(G8435,G8141,G1014);
  nand GNAME8436(G8436,G8434,G8435);
  nand GNAME8437(G8437,G8139,G8436);
  nand GNAME8438(G8438,G8280,G8434,G8435);
  nand GNAME8439(G8439,G8137,G1047);
  nand GNAME8440(G8440,G8138,G1015);
  nand GNAME8441(G8441,G8439,G8440);
  nand GNAME8442(G8442,G8136,G8441);
  nand GNAME8443(G8443,G8276,G8439,G8440);
  nand GNAME8444(G8444,G8134,G1048);
  nand GNAME8445(G8445,G8135,G1016);
  nand GNAME8446(G8446,G8444,G8445);
  nand GNAME8447(G8447,G8133,G8446);
  nand GNAME8448(G8448,G8272,G8444,G8445);
  nand GNAME8449(G8449,G8131,G1049);
  nand GNAME8450(G8450,G8132,G1017);
  nand GNAME8451(G8451,G8449,G8450);
  nand GNAME8452(G8452,G8130,G8451);
  nand GNAME8453(G8453,G8268,G8449,G8450);
  nand GNAME8454(G8454,G8128,G1050);
  nand GNAME8455(G8455,G8129,G1018);
  nand GNAME8456(G8456,G8454,G8455);
  nand GNAME8457(G8457,G8127,G8456);
  nand GNAME8458(G8458,G8264,G8454,G8455);
  nand GNAME8459(G8459,G8125,G1051);
  nand GNAME8460(G8460,G8126,G1019);
  nand GNAME8461(G8461,G8459,G8460);
  nand GNAME8462(G8462,G8124,G8461);
  nand GNAME8463(G8463,G8260,G8459,G8460);
  nand GNAME8464(G8464,G8122,G1052);
  nand GNAME8465(G8465,G8123,G1020);
  nand GNAME8466(G8466,G8464,G8465);
  nand GNAME8467(G8467,G8121,G8466);
  nand GNAME8468(G8468,G8256,G8464,G8465);
  nand GNAME8469(G8469,G8119,G1053);
  nand GNAME8470(G8470,G8120,G1021);
  nand GNAME8471(G8471,G8469,G8470);
  nand GNAME8472(G8472,G8118,G8471);
  nand GNAME8473(G8473,G8252,G8469,G8470);
  nand GNAME8474(G8474,G8116,G1054);
  nand GNAME8475(G8475,G8117,G1022);
  nand GNAME8476(G8476,G8474,G8475);
  nand GNAME8477(G8477,G8115,G8476);
  nand GNAME8478(G8478,G8248,G8474,G8475);
  nand GNAME8479(G8479,G8113,G1055);
  nand GNAME8480(G8480,G8114,G1023);
  nand GNAME8481(G8481,G8479,G8480);
  nand GNAME8482(G8482,G8112,G8481);
  nand GNAME8483(G8483,G8244,G8479,G8480);
  nand GNAME8484(G8484,G8634,G8630);
  nand GNAME8485(G8485,G8635,G8558);
  not GNAME8486(G8486,G4283);
  not GNAME8487(G8487,G4282);
  nand GNAME8488(G8488,G8562,G8563);
  not GNAME8489(G8489,G4271);
  not GNAME8490(G8490,G4158);
  nand GNAME8491(G8491,G8566,G8567);
  not GNAME8492(G8492,G4270);
  not GNAME8493(G8493,G4157);
  nand GNAME8494(G8494,G8570,G8571);
  not GNAME8495(G8495,G4269);
  not GNAME8496(G8496,G4156);
  nand GNAME8497(G8497,G8574,G8575);
  not GNAME8498(G8498,G4268);
  not GNAME8499(G8499,G4155);
  nand GNAME8500(G8500,G8578,G8579);
  not GNAME8501(G8501,G4267);
  not GNAME8502(G8502,G4154);
  nand GNAME8503(G8503,G8582,G8583);
  not GNAME8504(G8504,G4266);
  not GNAME8505(G8505,G4153);
  nand GNAME8506(G8506,G8586,G8587);
  not GNAME8507(G8507,G4265);
  not GNAME8508(G8508,G4152);
  not GNAME8509(G8509,G4151);
  not GNAME8510(G8510,G4264);
  nand GNAME8511(G8511,G8590,G8591);
  nand GNAME8512(G8512,G8594,G8595);
  not GNAME8513(G8513,G4281);
  not GNAME8514(G8514,G4168);
  nand GNAME8515(G8515,G8598,G8599);
  not GNAME8516(G8516,G4280);
  not GNAME8517(G8517,G4167);
  nand GNAME8518(G8518,G8602,G8603);
  not GNAME8519(G8519,G4279);
  not GNAME8520(G8520,G4166);
  nand GNAME8521(G8521,G8606,G8607);
  not GNAME8522(G8522,G4278);
  not GNAME8523(G8523,G4165);
  nand GNAME8524(G8524,G8610,G8611);
  not GNAME8525(G8525,G4277);
  not GNAME8526(G8526,G4164);
  nand GNAME8527(G8527,G8614,G8615);
  not GNAME8528(G8528,G4276);
  not GNAME8529(G8529,G4163);
  nand GNAME8530(G8530,G8618,G8619);
  not GNAME8531(G8531,G4275);
  not GNAME8532(G8532,G4162);
  nand GNAME8533(G8533,G8622,G8623);
  not GNAME8534(G8534,G4274);
  not GNAME8535(G8535,G4161);
  nand GNAME8536(G8536,G8626,G8627);
  not GNAME8537(G8537,G4160);
  not GNAME8538(G8538,G4273);
  nand GNAME8539(G8539,G8678,G8679);
  nand GNAME8540(G8540,G8639,G8640);
  nand GNAME8541(G8541,G8644,G8645);
  nand GNAME8542(G8542,G8649,G8650);
  nand GNAME8543(G8543,G8654,G8655);
  nand GNAME8544(G8544,G8659,G8660);
  nand GNAME8545(G8545,G8664,G8665);
  nand GNAME8546(G8546,G8669,G8670);
  nand GNAME8547(G8547,G8674,G8675);
  nand GNAME8548(G8548,G8686,G8687);
  nand GNAME8549(G8549,G8691,G8692);
  nand GNAME8550(G8550,G8696,G8697);
  nand GNAME8551(G8551,G8701,G8702);
  nand GNAME8552(G8552,G8706,G8707);
  nand GNAME8553(G8553,G8711,G8712);
  nand GNAME8554(G8554,G8716,G8717);
  nand GNAME8555(G8555,G8721,G8722);
  nand GNAME8556(G8556,G8726,G8727);
  and GNAME8557(G8557,G8676,G8677);
  or GNAME8558(G8558,G4169,G8486);
  not GNAME8559(G8559,G4175);
  not GNAME8560(G8560,G4272);
  or GNAME8561(G8561,G4159,G8487);
  nand GNAME8562(G8562,G8558,G8561);
  nand GNAME8563(G8563,G8487,G4159);
  not GNAME8564(G8564,G8488);
  nand GNAME8565(G8565,G8564,G4271);
  nand GNAME8566(G8566,G8565,G4158);
  nand GNAME8567(G8567,G8489,G8488);
  not GNAME8568(G8568,G8491);
  nand GNAME8569(G8569,G8568,G4270);
  nand GNAME8570(G8570,G8569,G4157);
  nand GNAME8571(G8571,G8492,G8491);
  not GNAME8572(G8572,G8494);
  nand GNAME8573(G8573,G8572,G4269);
  nand GNAME8574(G8574,G8573,G4156);
  nand GNAME8575(G8575,G8495,G8494);
  not GNAME8576(G8576,G8497);
  nand GNAME8577(G8577,G8576,G4268);
  nand GNAME8578(G8578,G8577,G4155);
  nand GNAME8579(G8579,G8498,G8497);
  not GNAME8580(G8580,G8500);
  nand GNAME8581(G8581,G8580,G4267);
  nand GNAME8582(G8582,G8581,G4154);
  nand GNAME8583(G8583,G8501,G8500);
  not GNAME8584(G8584,G8503);
  nand GNAME8585(G8585,G8584,G4266);
  nand GNAME8586(G8586,G8585,G4153);
  nand GNAME8587(G8587,G8504,G8503);
  not GNAME8588(G8588,G8506);
  nand GNAME8589(G8589,G8588,G4265);
  nand GNAME8590(G8590,G8589,G4152);
  nand GNAME8591(G8591,G8507,G8506);
  not GNAME8592(G8592,G8511);
  nand GNAME8593(G8593,G4264,G8592);
  nand GNAME8594(G8594,G8593,G4151);
  nand GNAME8595(G8595,G8510,G8511);
  not GNAME8596(G8596,G8512);
  nand GNAME8597(G8597,G8596,G4281);
  nand GNAME8598(G8598,G8597,G4168);
  nand GNAME8599(G8599,G8513,G8512);
  not GNAME8600(G8600,G8515);
  nand GNAME8601(G8601,G8600,G4280);
  nand GNAME8602(G8602,G8601,G4167);
  nand GNAME8603(G8603,G8516,G8515);
  not GNAME8604(G8604,G8518);
  nand GNAME8605(G8605,G8604,G4279);
  nand GNAME8606(G8606,G8605,G4166);
  nand GNAME8607(G8607,G8519,G8518);
  not GNAME8608(G8608,G8521);
  nand GNAME8609(G8609,G8608,G4278);
  nand GNAME8610(G8610,G8609,G4165);
  nand GNAME8611(G8611,G8522,G8521);
  not GNAME8612(G8612,G8524);
  nand GNAME8613(G8613,G8612,G4277);
  nand GNAME8614(G8614,G8613,G4164);
  nand GNAME8615(G8615,G8525,G8524);
  not GNAME8616(G8616,G8527);
  nand GNAME8617(G8617,G8616,G4276);
  nand GNAME8618(G8618,G8617,G4163);
  nand GNAME8619(G8619,G8528,G8527);
  not GNAME8620(G8620,G8530);
  nand GNAME8621(G8621,G8620,G4275);
  nand GNAME8622(G8622,G8621,G4162);
  nand GNAME8623(G8623,G8531,G8530);
  not GNAME8624(G8624,G8533);
  nand GNAME8625(G8625,G8624,G4274);
  nand GNAME8626(G8626,G8625,G4161);
  nand GNAME8627(G8627,G8534,G8533);
  not GNAME8628(G8628,G8536);
  nand GNAME8629(G8629,G8633,G4273);
  nand GNAME8630(G8630,G8682,G8629,G8631);
  nand GNAME8631(G8631,G8537,G8628);
  nand GNAME8632(G8632,G8538,G8631);
  nand GNAME8633(G8633,G8536,G4160);
  nand GNAME8634(G8634,G8680,G8681,G8632,G8633);
  nand GNAME8635(G8635,G8486,G4169);
  nand GNAME8636(G8636,G8510,G4151);
  nand GNAME8637(G8637,G8509,G4264);
  nand GNAME8638(G8638,G8636,G8637);
  nand GNAME8639(G8639,G8511,G8638);
  nand GNAME8640(G8640,G8592,G8636,G8637);
  nand GNAME8641(G8641,G8507,G4152);
  nand GNAME8642(G8642,G8508,G4265);
  nand GNAME8643(G8643,G8641,G8642);
  nand GNAME8644(G8644,G8506,G8643);
  nand GNAME8645(G8645,G8588,G8641,G8642);
  nand GNAME8646(G8646,G8504,G4153);
  nand GNAME8647(G8647,G8505,G4266);
  nand GNAME8648(G8648,G8646,G8647);
  nand GNAME8649(G8649,G8503,G8648);
  nand GNAME8650(G8650,G8584,G8646,G8647);
  nand GNAME8651(G8651,G8501,G4154);
  nand GNAME8652(G8652,G8502,G4267);
  nand GNAME8653(G8653,G8651,G8652);
  nand GNAME8654(G8654,G8500,G8653);
  nand GNAME8655(G8655,G8580,G8651,G8652);
  nand GNAME8656(G8656,G8498,G4155);
  nand GNAME8657(G8657,G8499,G4268);
  nand GNAME8658(G8658,G8656,G8657);
  nand GNAME8659(G8659,G8497,G8658);
  nand GNAME8660(G8660,G8576,G8656,G8657);
  nand GNAME8661(G8661,G8495,G4156);
  nand GNAME8662(G8662,G8496,G4269);
  nand GNAME8663(G8663,G8661,G8662);
  nand GNAME8664(G8664,G8494,G8663);
  nand GNAME8665(G8665,G8572,G8661,G8662);
  nand GNAME8666(G8666,G8492,G4157);
  nand GNAME8667(G8667,G8493,G4270);
  nand GNAME8668(G8668,G8666,G8667);
  nand GNAME8669(G8669,G8491,G8668);
  nand GNAME8670(G8670,G8568,G8666,G8667);
  nand GNAME8671(G8671,G8489,G4158);
  nand GNAME8672(G8672,G8490,G4271);
  nand GNAME8673(G8673,G8671,G8672);
  nand GNAME8674(G8674,G8488,G8673);
  nand GNAME8675(G8675,G8564,G8671,G8672);
  or GNAME8676(G8676,G4282,G8558);
  nand GNAME8677(G8677,G8558,G4282);
  nand GNAME8678(G8678,G4159,G8557);
  or GNAME8679(G8679,G4159,G8557);
  nand GNAME8680(G8680,G8560,G4175);
  nand GNAME8681(G8681,G8559,G4272);
  nand GNAME8682(G8682,G8680,G8681);
  nand GNAME8683(G8683,G8537,G4273);
  nand GNAME8684(G8684,G8538,G4160);
  nand GNAME8685(G8685,G8683,G8684);
  nand GNAME8686(G8686,G8536,G8685);
  nand GNAME8687(G8687,G8628,G8683,G8684);
  nand GNAME8688(G8688,G8534,G4161);
  nand GNAME8689(G8689,G8535,G4274);
  nand GNAME8690(G8690,G8688,G8689);
  nand GNAME8691(G8691,G8533,G8690);
  nand GNAME8692(G8692,G8624,G8688,G8689);
  nand GNAME8693(G8693,G8531,G4162);
  nand GNAME8694(G8694,G8532,G4275);
  nand GNAME8695(G8695,G8693,G8694);
  nand GNAME8696(G8696,G8530,G8695);
  nand GNAME8697(G8697,G8620,G8693,G8694);
  nand GNAME8698(G8698,G8528,G4163);
  nand GNAME8699(G8699,G8529,G4276);
  nand GNAME8700(G8700,G8698,G8699);
  nand GNAME8701(G8701,G8527,G8700);
  nand GNAME8702(G8702,G8616,G8698,G8699);
  nand GNAME8703(G8703,G8525,G4164);
  nand GNAME8704(G8704,G8526,G4277);
  nand GNAME8705(G8705,G8703,G8704);
  nand GNAME8706(G8706,G8524,G8705);
  nand GNAME8707(G8707,G8612,G8703,G8704);
  nand GNAME8708(G8708,G8522,G4165);
  nand GNAME8709(G8709,G8523,G4278);
  nand GNAME8710(G8710,G8708,G8709);
  nand GNAME8711(G8711,G8521,G8710);
  nand GNAME8712(G8712,G8608,G8708,G8709);
  nand GNAME8713(G8713,G8519,G4166);
  nand GNAME8714(G8714,G8520,G4279);
  nand GNAME8715(G8715,G8713,G8714);
  nand GNAME8716(G8716,G8518,G8715);
  nand GNAME8717(G8717,G8604,G8713,G8714);
  nand GNAME8718(G8718,G8516,G4167);
  nand GNAME8719(G8719,G8517,G4280);
  nand GNAME8720(G8720,G8718,G8719);
  nand GNAME8721(G8721,G8515,G8720);
  nand GNAME8722(G8722,G8600,G8718,G8719);
  nand GNAME8723(G8723,G8513,G4168);
  nand GNAME8724(G8724,G8514,G4281);
  nand GNAME8725(G8725,G8723,G8724);
  nand GNAME8726(G8726,G8512,G8725);
  nand GNAME8727(G8727,G8596,G8723,G8724);
  nand GNAME8728(G8728,G8851,G8854,G8855);
  not GNAME8729(G8729,G3740);
  not GNAME8730(G8730,G3773);
  not GNAME8731(G8731,G3736);
  not GNAME8732(G8732,G3771);
  not GNAME8733(G8733,G3732);
  not GNAME8734(G8734,G3769);
  not GNAME8735(G8735,G3728);
  not GNAME8736(G8736,G3767);
  not GNAME8737(G8737,G3724);
  not GNAME8738(G8738,G3765);
  not GNAME8739(G8739,G3720);
  not GNAME8740(G8740,G3763);
  not GNAME8741(G8741,G3716);
  not GNAME8742(G8742,G3761);
  not GNAME8743(G8743,G3712);
  not GNAME8744(G8744,G3759);
  not GNAME8745(G8745,G3708);
  not GNAME8746(G8746,G3757);
  not GNAME8747(G8747,G3704);
  not GNAME8748(G8748,G3755);
  not GNAME8749(G8749,G3700);
  not GNAME8750(G8750,G3753);
  not GNAME8751(G8751,G3696);
  not GNAME8752(G8752,G3751);
  not GNAME8753(G8753,G3692);
  not GNAME8754(G8754,G3749);
  not GNAME8755(G8755,G3688);
  not GNAME8756(G8756,G3747);
  not GNAME8757(G8757,G3684);
  not GNAME8758(G8758,G3682);
  not GNAME8759(G8759,G3744);
  not GNAME8760(G8760,G3742);
  or GNAME8761(G8761,G3774,G8729);
  nand GNAME8762(G8762,G3775,G8760,G8761);
  or GNAME8763(G8763,G3738,G8730);
  nand GNAME8764(G8764,G8729,G3774);
  nand GNAME8765(G8765,G8764,G8762,G8763);
  or GNAME8766(G8766,G3772,G8731);
  nand GNAME8767(G8767,G8730,G3738);
  nand GNAME8768(G8768,G8767,G8765,G8766);
  or GNAME8769(G8769,G3734,G8732);
  nand GNAME8770(G8770,G8731,G3772);
  nand GNAME8771(G8771,G8770,G8768,G8769);
  or GNAME8772(G8772,G3770,G8733);
  nand GNAME8773(G8773,G8732,G3734);
  nand GNAME8774(G8774,G8773,G8771,G8772);
  or GNAME8775(G8775,G3730,G8734);
  nand GNAME8776(G8776,G8733,G3770);
  nand GNAME8777(G8777,G8776,G8774,G8775);
  or GNAME8778(G8778,G3768,G8735);
  nand GNAME8779(G8779,G8734,G3730);
  nand GNAME8780(G8780,G8779,G8777,G8778);
  or GNAME8781(G8781,G3726,G8736);
  nand GNAME8782(G8782,G8735,G3768);
  nand GNAME8783(G8783,G8782,G8780,G8781);
  or GNAME8784(G8784,G3766,G8737);
  nand GNAME8785(G8785,G8736,G3726);
  nand GNAME8786(G8786,G8785,G8783,G8784);
  or GNAME8787(G8787,G3722,G8738);
  nand GNAME8788(G8788,G8737,G3766);
  nand GNAME8789(G8789,G8788,G8786,G8787);
  or GNAME8790(G8790,G3764,G8739);
  nand GNAME8791(G8791,G8738,G3722);
  nand GNAME8792(G8792,G8791,G8789,G8790);
  or GNAME8793(G8793,G3718,G8740);
  nand GNAME8794(G8794,G8739,G3764);
  nand GNAME8795(G8795,G8794,G8792,G8793);
  or GNAME8796(G8796,G3762,G8741);
  nand GNAME8797(G8797,G8740,G3718);
  nand GNAME8798(G8798,G8797,G8795,G8796);
  or GNAME8799(G8799,G3714,G8742);
  nand GNAME8800(G8800,G8741,G3762);
  nand GNAME8801(G8801,G8800,G8798,G8799);
  or GNAME8802(G8802,G3760,G8743);
  nand GNAME8803(G8803,G8742,G3714);
  nand GNAME8804(G8804,G8803,G8801,G8802);
  or GNAME8805(G8805,G3710,G8744);
  nand GNAME8806(G8806,G8743,G3760);
  nand GNAME8807(G8807,G8806,G8804,G8805);
  or GNAME8808(G8808,G3758,G8745);
  nand GNAME8809(G8809,G8744,G3710);
  nand GNAME8810(G8810,G8809,G8807,G8808);
  or GNAME8811(G8811,G3706,G8746);
  nand GNAME8812(G8812,G8745,G3758);
  nand GNAME8813(G8813,G8812,G8810,G8811);
  or GNAME8814(G8814,G3756,G8747);
  nand GNAME8815(G8815,G8746,G3706);
  nand GNAME8816(G8816,G8815,G8813,G8814);
  or GNAME8817(G8817,G3702,G8748);
  nand GNAME8818(G8818,G8747,G3756);
  nand GNAME8819(G8819,G8818,G8816,G8817);
  or GNAME8820(G8820,G3754,G8749);
  nand GNAME8821(G8821,G8748,G3702);
  nand GNAME8822(G8822,G8821,G8819,G8820);
  or GNAME8823(G8823,G3698,G8750);
  nand GNAME8824(G8824,G8749,G3754);
  nand GNAME8825(G8825,G8824,G8822,G8823);
  or GNAME8826(G8826,G3752,G8751);
  nand GNAME8827(G8827,G8750,G3698);
  nand GNAME8828(G8828,G8827,G8825,G8826);
  or GNAME8829(G8829,G3694,G8752);
  nand GNAME8830(G8830,G8751,G3752);
  nand GNAME8831(G8831,G8830,G8828,G8829);
  or GNAME8832(G8832,G3750,G8753);
  nand GNAME8833(G8833,G8752,G3694);
  nand GNAME8834(G8834,G8833,G8831,G8832);
  or GNAME8835(G8835,G3690,G8754);
  nand GNAME8836(G8836,G8753,G3750);
  nand GNAME8837(G8837,G8836,G8834,G8835);
  or GNAME8838(G8838,G3748,G8755);
  nand GNAME8839(G8839,G8754,G3690);
  nand GNAME8840(G8840,G8839,G8837,G8838);
  or GNAME8841(G8841,G3686,G8756);
  nand GNAME8842(G8842,G8755,G3748);
  nand GNAME8843(G8843,G8842,G8840,G8841);
  or GNAME8844(G8844,G3746,G8757);
  nand GNAME8845(G8845,G8756,G3686);
  nand GNAME8846(G8846,G8845,G8843,G8844);
  nand GNAME8847(G8847,G8758,G3745);
  nand GNAME8848(G8848,G8757,G3746);
  nand GNAME8849(G8849,G8848,G8846,G8847);
  or GNAME8850(G8850,G3745,G8758);
  nand GNAME8851(G8851,G8852,G8853,G8849,G8850);
  or GNAME8852(G8852,G3680,G8759);
  nand GNAME8853(G8853,G8759,G3680);
  or GNAME8854(G8854,G3680,G4050,G8759);
  nand GNAME8855(G8855,G3680,G8759,G4050);
  and GNAME8856(G8856,G8875,G8921);
  and GNAME8857(G8857,G8877,G8918);
  and GNAME8858(G8858,G8879,G8916);
  and GNAME8859(G8859,G8881,G8914);
  and GNAME8860(G8860,G8883,G8912);
  and GNAME8861(G8861,G8885,G8910);
  and GNAME8862(G8862,G8871,G8909);
  and GNAME8863(G8863,G8873,G8906);
  and GNAME8864(G8864,G8874,G8905);
  and GNAME8865(G8865,G8872,G8907);
  and GNAME8866(G8866,G8884,G8911);
  and GNAME8867(G8867,G8882,G8913);
  and GNAME8868(G8868,G8880,G8915);
  and GNAME8869(G8869,G8878,G8917);
  and GNAME8870(G8870,G8876,G8919);
  or GNAME8871(G8871,G22802,G22803,G22801);
  or GNAME8872(G8872,G8871,G22804,G22805);
  or GNAME8873(G8873,G8872,G22807,G22806);
  or GNAME8874(G8874,G8873,G22808,G22809);
  or GNAME8875(G8875,G8874,G22810,G22811);
  or GNAME8876(G8876,G8875,G22812,G22813);
  or GNAME8877(G8877,G8876,G22815,G22814);
  or GNAME8878(G8878,G8877,G22816,G22817);
  or GNAME8879(G8879,G8878,G22819,G22818);
  or GNAME8880(G8880,G8879,G22820,G22821);
  or GNAME8881(G8881,G8880,G22823,G22822);
  or GNAME8882(G8882,G8881,G22824,G22825);
  or GNAME8883(G8883,G8882,G22827,G22826);
  or GNAME8884(G8884,G8883,G22828,G22829);
  or GNAME8885(G8885,G22830,G8884);
  nand GNAME8886(G8886,G8941,G8942);
  not GNAME8887(G8887,G22810);
  and GNAME8888(G8888,G8922,G8920);
  and GNAME8889(G8889,G8923,G8924);
  and GNAME8890(G8890,G8925,G8926);
  and GNAME8891(G8891,G8927,G8928);
  and GNAME8892(G8892,G8929,G8930);
  and GNAME8893(G8893,G8931,G8932);
  and GNAME8894(G8894,G8933,G8934);
  and GNAME8895(G8895,G8935,G8936);
  and GNAME8896(G8896,G8937,G8938);
  and GNAME8897(G8897,G8939,G8940);
  not GNAME8898(G8898,G22801);
  and GNAME8899(G8899,G8943,G8944);
  and GNAME8900(G8900,G8945,G8946);
  and GNAME8901(G8901,G8947,G8948);
  and GNAME8902(G8902,G8949,G8950);
  and GNAME8903(G8903,G8951,G8952);
  not GNAME8904(G8904,G8874);
  nand GNAME8905(G8905,G8924,G22809);
  nand GNAME8906(G8906,G8926,G22807);
  nand GNAME8907(G8907,G8928,G22805);
  or GNAME8908(G8908,G22802,G22801);
  nand GNAME8909(G8909,G8908,G22803);
  nand GNAME8910(G8910,G8884,G22830);
  nand GNAME8911(G8911,G8934,G22829);
  nand GNAME8912(G8912,G8936,G22827);
  nand GNAME8913(G8913,G8938,G22825);
  nand GNAME8914(G8914,G8940,G22823);
  nand GNAME8915(G8915,G8944,G22821);
  nand GNAME8916(G8916,G8946,G22819);
  nand GNAME8917(G8917,G8948,G22817);
  nand GNAME8918(G8918,G8950,G22815);
  nand GNAME8919(G8919,G8952,G22813);
  nand GNAME8920(G8920,G8887,G8904);
  nand GNAME8921(G8921,G8920,G22811);
  nand GNAME8922(G8922,G8874,G22810);
  nand GNAME8923(G8923,G8873,G22808);
  or GNAME8924(G8924,G22808,G8873);
  nand GNAME8925(G8925,G8872,G22806);
  or GNAME8926(G8926,G22806,G8872);
  nand GNAME8927(G8927,G8871,G22804);
  or GNAME8928(G8928,G22804,G8871);
  nand GNAME8929(G8929,G8932,G22832);
  or GNAME8930(G8930,G22832,G8932);
  nand GNAME8931(G8931,G8885,G22831);
  or GNAME8932(G8932,G22831,G8885);
  nand GNAME8933(G8933,G8883,G22828);
  or GNAME8934(G8934,G22828,G8883);
  nand GNAME8935(G8935,G8882,G22826);
  or GNAME8936(G8936,G22826,G8882);
  nand GNAME8937(G8937,G8881,G22824);
  or GNAME8938(G8938,G22824,G8881);
  nand GNAME8939(G8939,G8880,G22822);
  or GNAME8940(G8940,G22822,G8880);
  or GNAME8941(G8941,G22802,G8898);
  nand GNAME8942(G8942,G8898,G22802);
  nand GNAME8943(G8943,G8879,G22820);
  or GNAME8944(G8944,G22820,G8879);
  nand GNAME8945(G8945,G8878,G22818);
  or GNAME8946(G8946,G22818,G8878);
  nand GNAME8947(G8947,G8877,G22816);
  or GNAME8948(G8948,G22816,G8877);
  nand GNAME8949(G8949,G8876,G22814);
  or GNAME8950(G8950,G22814,G8876);
  nand GNAME8951(G8951,G8875,G22812);
  or GNAME8952(G8952,G22812,G8875);
  and GNAME8953(G8953,G9218,G9219);
  and GNAME8954(G8954,G9214,G9215);
  and GNAME8955(G8955,G9139,G9140);
  not GNAME8956(G8956,G3776);
  not GNAME8957(G8957,G3833);
  not GNAME8958(G8958,G3834);
  not GNAME8959(G8959,G3837);
  not GNAME8960(G8960,G3838);
  not GNAME8961(G8961,G3839);
  not GNAME8962(G8962,G3836);
  not GNAME8963(G8963,G3835);
  not GNAME8964(G8964,G3832);
  not GNAME8965(G8965,G3831);
  not GNAME8966(G8966,G3830);
  and GNAME8967(G8967,G9127,G9097);
  not GNAME8968(G8968,G3829);
  not GNAME8969(G8969,G3828);
  not GNAME8970(G8970,G3827);
  not GNAME8971(G8971,G3826);
  not GNAME8972(G8972,G3825);
  not GNAME8973(G8973,G3824);
  not GNAME8974(G8974,G3823);
  not GNAME8975(G8975,G3822);
  not GNAME8976(G8976,G3821);
  not GNAME8977(G8977,G3820);
  not GNAME8978(G8978,G3819);
  not GNAME8979(G8979,G3818);
  not GNAME8980(G8980,G3817);
  not GNAME8981(G8981,G3816);
  not GNAME8982(G8982,G3815);
  not GNAME8983(G8983,G3814);
  not GNAME8984(G8984,G3813);
  not GNAME8985(G8985,G3812);
  not GNAME8986(G8986,G3811);
  not GNAME8987(G8987,G3809);
  and GNAME8988(G8988,G9119,G9099);
  and GNAME8989(G8989,G9168,G9101);
  and GNAME8990(G8990,G9313,G9314);
  nand GNAME8991(G8991,G9363,G9364);
  nand GNAME8992(G8992,G9254,G9255);
  nand GNAME8993(G8993,G9260,G9261);
  nand GNAME8994(G8994,G9319,G9320);
  nand GNAME8995(G8995,G9321,G9322);
  nand GNAME8996(G8996,G9355,G9356);
  nand GNAME8997(G8997,G9361,G9362);
  not GNAME8998(G8998,G3800);
  not GNAME8999(G8999,G3802);
  not GNAME9000(G9000,G3804);
  not GNAME9001(G9001,G3806);
  not GNAME9002(G9002,G3807);
  not GNAME9003(G9003,G3803);
  not GNAME9004(G9004,G3799);
  not GNAME9005(G9005,G3798);
  nand GNAME9006(G9006,G9134,G9132);
  and GNAME9007(G9007,G9136,G9135);
  and GNAME9008(G9008,G9250,G9251);
  nand GNAME9009(G9009,G9131,G9104);
  and GNAME9010(G9010,G9133,G9132);
  and GNAME9011(G9011,G9252,G9253);
  nor GNAME9012(G9012,G9366,G8967);
  nand GNAME9013(G9013,G9125,G9109);
  and GNAME9014(G9014,G9126,G9106);
  and GNAME9015(G9015,G9256,G9257);
  nand GNAME9016(G9016,G9123,G9110);
  and GNAME9017(G9017,G9124,G9109);
  and GNAME9018(G9018,G9258,G9259);
  nor GNAME9019(G9019,G9365,G8988);
  not GNAME9020(G9020,G3796);
  not GNAME9021(G9021,G3795);
  not GNAME9022(G9022,G3794);
  not GNAME9023(G9023,G3792);
  not GNAME9024(G9024,G3791);
  not GNAME9025(G9025,G3790);
  not GNAME9026(G9026,G3789);
  not GNAME9027(G9027,G3788);
  not GNAME9028(G9028,G3787);
  not GNAME9029(G9029,G3786);
  not GNAME9030(G9030,G3785);
  not GNAME9031(G9031,G3784);
  not GNAME9032(G9032,G3783);
  not GNAME9033(G9033,G3782);
  not GNAME9034(G9034,G3781);
  not GNAME9035(G9035,G3780);
  not GNAME9036(G9036,G3779);
  not GNAME9037(G9037,G3808);
  and GNAME9038(G9038,G9210,G9103);
  and GNAME9039(G9039,G9208,G9144);
  nand GNAME9040(G9040,G9206,G9145);
  and GNAME9041(G9041,G9207,G9144);
  and GNAME9042(G9042,G9323,G9324);
  nand GNAME9043(G9043,G9204,G9146);
  and GNAME9044(G9044,G9205,G9145);
  and GNAME9045(G9045,G9325,G9326);
  nand GNAME9046(G9046,G9202,G9147);
  and GNAME9047(G9047,G9203,G9146);
  and GNAME9048(G9048,G9327,G9328);
  nand GNAME9049(G9049,G9200,G9148);
  and GNAME9050(G9050,G9201,G9147);
  and GNAME9051(G9051,G9329,G9330);
  nand GNAME9052(G9052,G9198,G9149);
  and GNAME9053(G9053,G9199,G9148);
  and GNAME9054(G9054,G9331,G9332);
  nand GNAME9055(G9055,G9196,G9150);
  and GNAME9056(G9056,G9197,G9149);
  and GNAME9057(G9057,G9333,G9334);
  nand GNAME9058(G9058,G9194,G9151);
  and GNAME9059(G9059,G9195,G9150);
  and GNAME9060(G9060,G9335,G9336);
  nand GNAME9061(G9061,G9192,G9152);
  and GNAME9062(G9062,G9193,G9151);
  and GNAME9063(G9063,G9337,G9338);
  nand GNAME9064(G9064,G9190,G9153);
  and GNAME9065(G9065,G9191,G9152);
  and GNAME9066(G9066,G9339,G9340);
  nand GNAME9067(G9067,G9188,G9154);
  and GNAME9068(G9068,G9189,G9153);
  and GNAME9069(G9069,G9341,G9342);
  nand GNAME9070(G9070,G9117,G9115);
  and GNAME9071(G9071,G9118,G9112);
  and GNAME9072(G9072,G9343,G9344);
  nand GNAME9073(G9073,G9186,G9155);
  and GNAME9074(G9074,G9187,G9154);
  and GNAME9075(G9075,G9345,G9346);
  nand GNAME9076(G9076,G9184,G9156);
  and GNAME9077(G9077,G9185,G9155);
  and GNAME9078(G9078,G9347,G9348);
  nand GNAME9079(G9079,G9182,G9157);
  and GNAME9080(G9080,G9183,G9156);
  and GNAME9081(G9081,G9349,G9350);
  nand GNAME9082(G9082,G9180,G9158);
  and GNAME9083(G9083,G9181,G9157);
  and GNAME9084(G9084,G9351,G9352);
  nand GNAME9085(G9085,G9178,G9102);
  and GNAME9086(G9086,G9179,G9158);
  and GNAME9087(G9087,G9353,G9354);
  and GNAME9088(G9088,G9176,G9162);
  nand GNAME9089(G9089,G9174,G9163);
  and GNAME9090(G9090,G9175,G9162);
  and GNAME9091(G9091,G9357,G9358);
  nand GNAME9092(G9092,G9172,G9164);
  and GNAME9093(G9093,G9173,G9163);
  and GNAME9094(G9094,G9359,G9360);
  nor GNAME9095(G9095,G9367,G8989);
  and GNAME9096(G9096,G9116,G9115);
  nand GNAME9097(G9097,G9108,G8957,G9107);
  nand GNAME9098(G9098,G9142,G8987,G9141);
  nand GNAME9099(G9099,G9114,G8959,G9113);
  nand GNAME9100(G9100,G9160,G8972,G9159);
  nand GNAME9101(G9101,G9167,G8968,G9166);
  nand GNAME9102(G9102,G9161,G3825);
  nand GNAME9103(G9103,G9143,G3809);
  nand GNAME9104(G9104,G9243,G3832);
  nand GNAME9105(G9105,G8964,G9226,G9227);
  nand GNAME9106(G9106,G9230,G3834);
  or GNAME9107(G9107,G3801,G8956);
  nand GNAME9108(G9108,G8956,G3801);
  nand GNAME9109(G9109,G9242,G3835);
  nand GNAME9110(G9110,G9239,G3836);
  nand GNAME9111(G9111,G8962,G9231,G9232);
  nand GNAME9112(G9112,G9235,G3838);
  or GNAME9113(G9113,G3805,G8956);
  nand GNAME9114(G9114,G8956,G3805);
  nand GNAME9115(G9115,G9238,G3839);
  nand GNAME9116(G9116,G8961,G9236,G9237);
  nand GNAME9117(G9117,G9116,G3776);
  nand GNAME9118(G9118,G8960,G9233,G9234);
  nand GNAME9119(G9119,G9112,G9212);
  nand GNAME9120(G9120,G9113,G9114);
  nand GNAME9121(G9121,G9120,G3837);
  not GNAME9122(G9122,G9019);
  nand GNAME9123(G9123,G9111,G9122);
  nand GNAME9124(G9124,G8963,G9240,G9241);
  nand GNAME9125(G9125,G9016,G9124);
  nand GNAME9126(G9126,G8958,G9228,G9229);
  nand GNAME9127(G9127,G9106,G9137);
  nand GNAME9128(G9128,G9107,G9108);
  nand GNAME9129(G9129,G9128,G3833);
  not GNAME9130(G9130,G9012);
  nand GNAME9131(G9131,G9105,G9130);
  nand GNAME9132(G9132,G9246,G3831);
  nand GNAME9133(G9133,G8965,G9244,G9245);
  nand GNAME9134(G9134,G9009,G9133);
  nand GNAME9135(G9135,G9249,G3830);
  nand GNAME9136(G9136,G8966,G9247,G9248);
  nand GNAME9137(G9137,G9013,G9126);
  nand GNAME9138(G9138,G9097,G9129);
  nand GNAME9139(G9139,G9138,G9106,G9137);
  nand GNAME9140(G9140,G9129,G8967);
  or GNAME9141(G9141,G3777,G8956);
  nand GNAME9142(G9142,G8956,G3777);
  nand GNAME9143(G9143,G9142,G9141);
  nand GNAME9144(G9144,G9315,G3810);
  nand GNAME9145(G9145,G9312,G3811);
  nand GNAME9146(G9146,G9309,G3812);
  nand GNAME9147(G9147,G9306,G3813);
  nand GNAME9148(G9148,G9303,G3814);
  nand GNAME9149(G9149,G9300,G3815);
  nand GNAME9150(G9150,G9297,G3816);
  nand GNAME9151(G9151,G9294,G3817);
  nand GNAME9152(G9152,G9291,G3818);
  nand GNAME9153(G9153,G9288,G3819);
  nand GNAME9154(G9154,G9285,G3820);
  nand GNAME9155(G9155,G9282,G3821);
  nand GNAME9156(G9156,G9279,G3822);
  nand GNAME9157(G9157,G9276,G3823);
  nand GNAME9158(G9158,G9273,G3824);
  or GNAME9159(G9159,G3793,G8956);
  nand GNAME9160(G9160,G8956,G3793);
  nand GNAME9161(G9161,G9160,G9159);
  nand GNAME9162(G9162,G9270,G3826);
  nand GNAME9163(G9163,G9267,G3827);
  nand GNAME9164(G9164,G9264,G3828);
  nand GNAME9165(G9165,G8969,G9262,G9263);
  or GNAME9166(G9166,G3797,G8956);
  nand GNAME9167(G9167,G8956,G3797);
  nand GNAME9168(G9168,G9135,G9217);
  nand GNAME9169(G9169,G9166,G9167);
  nand GNAME9170(G9170,G9169,G3829);
  not GNAME9171(G9171,G9095);
  nand GNAME9172(G9172,G9165,G9171);
  nand GNAME9173(G9173,G8970,G9265,G9266);
  nand GNAME9174(G9174,G9092,G9173);
  nand GNAME9175(G9175,G8971,G9268,G9269);
  nand GNAME9176(G9176,G9089,G9175);
  not GNAME9177(G9177,G9088);
  nand GNAME9178(G9178,G9100,G9177);
  nand GNAME9179(G9179,G8973,G9271,G9272);
  nand GNAME9180(G9180,G9085,G9179);
  nand GNAME9181(G9181,G8974,G9274,G9275);
  nand GNAME9182(G9182,G9082,G9181);
  nand GNAME9183(G9183,G8975,G9277,G9278);
  nand GNAME9184(G9184,G9079,G9183);
  nand GNAME9185(G9185,G8976,G9280,G9281);
  nand GNAME9186(G9186,G9076,G9185);
  nand GNAME9187(G9187,G8977,G9283,G9284);
  nand GNAME9188(G9188,G9073,G9187);
  nand GNAME9189(G9189,G8978,G9286,G9287);
  nand GNAME9190(G9190,G9067,G9189);
  nand GNAME9191(G9191,G8979,G9289,G9290);
  nand GNAME9192(G9192,G9064,G9191);
  nand GNAME9193(G9193,G8980,G9292,G9293);
  nand GNAME9194(G9194,G9061,G9193);
  nand GNAME9195(G9195,G8981,G9295,G9296);
  nand GNAME9196(G9196,G9058,G9195);
  nand GNAME9197(G9197,G8982,G9298,G9299);
  nand GNAME9198(G9198,G9055,G9197);
  nand GNAME9199(G9199,G8983,G9301,G9302);
  nand GNAME9200(G9200,G9052,G9199);
  nand GNAME9201(G9201,G8984,G9304,G9305);
  nand GNAME9202(G9202,G9049,G9201);
  nand GNAME9203(G9203,G8985,G9307,G9308);
  nand GNAME9204(G9204,G9046,G9203);
  nand GNAME9205(G9205,G8986,G9310,G9311);
  nand GNAME9206(G9206,G9043,G9205);
  or GNAME9207(G9207,G3810,G9315);
  nand GNAME9208(G9208,G9040,G9207);
  not GNAME9209(G9209,G9039);
  nand GNAME9210(G9210,G9098,G9209);
  not GNAME9211(G9211,G9038);
  nand GNAME9212(G9212,G9070,G9118);
  nand GNAME9213(G9213,G9099,G9121);
  nand GNAME9214(G9214,G9213,G9112,G9212);
  nand GNAME9215(G9215,G9121,G8988);
  nand GNAME9216(G9216,G9101,G9170);
  nand GNAME9217(G9217,G9006,G9136);
  nand GNAME9218(G9218,G9217,G9135,G9216);
  nand GNAME9219(G9219,G9170,G8989);
  not GNAME9220(G9220,G9096);
  nand GNAME9221(G9221,G9104,G9105);
  nand GNAME9222(G9222,G9110,G9111);
  nand GNAME9223(G9223,G9098,G9103);
  nand GNAME9224(G9224,G9100,G9102);
  nand GNAME9225(G9225,G9164,G9165);
  or GNAME9226(G9226,G3800,G8956);
  or GNAME9227(G9227,G3776,G8998);
  or GNAME9228(G9228,G3802,G8956);
  or GNAME9229(G9229,G3776,G8999);
  nand GNAME9230(G9230,G9228,G9229);
  or GNAME9231(G9231,G3804,G8956);
  or GNAME9232(G9232,G3776,G9000);
  or GNAME9233(G9233,G3806,G8956);
  or GNAME9234(G9234,G3776,G9001);
  nand GNAME9235(G9235,G9233,G9234);
  or GNAME9236(G9236,G3807,G8956);
  or GNAME9237(G9237,G3776,G9002);
  nand GNAME9238(G9238,G9236,G9237);
  nand GNAME9239(G9239,G9231,G9232);
  or GNAME9240(G9240,G3803,G8956);
  or GNAME9241(G9241,G3776,G9003);
  nand GNAME9242(G9242,G9240,G9241);
  nand GNAME9243(G9243,G9226,G9227);
  or GNAME9244(G9244,G3799,G8956);
  or GNAME9245(G9245,G3776,G9004);
  nand GNAME9246(G9246,G9244,G9245);
  or GNAME9247(G9247,G3798,G8956);
  or GNAME9248(G9248,G3776,G9005);
  nand GNAME9249(G9249,G9247,G9248);
  or GNAME9250(G9250,G9007,G9006);
  nand GNAME9251(G9251,G9006,G9007);
  or GNAME9252(G9252,G9010,G9009);
  nand GNAME9253(G9253,G9009,G9010);
  nand GNAME9254(G9254,G9130,G9221);
  nand GNAME9255(G9255,G9012,G9104,G9105);
  or GNAME9256(G9256,G9014,G9013);
  nand GNAME9257(G9257,G9013,G9014);
  or GNAME9258(G9258,G9017,G9016);
  nand GNAME9259(G9259,G9016,G9017);
  nand GNAME9260(G9260,G9122,G9222);
  nand GNAME9261(G9261,G9019,G9110,G9111);
  or GNAME9262(G9262,G3796,G8956);
  or GNAME9263(G9263,G3776,G9020);
  nand GNAME9264(G9264,G9262,G9263);
  or GNAME9265(G9265,G3795,G8956);
  or GNAME9266(G9266,G3776,G9021);
  nand GNAME9267(G9267,G9265,G9266);
  or GNAME9268(G9268,G3794,G8956);
  or GNAME9269(G9269,G3776,G9022);
  nand GNAME9270(G9270,G9268,G9269);
  or GNAME9271(G9271,G3792,G8956);
  or GNAME9272(G9272,G3776,G9023);
  nand GNAME9273(G9273,G9271,G9272);
  or GNAME9274(G9274,G3791,G8956);
  or GNAME9275(G9275,G3776,G9024);
  nand GNAME9276(G9276,G9274,G9275);
  or GNAME9277(G9277,G3790,G8956);
  or GNAME9278(G9278,G3776,G9025);
  nand GNAME9279(G9279,G9277,G9278);
  or GNAME9280(G9280,G3789,G8956);
  or GNAME9281(G9281,G3776,G9026);
  nand GNAME9282(G9282,G9280,G9281);
  or GNAME9283(G9283,G3788,G8956);
  or GNAME9284(G9284,G3776,G9027);
  nand GNAME9285(G9285,G9283,G9284);
  or GNAME9286(G9286,G3787,G8956);
  or GNAME9287(G9287,G3776,G9028);
  nand GNAME9288(G9288,G9286,G9287);
  or GNAME9289(G9289,G3786,G8956);
  or GNAME9290(G9290,G3776,G9029);
  nand GNAME9291(G9291,G9289,G9290);
  or GNAME9292(G9292,G3785,G8956);
  or GNAME9293(G9293,G3776,G9030);
  nand GNAME9294(G9294,G9292,G9293);
  or GNAME9295(G9295,G3784,G8956);
  or GNAME9296(G9296,G3776,G9031);
  nand GNAME9297(G9297,G9295,G9296);
  or GNAME9298(G9298,G3783,G8956);
  or GNAME9299(G9299,G3776,G9032);
  nand GNAME9300(G9300,G9298,G9299);
  or GNAME9301(G9301,G3782,G8956);
  or GNAME9302(G9302,G3776,G9033);
  nand GNAME9303(G9303,G9301,G9302);
  or GNAME9304(G9304,G3781,G8956);
  or GNAME9305(G9305,G3776,G9034);
  nand GNAME9306(G9306,G9304,G9305);
  or GNAME9307(G9307,G3780,G8956);
  or GNAME9308(G9308,G3776,G9035);
  nand GNAME9309(G9309,G9307,G9308);
  or GNAME9310(G9310,G3779,G8956);
  or GNAME9311(G9311,G3776,G9036);
  nand GNAME9312(G9312,G9310,G9311);
  or GNAME9313(G9313,G3778,G8956);
  nand GNAME9314(G9314,G8956,G3778);
  not GNAME9315(G9315,G8990);
  or GNAME9316(G9316,G9038,G9037);
  or GNAME9317(G9317,G3808,G9211);
  nand GNAME9318(G9318,G9316,G9317);
  nand GNAME9319(G9319,G8990,G9316,G9317);
  nand GNAME9320(G9320,G9315,G9318);
  nand GNAME9321(G9321,G9209,G9223);
  nand GNAME9322(G9322,G9039,G9098,G9103);
  or GNAME9323(G9323,G9041,G9040);
  nand GNAME9324(G9324,G9040,G9041);
  or GNAME9325(G9325,G9044,G9043);
  nand GNAME9326(G9326,G9043,G9044);
  or GNAME9327(G9327,G9047,G9046);
  nand GNAME9328(G9328,G9046,G9047);
  or GNAME9329(G9329,G9050,G9049);
  nand GNAME9330(G9330,G9049,G9050);
  or GNAME9331(G9331,G9053,G9052);
  nand GNAME9332(G9332,G9052,G9053);
  or GNAME9333(G9333,G9056,G9055);
  nand GNAME9334(G9334,G9055,G9056);
  or GNAME9335(G9335,G9059,G9058);
  nand GNAME9336(G9336,G9058,G9059);
  or GNAME9337(G9337,G9062,G9061);
  nand GNAME9338(G9338,G9061,G9062);
  or GNAME9339(G9339,G9065,G9064);
  nand GNAME9340(G9340,G9064,G9065);
  or GNAME9341(G9341,G9068,G9067);
  nand GNAME9342(G9342,G9067,G9068);
  or GNAME9343(G9343,G9071,G9070);
  nand GNAME9344(G9344,G9070,G9071);
  or GNAME9345(G9345,G9074,G9073);
  nand GNAME9346(G9346,G9073,G9074);
  or GNAME9347(G9347,G9077,G9076);
  nand GNAME9348(G9348,G9076,G9077);
  or GNAME9349(G9349,G9080,G9079);
  nand GNAME9350(G9350,G9079,G9080);
  or GNAME9351(G9351,G9083,G9082);
  nand GNAME9352(G9352,G9082,G9083);
  or GNAME9353(G9353,G9086,G9085);
  nand GNAME9354(G9354,G9085,G9086);
  nand GNAME9355(G9355,G9177,G9224);
  nand GNAME9356(G9356,G9088,G9100,G9102);
  or GNAME9357(G9357,G9090,G9089);
  nand GNAME9358(G9358,G9089,G9090);
  or GNAME9359(G9359,G9093,G9092);
  nand GNAME9360(G9360,G9092,G9093);
  nand GNAME9361(G9361,G9171,G9225);
  nand GNAME9362(G9362,G9095,G9164,G9165);
  or GNAME9363(G9363,G9096,G8956);
  or GNAME9364(G9364,G3776,G9220);
  not GNAME9365(G9365,G9121);
  not GNAME9366(G9366,G9129);
  not GNAME9367(G9367,G9170);
  not GNAME9368(G9368,G3683);
  and GNAME9369(G9369,G9370,G9371);
  or GNAME9370(G9370,G9368,G3681);
  nand GNAME9371(G9371,G9368,G3681);
  nand GNAME9372(G9372,G6384,G9417);
  nand GNAME9373(G9373,G6377,G9410);
  nand GNAME9374(G9374,G6392,G9400);
  nand GNAME9375(G9375,G6372,G9405);
  nand GNAME9376(G9376,G6385,G9418);
  nand GNAME9377(G9377,G6379,G9412);
  nand GNAME9378(G9378,G6394,G9402);
  nand GNAME9379(G9379,G6371,G9404);
  nand GNAME9380(G9380,G6395,G9403);
  nand GNAME9381(G9381,G6380,G9413);
  nand GNAME9382(G9382,G6386,G9419);
  nand GNAME9383(G9383,G6383,G9416);
  nand GNAME9384(G9384,G6393,G9401);
  nand GNAME9385(G9385,G6378,G9411);
  nand GNAME9386(G9386,G6381,G9414);
  nand GNAME9387(G9387,G6376,G9409);
  nand GNAME9388(G9388,G6391,G9399);
  nand GNAME9389(G9389,G6388,G6397);
  nand GNAME9390(G9390,G6373,G9406);
  nand GNAME9391(G9391,G6374,G9407);
  not GNAME9392(G9392,G23037);
  nand GNAME9393(G9393,G6387,G6398);
  nand GNAME9394(G9394,G6382,G9415);
  or GNAME9395(G9395,G6389,G6396);
  nand GNAME9396(G9396,G6390,G9398);
  nand GNAME9397(G9397,G6375,G9408);
  or GNAME9398(G9398,G23037,G23025);
  or GNAME9399(G9399,G23028,G9398);
  or GNAME9400(G9400,G23016,G9399);
  or GNAME9401(G9401,G23042,G9400);
  or GNAME9402(G9402,G23034,G9401);
  or GNAME9403(G9403,G23024,G9402);
  or GNAME9404(G9404,G23038,G9403);
  or GNAME9405(G9405,G23019,G9404);
  or GNAME9406(G9406,G23031,G9405);
  or GNAME9407(G9407,G23021,G9406);
  or GNAME9408(G9408,G23040,G9407);
  or GNAME9409(G9409,G23014,G9408);
  or GNAME9410(G9410,G23029,G9409);
  or GNAME9411(G9411,G23027,G9410);
  or GNAME9412(G9412,G23017,G9411);
  or GNAME9413(G9413,G23036,G9412);
  or GNAME9414(G9414,G23022,G9413);
  or GNAME9415(G9415,G23032,G9414);
  or GNAME9416(G9416,G23020,G9415);
  or GNAME9417(G9417,G23039,G9416);
  or GNAME9418(G9418,G23026,G9417);
  or GNAME9419(G9419,G23030,G9418);

endmodule