module b22s(CK,G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G10148,G10226,G10228,G10230,G10232,G10234,G10236,G10238,G10240,G10242,G10208,G10210,G10212,G10214,G10216,G10218,G10220,G10222,G10188,G10149,G792,G793);
input CK,G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32;
output G10148,G10226,G10228,G10230,G10232,G10234,G10236,G10238,G10240,G10242,G10208,G10210,G10212,G10214,G10216,G10218,G10220,G10222,G10188,G10149,G792,G793;

  wire G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,
       G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,G40,
       G41,G42,G43,G44,G45,G46,G47,G48,G49,G50,G51,G52,G53,G54,G55,G56,G57,G58,G59,G60,
       G61,G62,G63,G64,G65,G66,G67,G68,G69,G70,G71,G72,G73,G74,G75,G76,G77,G78,G79,G80,
       G81,G82,G83,G84,G85,G86,G87,G88,G89,G90,G91,G92,G93,G94,G95,G96,G97,G98,G99,G100,
       G101,G102,G103,G104,G105,G106,G107,G108,G109,G110,G111,G112,G113,G114,G115,G116,G117,G118,G119,G120,
       G121,G122,G123,G124,G125,G126,G127,G128,G129,G130,G131,G132,G133,G134,G135,G136,G137,G138,G139,G140,
       G141,G142,G143,G144,G145,G146,G147,G148,G149,G150,G151,G152,G153,G154,G155,G156,G157,G158,G159,G160,
       G161,G162,G163,G164,G165,G166,G167,G168,G169,G170,G171,G172,G173,G174,G175,G176,G177,G178,G179,G180,
       G181,G182,G183,G184,G185,G186,G187,G188,G189,G190,G191,G192,G193,G194,G195,G196,G197,G198,G199,G200,
       G201,G202,G203,G204,G205,G206,G207,G208,G209,G210,G211,G212,G213,G214,G215,G216,G217,G218,G219,G220,
       G221,G222,G223,G224,G225,G226,G227,G228,G229,G230,G231,G232,G233,G234,G235,G236,G237,G238,G239,G240,
       G241,G242,G243,G244,G245,G246,G247,G248,G249,G250,G251,G252,G253,G254,G255,G256,G257,G258,G259,G260,
       G261,G262,G263,G264,G265,G266,G267,G268,G269,G270,G271,G272,G273,G274,G275,G276,G277,G278,G279,G280,
       G281,G282,G283,G284,G285,G286,G287,G288,G289,G290,G291,G292,G293,G294,G295,G296,G297,G298,G299,G300,
       G301,G302,G303,G304,G305,G306,G307,G308,G309,G310,G311,G312,G313,G314,G315,G316,G317,G318,G319,G320,
       G321,G322,G323,G324,G325,G326,G327,G328,G329,G330,G331,G332,G333,G334,G335,G336,G337,G338,G339,G340,
       G341,G342,G343,G344,G345,G346,G347,G348,G349,G350,G351,G352,G353,G354,G355,G356,G357,G358,G359,G360,
       G361,G362,G363,G364,G365,G366,G367,G368,G369,G370,G371,G372,G373,G374,G375,G376,G377,G378,G379,G380,
       G381,G382,G383,G384,G385,G386,G387,G388,G389,G390,G391,G392,G393,G394,G395,G396,G397,G398,G399,G400,
       G401,G402,G403,G404,G405,G406,G407,G408,G409,G410,G411,G412,G413,G414,G415,G416,G417,G418,G419,G420,
       G421,G422,G423,G424,G425,G426,G427,G428,G429,G430,G431,G432,G433,G434,G435,G436,G437,G438,G439,G440,
       G441,G442,G443,G444,G445,G446,G447,G448,G449,G450,G451,G452,G453,G454,G455,G456,G457,G458,G459,G460,
       G461,G462,G463,G464,G465,G466,G467,G468,G469,G470,G471,G472,G473,G474,G475,G476,G477,G478,G479,G480,
       G481,G482,G483,G484,G485,G486,G487,G488,G489,G490,G491,G492,G493,G494,G495,G496,G497,G498,G499,G500,
       G501,G502,G503,G504,G505,G506,G507,G508,G509,G510,G511,G512,G513,G514,G515,G516,G517,G518,G519,G520,
       G521,G522,G523,G524,G525,G526,G527,G528,G529,G530,G531,G532,G533,G534,G535,G536,G537,G538,G539,G540,
       G541,G542,G543,G544,G545,G546,G547,G548,G549,G550,G551,G552,G553,G554,G555,G556,G557,G558,G559,G560,
       G561,G562,G563,G564,G565,G566,G567,G568,G569,G570,G571,G572,G573,G574,G575,G576,G577,G578,G579,G580,
       G581,G582,G583,G584,G585,G586,G587,G588,G589,G590,G591,G592,G593,G594,G595,G596,G597,G598,G599,G600,
       G601,G602,G603,G604,G605,G606,G607,G608,G609,G610,G611,G612,G613,G614,G615,G616,G617,G618,G619,G620,
       G621,G622,G623,G624,G625,G626,G627,G628,G629,G630,G631,G632,G633,G634,G635,G636,G637,G638,G639,G640,
       G641,G642,G643,G644,G645,G646,G647,G648,G649,G650,G651,G652,G653,G654,G655,G656,G657,G658,G659,G660,
       G661,G662,G663,G664,G665,G666,G667,G668,G669,G670,G671,G672,G673,G674,G675,G676,G677,G678,G679,G680,
       G681,G682,G683,G684,G685,G686,G687,G688,G689,G690,G691,G692,G693,G694,G695,G696,G697,G698,G699,G700,
       G701,G702,G703,G704,G705,G706,G707,G708,G709,G710,G711,G712,G713,G714,G715,G716,G717,G718,G719,G720,
       G721,G722,G723,G724,G725,G726,G727,G728,G729,G730,G731,G732,G733,G734,G735,G736,G737,G738,G739,G740,
       G741,G742,G743,G744,G745,G746,G747,G748,G749,G750,G751,G752,G753,G754,G755,G756,G757,G758,G759,G760,
       G761,G762,G763,G764,G765,G766,G767,G768,G769,G770,G771,G772,G773,G774,G775,G776,G777,G778,G779,G780,
       G781,G782,G783,G784,G785,G786,G787,G788,G789,G790,G791,G792,G793,G794,G795,G796,G797,G798,G799,G800,
       G801,G802,G803,G804,G805,G806,G807,G808,G809,G810,G811,G812,G813,G814,G815,G816,G817,G818,G819,G820,
       G821,G822,G823,G824,G825,G826,G827,G828,G829,G830,G831,G832,G833,G834,G835,G836,G837,G838,G839,G840,
       G841,G842,G843,G844,G845,G846,G847,G848,G849,G850,G851,G852,G853,G854,G855,G856,G857,G858,G859,G860,
       G861,G862,G863,G864,G865,G866,G867,G868,G869,G870,G871,G872,G873,G874,G875,G876,G877,G878,G879,G880,
       G881,G882,G883,G884,G885,G886,G887,G888,G889,G890,G891,G892,G893,G894,G895,G896,G897,G898,G899,G900,
       G901,G902,G903,G904,G905,G906,G907,G908,G909,G910,G911,G912,G913,G914,G915,G916,G917,G918,G919,G920,
       G921,G922,G923,G924,G925,G926,G927,G928,G929,G930,G931,G932,G933,G934,G935,G936,G937,G938,G939,G940,
       G941,G942,G943,G944,G945,G946,G947,G948,G949,G950,G951,G952,G953,G954,G955,G956,G957,G958,G959,G960,
       G961,G962,G963,G964,G965,G966,G967,G968,G969,G970,G971,G972,G973,G974,G975,G976,G977,G978,G979,G980,
       G981,G982,G983,G984,G985,G986,G987,G988,G989,G990,G991,G992,G993,G994,G995,G996,G997,G998,G999,G1000,
       G1001,G1002,G1003,G1004,G1005,G1006,G1007,G1008,G1009,G1010,G1011,G1012,G1013,G1014,G1015,G1016,G1017,G1018,G1019,G1020,
       G1021,G1022,G1023,G1024,G1025,G1026,G1027,G1028,G1029,G1030,G1031,G1032,G1033,G1034,G1035,G1036,G1037,G1038,G1039,G1040,
       G1041,G1042,G1043,G1044,G1045,G1046,G1047,G1048,G1049,G1050,G1051,G1052,G1053,G1054,G1055,G1056,G1057,G1058,G1059,G1060,
       G1061,G1062,G1063,G1064,G1065,G1066,G1067,G1068,G1069,G1070,G1071,G1072,G1073,G1074,G1075,G1076,G1077,G1078,G1079,G1080,
       G1081,G1082,G1083,G1084,G1085,G1086,G1087,G1088,G1089,G1090,G1091,G1092,G1093,G1094,G1095,G1096,G1097,G1098,G1099,G1100,
       G1101,G1102,G1103,G1104,G1105,G1106,G1107,G1108,G1109,G1110,G1111,G1112,G1113,G1114,G1115,G1116,G1117,G1118,G1119,G1120,
       G1121,G1122,G1123,G1124,G1125,G1126,G1127,G1128,G1129,G1130,G1131,G1132,G1133,G1134,G1135,G1136,G1137,G1138,G1139,G1140,
       G1141,G1142,G1143,G1144,G1145,G1146,G1147,G1148,G1149,G1150,G1151,G1152,G1153,G1154,G1155,G1156,G1157,G1158,G1159,G1160,
       G1161,G1162,G1163,G1164,G1165,G1166,G1167,G1168,G1169,G1170,G1171,G1172,G1173,G1174,G1175,G1176,G1177,G1178,G1179,G1180,
       G1181,G1182,G1183,G1184,G1185,G1186,G1187,G1188,G1189,G1190,G1191,G1192,G1193,G1194,G1195,G1196,G1197,G1198,G1199,G1200,
       G1201,G1202,G1203,G1204,G1205,G1206,G1207,G1208,G1209,G1210,G1211,G1212,G1213,G1214,G1215,G1216,G1217,G1218,G1219,G1220,
       G1221,G1222,G1223,G1224,G1225,G1226,G1227,G1228,G1229,G1230,G1231,G1232,G1233,G1234,G1235,G1236,G1237,G1238,G1239,G1240,
       G1241,G1242,G1243,G1244,G1245,G1246,G1247,G1248,G1249,G1250,G1251,G1252,G1253,G1254,G1255,G1256,G1257,G1258,G1259,G1260,
       G1261,G1262,G1263,G1264,G1265,G1266,G1267,G1268,G1269,G1270,G1271,G1272,G1273,G1274,G1275,G1276,G1277,G1278,G1279,G1280,
       G1281,G1282,G1283,G1284,G1285,G1286,G1287,G1288,G1289,G1290,G1291,G1292,G1293,G1294,G1295,G1296,G1297,G1298,G1299,G1300,
       G1301,G1302,G1303,G1304,G1305,G1306,G1307,G1308,G1309,G1310,G1311,G1312,G1313,G1314,G1315,G1316,G1317,G1318,G1319,G1320,
       G1321,G1322,G1323,G1324,G1325,G1326,G1327,G1328,G1329,G1330,G1331,G1332,G1333,G1334,G1335,G1336,G1337,G1338,G1339,G1340,
       G1341,G1342,G1343,G1344,G1345,G1346,G1347,G1348,G1349,G1350,G1351,G1352,G1353,G1354,G1355,G1356,G1357,G1358,G1359,G1360,
       G1361,G1362,G1363,G1364,G1365,G1366,G1367,G1368,G1369,G1370,G1371,G1372,G1373,G1374,G1375,G1376,G1377,G1378,G1379,G1380,
       G1381,G1382,G1383,G1384,G1385,G1386,G1387,G1388,G1389,G1390,G1391,G1392,G1393,G1394,G1395,G1396,G1397,G1398,G1399,G1400,
       G1401,G1402,G1403,G1404,G1405,G1406,G1407,G1408,G1409,G1410,G1411,G1412,G1413,G1414,G1415,G1416,G1417,G1418,G1419,G1420,
       G1421,G1422,G1423,G1424,G1425,G1426,G1427,G1428,G1429,G1430,G1431,G1432,G1433,G1434,G1435,G1436,G1437,G1438,G1439,G1440,
       G1441,G1442,G1443,G1444,G1445,G1446,G1447,G1448,G1449,G1450,G1451,G1452,G1453,G1454,G1455,G1456,G1457,G1458,G1459,G1460,
       G1461,G1462,G1463,G1464,G1465,G1466,G1467,G1468,G1469,G1470,G1471,G1472,G1473,G1474,G1475,G1476,G1477,G1478,G1479,G1480,
       G1481,G1482,G1483,G1484,G1485,G1486,G1487,G1488,G1489,G1490,G1491,G1492,G1493,G1494,G1495,G1496,G1497,G1498,G1499,G1500,
       G1501,G1502,G1503,G1504,G1505,G1506,G1507,G1508,G1509,G1510,G1511,G1512,G1513,G1514,G1515,G1516,G1517,G1518,G1519,G1520,
       G1521,G1522,G1523,G1524,G1525,G1526,G1527,G1528,G1529,G1530,G1531,G1532,G1533,G1534,G1535,G1536,G1537,G1538,G1539,G1540,
       G1541,G1542,G1543,G1544,G1545,G1546,G1547,G1548,G1549,G1550,G1551,G1552,G1553,G1554,G1555,G1556,G1557,G1558,G1559,G1560,
       G1561,G1562,G1563,G1564,G1565,G1566,G1567,G1568,G1569,G1570,G1571,G1572,G1573,G1574,G1575,G1576,G1577,G1578,G1579,G1580,
       G1581,G1582,G1583,G1584,G1585,G1586,G1587,G1588,G1589,G1590,G1591,G1592,G1593,G1594,G1595,G1596,G1597,G1598,G1599,G1600,
       G1601,G1602,G1603,G1604,G1605,G1606,G1607,G1608,G1609,G1610,G1611,G1612,G1613,G1614,G1615,G1616,G1617,G1618,G1619,G1620,
       G1621,G1622,G1623,G1624,G1625,G1626,G1627,G1628,G1629,G1630,G1631,G1632,G1633,G1634,G1635,G1636,G1637,G1638,G1639,G1640,
       G1641,G1642,G1643,G1644,G1645,G1646,G1647,G1648,G1649,G1650,G1651,G1652,G1653,G1654,G1655,G1656,G1657,G1658,G1659,G1660,
       G1661,G1662,G1663,G1664,G1665,G1666,G1667,G1668,G1669,G1670,G1671,G1672,G1673,G1674,G1675,G1676,G1677,G1678,G1679,G1680,
       G1681,G1682,G1683,G1684,G1685,G1686,G1687,G1688,G1689,G1690,G1691,G1692,G1693,G1694,G1695,G1696,G1697,G1698,G1699,G1700,
       G1701,G1702,G1703,G1704,G1705,G1706,G1707,G1708,G1709,G1710,G1711,G1712,G1713,G1714,G1715,G1716,G1717,G1718,G1719,G1720,
       G1721,G1722,G1723,G1724,G1725,G1726,G1727,G1728,G1729,G1730,G1731,G1732,G1733,G1734,G1735,G1736,G1737,G1738,G1739,G1740,
       G1741,G1742,G1743,G1744,G1745,G1746,G1747,G1748,G1749,G1750,G1751,G1752,G1753,G1754,G1755,G1756,G1757,G1758,G1759,G1760,
       G1761,G1762,G1763,G1764,G1765,G1766,G1767,G1768,G1769,G1770,G1771,G1772,G1773,G1774,G1775,G1776,G1777,G1778,G1779,G1780,
       G1781,G1782,G1783,G1784,G1785,G1786,G1787,G1788,G1789,G1790,G1791,G1792,G1793,G1794,G1795,G1796,G1797,G1798,G1799,G1800,
       G1801,G1802,G1803,G1804,G1805,G1806,G1807,G1808,G1809,G1810,G1811,G1812,G1813,G1814,G1815,G1816,G1817,G1818,G1819,G1820,
       G1821,G1822,G1823,G1824,G1825,G1826,G1827,G1828,G1829,G1830,G1831,G1832,G1833,G1834,G1835,G1836,G1837,G1838,G1839,G1840,
       G1841,G1842,G1843,G1844,G1845,G1846,G1847,G1848,G1849,G1850,G1851,G1852,G1853,G1854,G1855,G1856,G1857,G1858,G1859,G1860,
       G1861,G1862,G1863,G1864,G1865,G1866,G1867,G1868,G1869,G1870,G1871,G1872,G1873,G1874,G1875,G1876,G1877,G1878,G1879,G1880,
       G1881,G1882,G1883,G1884,G1885,G1886,G1887,G1888,G1889,G1890,G1891,G1892,G1893,G1894,G1895,G1896,G1897,G1898,G1899,G1900,
       G1901,G1902,G1903,G1904,G1905,G1906,G1907,G1908,G1909,G1910,G1911,G1912,G1913,G1914,G1915,G1916,G1917,G1918,G1919,G1920,
       G1921,G1922,G1923,G1924,G1925,G1926,G1927,G1928,G1929,G1930,G1931,G1932,G1933,G1934,G1935,G1936,G1937,G1938,G1939,G1940,
       G1941,G1942,G1943,G1944,G1945,G1946,G1947,G1948,G1949,G1950,G1951,G1952,G1953,G1954,G1955,G1956,G1957,G1958,G1959,G1960,
       G1961,G1962,G1963,G1964,G1965,G1966,G1967,G1968,G1969,G1970,G1971,G1972,G1973,G1974,G1975,G1976,G1977,G1978,G1979,G1980,
       G1981,G1982,G1983,G1984,G1985,G1986,G1987,G1988,G1989,G1990,G1991,G1992,G1993,G1994,G1995,G1996,G1997,G1998,G1999,G2000,
       G2001,G2002,G2003,G2004,G2005,G2006,G2007,G2008,G2009,G2010,G2011,G2012,G2013,G2014,G2015,G2016,G2017,G2018,G2019,G2020,
       G2021,G2022,G2023,G2024,G2025,G2026,G2027,G2028,G2029,G2030,G2031,G2032,G2033,G2034,G2035,G2036,G2037,G2038,G2039,G2040,
       G2041,G2042,G2043,G2044,G2045,G2046,G2047,G2048,G2049,G2050,G2051,G2052,G2053,G2054,G2055,G2056,G2057,G2058,G2059,G2060,
       G2061,G2062,G2063,G2064,G2065,G2066,G2067,G2068,G2069,G2070,G2071,G2072,G2073,G2074,G2075,G2076,G2077,G2078,G2079,G2080,
       G2081,G2082,G2083,G2084,G2085,G2086,G2087,G2088,G2089,G2090,G2091,G2092,G2093,G2094,G2095,G2096,G2097,G2098,G2099,G2100,
       G2101,G2102,G2103,G2104,G2105,G2106,G2107,G2108,G2109,G2110,G2111,G2112,G2113,G2114,G2115,G2116,G2117,G2118,G2119,G2120,
       G2121,G2122,G2123,G2124,G2125,G2126,G2127,G2128,G2129,G2130,G2131,G2132,G2133,G2134,G2135,G2136,G2137,G2138,G2139,G2140,
       G2141,G2142,G2143,G2144,G2145,G2146,G2147,G2148,G2149,G2150,G2151,G2152,G2153,G2154,G2155,G2156,G2157,G2158,G2159,G2160,
       G2161,G2162,G2163,G2164,G2165,G2166,G2167,G2168,G2169,G2170,G2171,G2172,G2173,G2174,G2175,G2176,G2177,G2178,G2179,G2180,
       G2181,G2182,G2183,G2184,G2185,G2186,G2187,G2188,G2189,G2190,G2191,G2192,G2193,G2194,G2195,G2196,G2197,G2198,G2199,G2200,
       G2201,G2202,G2203,G2204,G2205,G2206,G2207,G2208,G2209,G2210,G2211,G2212,G2213,G2214,G2215,G2216,G2217,G2218,G2219,G2220,
       G2221,G2222,G2223,G2224,G2225,G2226,G2227,G2228,G2229,G2230,G2231,G2232,G2233,G2234,G2235,G2236,G2237,G2238,G2239,G2240,
       G2241,G2242,G2243,G2244,G2245,G2246,G2247,G2248,G2249,G2250,G2251,G2252,G2253,G2254,G2255,G2256,G2257,G2258,G2259,G2260,
       G2261,G2262,G2263,G2264,G2265,G2266,G2267,G2268,G2269,G2270,G2271,G2272,G2273,G2274,G2275,G2276,G2277,G2278,G2279,G2280,
       G2281,G2282,G2283,G2284,G2285,G2286,G2287,G2288,G2289,G2290,G2291,G2292,G2293,G2294,G2295,G2296,G2297,G2298,G2299,G2300,
       G2301,G2302,G2303,G2304,G2305,G2306,G2307,G2308,G2309,G2310,G2311,G2312,G2313,G2314,G2315,G2316,G2317,G2318,G2319,G2320,
       G2321,G2322,G2323,G2324,G2325,G2326,G2327,G2328,G2329,G2330,G2331,G2332,G2333,G2334,G2335,G2336,G2337,G2338,G2339,G2340,
       G2341,G2342,G2343,G2344,G2345,G2346,G2347,G2348,G2349,G2350,G2351,G2352,G2353,G2354,G2355,G2356,G2357,G2358,G2359,G2360,
       G2361,G2362,G2363,G2364,G2365,G2366,G2367,G2368,G2369,G2370,G2371,G2372,G2373,G2374,G2375,G2376,G2377,G2378,G2379,G2380,
       G2381,G2382,G2383,G2384,G2385,G2386,G2387,G2388,G2389,G2390,G2391,G2392,G2393,G2394,G2395,G2396,G2397,G2398,G2399,G2400,
       G2401,G2402,G2403,G2404,G2405,G2406,G2407,G2408,G2409,G2410,G2411,G2412,G2413,G2414,G2415,G2416,G2417,G2418,G2419,G2420,
       G2421,G2422,G2423,G2424,G2425,G2426,G2427,G2428,G2429,G2430,G2431,G2432,G2433,G2434,G2435,G2436,G2437,G2438,G2439,G2440,
       G2441,G2442,G2443,G2444,G2445,G2446,G2447,G2448,G2449,G2450,G2451,G2452,G2453,G2454,G2455,G2456,G2457,G2458,G2459,G2460,
       G2461,G2462,G2463,G2464,G2465,G2466,G2467,G2468,G2469,G2470,G2471,G2472,G2473,G2474,G2475,G2476,G2477,G2478,G2479,G2480,
       G2481,G2482,G2483,G2484,G2485,G2486,G2487,G2488,G2489,G2490,G2491,G2492,G2493,G2494,G2495,G2496,G2497,G2498,G2499,G2500,
       G2501,G2502,G2503,G2504,G2505,G2506,G2507,G2508,G2509,G2510,G2511,G2512,G2513,G2514,G2515,G2516,G2517,G2518,G2519,G2520,
       G2521,G2522,G2523,G2524,G2525,G2526,G2527,G2528,G2529,G2530,G2531,G2532,G2533,G2534,G2535,G2536,G2537,G2538,G2539,G2540,
       G2541,G2542,G2543,G2544,G2545,G2546,G2547,G2548,G2549,G2550,G2551,G2552,G2553,G2554,G2555,G2556,G2557,G2558,G2559,G2560,
       G2561,G2562,G2563,G2564,G2565,G2566,G2567,G2568,G2569,G2570,G2571,G2572,G2573,G2574,G2575,G2576,G2577,G2578,G2579,G2580,
       G2581,G2582,G2583,G2584,G2585,G2586,G2587,G2588,G2589,G2590,G2591,G2592,G2593,G2594,G2595,G2596,G2597,G2598,G2599,G2600,
       G2601,G2602,G2603,G2604,G2605,G2606,G2607,G2608,G2609,G2610,G2611,G2612,G2613,G2614,G2615,G2616,G2617,G2618,G2619,G2620,
       G2621,G2622,G2623,G2624,G2625,G2626,G2627,G2628,G2629,G2630,G2631,G2632,G2633,G2634,G2635,G2636,G2637,G2638,G2639,G2640,
       G2641,G2642,G2643,G2644,G2645,G2646,G2647,G2648,G2649,G2650,G2651,G2652,G2653,G2654,G2655,G2656,G2657,G2658,G2659,G2660,
       G2661,G2662,G2663,G2664,G2665,G2666,G2667,G2668,G2669,G2670,G2671,G2672,G2673,G2674,G2675,G2676,G2677,G2678,G2679,G2680,
       G2681,G2682,G2683,G2684,G2685,G2686,G2687,G2688,G2689,G2690,G2691,G2692,G2693,G2694,G2695,G2696,G2697,G2698,G2699,G2700,
       G2701,G2702,G2703,G2704,G2705,G2706,G2707,G2708,G2709,G2710,G2711,G2712,G2713,G2714,G2715,G2716,G2717,G2718,G2719,G2720,
       G2721,G2722,G2723,G2724,G2725,G2726,G2727,G2728,G2729,G2730,G2731,G2732,G2733,G2734,G2735,G2736,G2737,G2738,G2739,G2740,
       G2741,G2742,G2743,G2744,G2745,G2746,G2747,G2748,G2749,G2750,G2751,G2752,G2753,G2754,G2755,G2756,G2757,G2758,G2759,G2760,
       G2761,G2762,G2763,G2764,G2765,G2766,G2767,G2768,G2769,G2770,G2771,G2772,G2773,G2774,G2775,G2776,G2777,G2778,G2779,G2780,
       G2781,G2782,G2783,G2784,G2785,G2786,G2787,G2788,G2789,G2790,G2791,G2792,G2793,G2794,G2795,G2796,G2797,G2798,G2799,G2800,
       G2801,G2802,G2803,G2804,G2805,G2806,G2807,G2808,G2809,G2810,G2811,G2812,G2813,G2814,G2815,G2816,G2817,G2818,G2819,G2820,
       G2821,G2822,G2823,G2824,G2825,G2826,G2827,G2828,G2829,G2830,G2831,G2832,G2833,G2834,G2835,G2836,G2837,G2838,G2839,G2840,
       G2841,G2842,G2843,G2844,G2845,G2846,G2847,G2848,G2849,G2850,G2851,G2852,G2853,G2854,G2855,G2856,G2857,G2858,G2859,G2860,
       G2861,G2862,G2863,G2864,G2865,G2866,G2867,G2868,G2869,G2870,G2871,G2872,G2873,G2874,G2875,G2876,G2877,G2878,G2879,G2880,
       G2881,G2882,G2883,G2884,G2885,G2886,G2887,G2888,G2889,G2890,G2891,G2892,G2893,G2894,G2895,G2896,G2897,G2898,G2899,G2900,
       G2901,G2902,G2903,G2904,G2905,G2906,G2907,G2908,G2909,G2910,G2911,G2912,G2913,G2914,G2915,G2916,G2917,G2918,G2919,G2920,
       G2921,G2922,G2923,G2924,G2925,G2926,G2927,G2928,G2929,G2930,G2931,G2932,G2933,G2934,G2935,G2936,G2937,G2938,G2939,G2940,
       G2941,G2942,G2943,G2944,G2945,G2946,G2947,G2948,G2949,G2950,G2951,G2952,G2953,G2954,G2955,G2956,G2957,G2958,G2959,G2960,
       G2961,G2962,G2963,G2964,G2965,G2966,G2967,G2968,G2969,G2970,G2971,G2972,G2973,G2974,G2975,G2976,G2977,G2978,G2979,G2980,
       G2981,G2982,G2983,G2984,G2985,G2986,G2987,G2988,G2989,G2990,G2991,G2992,G2993,G2994,G2995,G2996,G2997,G2998,G2999,G3000,
       G3001,G3002,G3003,G3004,G3005,G3006,G3007,G3008,G3009,G3010,G3011,G3012,G3013,G3014,G3015,G3016,G3017,G3018,G3019,G3020,
       G3021,G3022,G3023,G3024,G3025,G3026,G3027,G3028,G3029,G3030,G3031,G3032,G3033,G3034,G3035,G3036,G3037,G3038,G3039,G3040,
       G3041,G3042,G3043,G3044,G3045,G3046,G3047,G3048,G3049,G3050,G3051,G3052,G3053,G3054,G3055,G3056,G3057,G3058,G3059,G3060,
       G3061,G3062,G3063,G3064,G3065,G3066,G3067,G3068,G3069,G3070,G3071,G3072,G3073,G3074,G3075,G3076,G3077,G3078,G3079,G3080,
       G3081,G3082,G3083,G3084,G3085,G3086,G3087,G3088,G3089,G3090,G3091,G3092,G3093,G3094,G3095,G3096,G3097,G3098,G3099,G3100,
       G3101,G3102,G3103,G3104,G3105,G3106,G3107,G3108,G3109,G3110,G3111,G3112,G3113,G3114,G3115,G3116,G3117,G3118,G3119,G3120,
       G3121,G3122,G3123,G3124,G3125,G3126,G3127,G3128,G3129,G3130,G3131,G3132,G3133,G3134,G3135,G3136,G3137,G3138,G3139,G3140,
       G3141,G3142,G3143,G3144,G3145,G3146,G3147,G3148,G3149,G3150,G3151,G3152,G3153,G3154,G3155,G3156,G3157,G3158,G3159,G3160,
       G3161,G3162,G3163,G3164,G3165,G3166,G3167,G3168,G3169,G3170,G3171,G3172,G3173,G3174,G3175,G3176,G3177,G3178,G3179,G3180,
       G3181,G3182,G3183,G3184,G3185,G3186,G3187,G3188,G3189,G3190,G3191,G3192,G3193,G3194,G3195,G3196,G3197,G3198,G3199,G3200,
       G3201,G3202,G3203,G3204,G3205,G3206,G3207,G3208,G3209,G3210,G3211,G3212,G3213,G3214,G3215,G3216,G3217,G3218,G3219,G3220,
       G3221,G3222,G3223,G3224,G3225,G3226,G3227,G3228,G3229,G3230,G3231,G3232,G3233,G3234,G3235,G3236,G3237,G3238,G3239,G3240,
       G3241,G3242,G3243,G3244,G3245,G3246,G3247,G3248,G3249,G3250,G3251,G3252,G3253,G3254,G3255,G3256,G3257,G3258,G3259,G3260,
       G3261,G3262,G3263,G3264,G3265,G3266,G3267,G3268,G3269,G3270,G3271,G3272,G3273,G3274,G3275,G3276,G3277,G3278,G3279,G3280,
       G3281,G3282,G3283,G3284,G3285,G3286,G3287,G3288,G3289,G3290,G3291,G3292,G3293,G3294,G3295,G3296,G3297,G3298,G3299,G3300,
       G3301,G3302,G3303,G3304,G3305,G3306,G3307,G3308,G3309,G3310,G3311,G3312,G3313,G3314,G3315,G3316,G3317,G3318,G3319,G3320,
       G3321,G3322,G3323,G3324,G3325,G3326,G3327,G3328,G3329,G3330,G3331,G3332,G3333,G3334,G3335,G3336,G3337,G3338,G3339,G3340,
       G3341,G3342,G3343,G3344,G3345,G3346,G3347,G3348,G3349,G3350,G3351,G3352,G3353,G3354,G3355,G3356,G3357,G3358,G3359,G3360,
       G3361,G3362,G3363,G3364,G3365,G3366,G3367,G3368,G3369,G3370,G3371,G3372,G3373,G3374,G3375,G3376,G3377,G3378,G3379,G3380,
       G3381,G3382,G3383,G3384,G3385,G3386,G3387,G3388,G3389,G3390,G3391,G3392,G3393,G3394,G3395,G3396,G3397,G3398,G3399,G3400,
       G3401,G3402,G3403,G3404,G3405,G3406,G3407,G3408,G3409,G3410,G3411,G3412,G3413,G3414,G3415,G3416,G3417,G3418,G3419,G3420,
       G3421,G3422,G3423,G3424,G3425,G3426,G3427,G3428,G3429,G3430,G3431,G3432,G3433,G3434,G3435,G3436,G3437,G3438,G3439,G3440,
       G3441,G3442,G3443,G3444,G3445,G3446,G3447,G3448,G3449,G3450,G3451,G3452,G3453,G3454,G3455,G3456,G3457,G3458,G3459,G3460,
       G3461,G3462,G3463,G3464,G3465,G3466,G3467,G3468,G3469,G3470,G3471,G3472,G3473,G3474,G3475,G3476,G3477,G3478,G3479,G3480,
       G3481,G3482,G3483,G3484,G3485,G3486,G3487,G3488,G3489,G3490,G3491,G3492,G3493,G3494,G3495,G3496,G3497,G3498,G3499,G3500,
       G3501,G3502,G3503,G3504,G3505,G3506,G3507,G3508,G3509,G3510,G3511,G3512,G3513,G3514,G3515,G3516,G3517,G3518,G3519,G3520,
       G3521,G3522,G3523,G3524,G3525,G3526,G3527,G3528,G3529,G3530,G3531,G3532,G3533,G3534,G3535,G3536,G3537,G3538,G3539,G3540,
       G3541,G3542,G3543,G3544,G3545,G3546,G3547,G3548,G3549,G3550,G3551,G3552,G3553,G3554,G3555,G3556,G3557,G3558,G3559,G3560,
       G3561,G3562,G3563,G3564,G3565,G3566,G3567,G3568,G3569,G3570,G3571,G3572,G3573,G3574,G3575,G3576,G3577,G3578,G3579,G3580,
       G3581,G3582,G3583,G3584,G3585,G3586,G3587,G3588,G3589,G3590,G3591,G3592,G3593,G3594,G3595,G3596,G3597,G3598,G3599,G3600,
       G3601,G3602,G3603,G3604,G3605,G3606,G3607,G3608,G3609,G3610,G3611,G3612,G3613,G3614,G3615,G3616,G3617,G3618,G3619,G3620,
       G3621,G3622,G3623,G3624,G3625,G3626,G3627,G3628,G3629,G3630,G3631,G3632,G3633,G3634,G3635,G3636,G3637,G3638,G3639,G3640,
       G3641,G3642,G3643,G3644,G3645,G3646,G3647,G3648,G3649,G3650,G3651,G3652,G3653,G3654,G3655,G3656,G3657,G3658,G3659,G3660,
       G3661,G3662,G3663,G3664,G3665,G3666,G3667,G3668,G3669,G3670,G3671,G3672,G3673,G3674,G3675,G3676,G3677,G3678,G3679,G3680,
       G3681,G3682,G3683,G3684,G3685,G3686,G3687,G3688,G3689,G3690,G3691,G3692,G3693,G3694,G3695,G3696,G3697,G3698,G3699,G3700,
       G3701,G3702,G3703,G3704,G3705,G3706,G3707,G3708,G3709,G3710,G3711,G3712,G3713,G3714,G3715,G3716,G3717,G3718,G3719,G3720,
       G3721,G3722,G3723,G3724,G3725,G3726,G3727,G3728,G3729,G3730,G3731,G3732,G3733,G3734,G3735,G3736,G3737,G3738,G3739,G3740,
       G3741,G3742,G3743,G3744,G3745,G3746,G3747,G3748,G3749,G3750,G3751,G3752,G3753,G3754,G3755,G3756,G3757,G3758,G3759,G3760,
       G3761,G3762,G3763,G3764,G3765,G3766,G3767,G3768,G3769,G3770,G3771,G3772,G3773,G3774,G3775,G3776,G3777,G3778,G3779,G3780,
       G3781,G3782,G3783,G3784,G3785,G3786,G3787,G3788,G3789,G3790,G3791,G3792,G3793,G3794,G3795,G3796,G3797,G3798,G3799,G3800,
       G3801,G3802,G3803,G3804,G3805,G3806,G3807,G3808,G3809,G3810,G3811,G3812,G3813,G3814,G3815,G3816,G3817,G3818,G3819,G3820,
       G3821,G3822,G3823,G3824,G3825,G3826,G3827,G3828,G3829,G3830,G3831,G3832,G3833,G3834,G3835,G3836,G3837,G3838,G3839,G3840,
       G3841,G3842,G3843,G3844,G3845,G3846,G3847,G3848,G3849,G3850,G3851,G3852,G3853,G3854,G3855,G3856,G3857,G3858,G3859,G3860,
       G3861,G3862,G3863,G3864,G3865,G3866,G3867,G3868,G3869,G3870,G3871,G3872,G3873,G3874,G3875,G3876,G3877,G3878,G3879,G3880,
       G3881,G3882,G3883,G3884,G3885,G3886,G3887,G3888,G3889,G3890,G3891,G3892,G3893,G3894,G3895,G3896,G3897,G3898,G3899,G3900,
       G3901,G3902,G3903,G3904,G3905,G3906,G3907,G3908,G3909,G3910,G3911,G3912,G3913,G3914,G3915,G3916,G3917,G3918,G3919,G3920,
       G3921,G3922,G3923,G3924,G3925,G3926,G3927,G3928,G3929,G3930,G3931,G3932,G3933,G3934,G3935,G3936,G3937,G3938,G3939,G3940,
       G3941,G3942,G3943,G3944,G3945,G3946,G3947,G3948,G3949,G3950,G3951,G3952,G3953,G3954,G3955,G3956,G3957,G3958,G3959,G3960,
       G3961,G3962,G3963,G3964,G3965,G3966,G3967,G3968,G3969,G3970,G3971,G3972,G3973,G3974,G3975,G3976,G3977,G3978,G3979,G3980,
       G3981,G3982,G3983,G3984,G3985,G3986,G3987,G3988,G3989,G3990,G3991,G3992,G3993,G3994,G3995,G3996,G3997,G3998,G3999,G4000,
       G4001,G4002,G4003,G4004,G4005,G4006,G4007,G4008,G4009,G4010,G4011,G4012,G4013,G4014,G4015,G4016,G4017,G4018,G4019,G4020,
       G4021,G4022,G4023,G4024,G4025,G4026,G4027,G4028,G4029,G4030,G4031,G4032,G4033,G4034,G4035,G4036,G4037,G4038,G4039,G4040,
       G4041,G4042,G4043,G4044,G4045,G4046,G4047,G4048,G4049,G4050,G4051,G4052,G4053,G4054,G4055,G4056,G4057,G4058,G4059,G4060,
       G4061,G4062,G4063,G4064,G4065,G4066,G4067,G4068,G4069,G4070,G4071,G4072,G4073,G4074,G4075,G4076,G4077,G4078,G4079,G4080,
       G4081,G4082,G4083,G4084,G4085,G4086,G4087,G4088,G4089,G4090,G4091,G4092,G4093,G4094,G4095,G4096,G4097,G4098,G4099,G4100,
       G4101,G4102,G4103,G4104,G4105,G4106,G4107,G4108,G4109,G4110,G4111,G4112,G4113,G4114,G4115,G4116,G4117,G4118,G4119,G4120,
       G4121,G4122,G4123,G4124,G4125,G4126,G4127,G4128,G4129,G4130,G4131,G4132,G4133,G4134,G4135,G4136,G4137,G4138,G4139,G4140,
       G4141,G4142,G4143,G4144,G4145,G4146,G4147,G4148,G4149,G4150,G4151,G4152,G4153,G4154,G4155,G4156,G4157,G4158,G4159,G4160,
       G4161,G4162,G4163,G4164,G4165,G4166,G4167,G4168,G4169,G4170,G4171,G4172,G4173,G4174,G4175,G4176,G4177,G4178,G4179,G4180,
       G4181,G4182,G4183,G4184,G4185,G4186,G4187,G4188,G4189,G4190,G4191,G4192,G4193,G4194,G4195,G4196,G4197,G4198,G4199,G4200,
       G4201,G4202,G4203,G4204,G4205,G4206,G4207,G4208,G4209,G4210,G4211,G4212,G4213,G4214,G4215,G4216,G4217,G4218,G4219,G4220,
       G4221,G4222,G4223,G4224,G4225,G4226,G4227,G4228,G4229,G4230,G4231,G4232,G4233,G4234,G4235,G4236,G4237,G4238,G4239,G4240,
       G4241,G4242,G4243,G4244,G4245,G4246,G4247,G4248,G4249,G4250,G4251,G4252,G4253,G4254,G4255,G4256,G4257,G4258,G4259,G4260,
       G4261,G4262,G4263,G4264,G4265,G4266,G4267,G4268,G4269,G4270,G4271,G4272,G4273,G4274,G4275,G4276,G4277,G4278,G4279,G4280,
       G4281,G4282,G4283,G4284,G4285,G4286,G4287,G4288,G4289,G4290,G4291,G4292,G4293,G4294,G4295,G4296,G4297,G4298,G4299,G4300,
       G4301,G4302,G4303,G4304,G4305,G4306,G4307,G4308,G4309,G4310,G4311,G4312,G4313,G4314,G4315,G4316,G4317,G4318,G4319,G4320,
       G4321,G4322,G4323,G4324,G4325,G4326,G4327,G4328,G4329,G4330,G4331,G4332,G4333,G4334,G4335,G4336,G4337,G4338,G4339,G4340,
       G4341,G4342,G4343,G4344,G4345,G4346,G4347,G4348,G4349,G4350,G4351,G4352,G4353,G4354,G4355,G4356,G4357,G4358,G4359,G4360,
       G4361,G4362,G4363,G4364,G4365,G4366,G4367,G4368,G4369,G4370,G4371,G4372,G4373,G4374,G4375,G4376,G4377,G4378,G4379,G4380,
       G4381,G4382,G4383,G4384,G4385,G4386,G4387,G4388,G4389,G4390,G4391,G4392,G4393,G4394,G4395,G4396,G4397,G4398,G4399,G4400,
       G4401,G4402,G4403,G4404,G4405,G4406,G4407,G4408,G4409,G4410,G4411,G4412,G4413,G4414,G4415,G4416,G4417,G4418,G4419,G4420,
       G4421,G4422,G4423,G4424,G4425,G4426,G4427,G4428,G4429,G4430,G4431,G4432,G4433,G4434,G4435,G4436,G4437,G4438,G4439,G4440,
       G4441,G4442,G4443,G4444,G4445,G4446,G4447,G4448,G4449,G4450,G4451,G4452,G4453,G4454,G4455,G4456,G4457,G4458,G4459,G4460,
       G4461,G4462,G4463,G4464,G4465,G4466,G4467,G4468,G4469,G4470,G4471,G4472,G4473,G4474,G4475,G4476,G4477,G4478,G4479,G4480,
       G4481,G4482,G4483,G4484,G4485,G4486,G4487,G4488,G4489,G4490,G4491,G4492,G4493,G4494,G4495,G4496,G4497,G4498,G4499,G4500,
       G4501,G4502,G4503,G4504,G4505,G4506,G4507,G4508,G4509,G4510,G4511,G4512,G4513,G4514,G4515,G4516,G4517,G4518,G4519,G4520,
       G4521,G4522,G4523,G4524,G4525,G4526,G4527,G4528,G4529,G4530,G4531,G4532,G4533,G4534,G4535,G4536,G4537,G4538,G4539,G4540,
       G4541,G4542,G4543,G4544,G4545,G4546,G4547,G4548,G4549,G4550,G4551,G4552,G4553,G4554,G4555,G4556,G4557,G4558,G4559,G4560,
       G4561,G4562,G4563,G4564,G4565,G4566,G4567,G4568,G4569,G4570,G4571,G4572,G4573,G4574,G4575,G4576,G4577,G4578,G4579,G4580,
       G4581,G4582,G4583,G4584,G4585,G4586,G4587,G4588,G4589,G4590,G4591,G4592,G4593,G4594,G4595,G4596,G4597,G4598,G4599,G4600,
       G4601,G4602,G4603,G4604,G4605,G4606,G4607,G4608,G4609,G4610,G4611,G4612,G4613,G4614,G4615,G4616,G4617,G4618,G4619,G4620,
       G4621,G4622,G4623,G4624,G4625,G4626,G4627,G4628,G4629,G4630,G4631,G4632,G4633,G4634,G4635,G4636,G4637,G4638,G4639,G4640,
       G4641,G4642,G4643,G4644,G4645,G4646,G4647,G4648,G4649,G4650,G4651,G4652,G4653,G4654,G4655,G4656,G4657,G4658,G4659,G4660,
       G4661,G4662,G4663,G4664,G4665,G4666,G4667,G4668,G4669,G4670,G4671,G4672,G4673,G4674,G4675,G4676,G4677,G4678,G4679,G4680,
       G4681,G4682,G4683,G4684,G4685,G4686,G4687,G4688,G4689,G4690,G4691,G4692,G4693,G4694,G4695,G4696,G4697,G4698,G4699,G4700,
       G4701,G4702,G4703,G4704,G4705,G4706,G4707,G4708,G4709,G4710,G4711,G4712,G4713,G4714,G4715,G4716,G4717,G4718,G4719,G4720,
       G4721,G4722,G4723,G4724,G4725,G4726,G4727,G4728,G4729,G4730,G4731,G4732,G4733,G4734,G4735,G4736,G4737,G4738,G4739,G4740,
       G4741,G4742,G4743,G4744,G4745,G4746,G4747,G4748,G4749,G4750,G4751,G4752,G4753,G4754,G4755,G4756,G4757,G4758,G4759,G4760,
       G4761,G4762,G4763,G4764,G4765,G4766,G4767,G4768,G4769,G4770,G4771,G4772,G4773,G4774,G4775,G4776,G4777,G4778,G4779,G4780,
       G4781,G4782,G4783,G4784,G4785,G4786,G4787,G4788,G4789,G4790,G4791,G4792,G4793,G4794,G4795,G4796,G4797,G4798,G4799,G4800,
       G4801,G4802,G4803,G4804,G4805,G4806,G4807,G4808,G4809,G4810,G4811,G4812,G4813,G4814,G4815,G4816,G4817,G4818,G4819,G4820,
       G4821,G4822,G4823,G4824,G4825,G4826,G4827,G4828,G4829,G4830,G4831,G4832,G4833,G4834,G4835,G4836,G4837,G4838,G4839,G4840,
       G4841,G4842,G4843,G4844,G4845,G4846,G4847,G4848,G4849,G4850,G4851,G4852,G4853,G4854,G4855,G4856,G4857,G4858,G4859,G4860,
       G4861,G4862,G4863,G4864,G4865,G4866,G4867,G4868,G4869,G4870,G4871,G4872,G4873,G4874,G4875,G4876,G4877,G4878,G4879,G4880,
       G4881,G4882,G4883,G4884,G4885,G4886,G4887,G4888,G4889,G4890,G4891,G4892,G4893,G4894,G4895,G4896,G4897,G4898,G4899,G4900,
       G4901,G4902,G4903,G4904,G4905,G4906,G4907,G4908,G4909,G4910,G4911,G4912,G4913,G4914,G4915,G4916,G4917,G4918,G4919,G4920,
       G4921,G4922,G4923,G4924,G4925,G4926,G4927,G4928,G4929,G4930,G4931,G4932,G4933,G4934,G4935,G4936,G4937,G4938,G4939,G4940,
       G4941,G4942,G4943,G4944,G4945,G4946,G4947,G4948,G4949,G4950,G4951,G4952,G4953,G4954,G4955,G4956,G4957,G4958,G4959,G4960,
       G4961,G4962,G4963,G4964,G4965,G4966,G4967,G4968,G4969,G4970,G4971,G4972,G4973,G4974,G4975,G4976,G4977,G4978,G4979,G4980,
       G4981,G4982,G4983,G4984,G4985,G4986,G4987,G4988,G4989,G4990,G4991,G4992,G4993,G4994,G4995,G4996,G4997,G4998,G4999,G5000,
       G5001,G5002,G5003,G5004,G5005,G5006,G5007,G5008,G5009,G5010,G5011,G5012,G5013,G5014,G5015,G5016,G5017,G5018,G5019,G5020,
       G5021,G5022,G5023,G5024,G5025,G5026,G5027,G5028,G5029,G5030,G5031,G5032,G5033,G5034,G5035,G5036,G5037,G5038,G5039,G5040,
       G5041,G5042,G5043,G5044,G5045,G5046,G5047,G5048,G5049,G5050,G5051,G5052,G5053,G5054,G5055,G5056,G5057,G5058,G5059,G5060,
       G5061,G5062,G5063,G5064,G5065,G5066,G5067,G5068,G5069,G5070,G5071,G5072,G5073,G5074,G5075,G5076,G5077,G5078,G5079,G5080,
       G5081,G5082,G5083,G5084,G5085,G5086,G5087,G5088,G5089,G5090,G5091,G5092,G5093,G5094,G5095,G5096,G5097,G5098,G5099,G5100,
       G5101,G5102,G5103,G5104,G5105,G5106,G5107,G5108,G5109,G5110,G5111,G5112,G5113,G5114,G5115,G5116,G5117,G5118,G5119,G5120,
       G5121,G5122,G5123,G5124,G5125,G5126,G5127,G5128,G5129,G5130,G5131,G5132,G5133,G5134,G5135,G5136,G5137,G5138,G5139,G5140,
       G5141,G5142,G5143,G5144,G5145,G5146,G5147,G5148,G5149,G5150,G5151,G5152,G5153,G5154,G5155,G5156,G5157,G5158,G5159,G5160,
       G5161,G5162,G5163,G5164,G5165,G5166,G5167,G5168,G5169,G5170,G5171,G5172,G5173,G5174,G5175,G5176,G5177,G5178,G5179,G5180,
       G5181,G5182,G5183,G5184,G5185,G5186,G5187,G5188,G5189,G5190,G5191,G5192,G5193,G5194,G5195,G5196,G5197,G5198,G5199,G5200,
       G5201,G5202,G5203,G5204,G5205,G5206,G5207,G5208,G5209,G5210,G5211,G5212,G5213,G5214,G5215,G5216,G5217,G5218,G5219,G5220,
       G5221,G5222,G5223,G5224,G5225,G5226,G5227,G5228,G5229,G5230,G5231,G5232,G5233,G5234,G5235,G5236,G5237,G5238,G5239,G5240,
       G5241,G5242,G5243,G5244,G5245,G5246,G5247,G5248,G5249,G5250,G5251,G5252,G5253,G5254,G5255,G5256,G5257,G5258,G5259,G5260,
       G5261,G5262,G5263,G5264,G5265,G5266,G5267,G5268,G5269,G5270,G5271,G5272,G5273,G5274,G5275,G5276,G5277,G5278,G5279,G5280,
       G5281,G5282,G5283,G5284,G5285,G5286,G5287,G5288,G5289,G5290,G5291,G5292,G5293,G5294,G5295,G5296,G5297,G5298,G5299,G5300,
       G5301,G5302,G5303,G5304,G5305,G5306,G5307,G5308,G5309,G5310,G5311,G5312,G5313,G5314,G5315,G5316,G5317,G5318,G5319,G5320,
       G5321,G5322,G5323,G5324,G5325,G5326,G5327,G5328,G5329,G5330,G5331,G5332,G5333,G5334,G5335,G5336,G5337,G5338,G5339,G5340,
       G5341,G5342,G5343,G5344,G5345,G5346,G5347,G5348,G5349,G5350,G5351,G5352,G5353,G5354,G5355,G5356,G5357,G5358,G5359,G5360,
       G5361,G5362,G5363,G5364,G5365,G5366,G5367,G5368,G5369,G5370,G5371,G5372,G5373,G5374,G5375,G5376,G5377,G5378,G5379,G5380,
       G5381,G5382,G5383,G5384,G5385,G5386,G5387,G5388,G5389,G5390,G5391,G5392,G5393,G5394,G5395,G5396,G5397,G5398,G5399,G5400,
       G5401,G5402,G5403,G5404,G5405,G5406,G5407,G5408,G5409,G5410,G5411,G5412,G5413,G5414,G5415,G5416,G5417,G5418,G5419,G5420,
       G5421,G5422,G5423,G5424,G5425,G5426,G5427,G5428,G5429,G5430,G5431,G5432,G5433,G5434,G5435,G5436,G5437,G5438,G5439,G5440,
       G5441,G5442,G5443,G5444,G5445,G5446,G5447,G5448,G5449,G5450,G5451,G5452,G5453,G5454,G5455,G5456,G5457,G5458,G5459,G5460,
       G5461,G5462,G5463,G5464,G5465,G5466,G5467,G5468,G5469,G5470,G5471,G5472,G5473,G5474,G5475,G5476,G5477,G5478,G5479,G5480,
       G5481,G5482,G5483,G5484,G5485,G5486,G5487,G5488,G5489,G5490,G5491,G5492,G5493,G5494,G5495,G5496,G5497,G5498,G5499,G5500,
       G5501,G5502,G5503,G5504,G5505,G5506,G5507,G5508,G5509,G5510,G5511,G5512,G5513,G5514,G5515,G5516,G5517,G5518,G5519,G5520,
       G5521,G5522,G5523,G5524,G5525,G5526,G5527,G5528,G5529,G5530,G5531,G5532,G5533,G5534,G5535,G5536,G5537,G5538,G5539,G5540,
       G5541,G5542,G5543,G5544,G5545,G5546,G5547,G5548,G5549,G5550,G5551,G5552,G5553,G5554,G5555,G5556,G5557,G5558,G5559,G5560,
       G5561,G5562,G5563,G5564,G5565,G5566,G5567,G5568,G5569,G5570,G5571,G5572,G5573,G5574,G5575,G5576,G5577,G5578,G5579,G5580,
       G5581,G5582,G5583,G5584,G5585,G5586,G5587,G5588,G5589,G5590,G5591,G5592,G5593,G5594,G5595,G5596,G5597,G5598,G5599,G5600,
       G5601,G5602,G5603,G5604,G5605,G5606,G5607,G5608,G5609,G5610,G5611,G5612,G5613,G5614,G5615,G5616,G5617,G5618,G5619,G5620,
       G5621,G5622,G5623,G5624,G5625,G5626,G5627,G5628,G5629,G5630,G5631,G5632,G5633,G5634,G5635,G5636,G5637,G5638,G5639,G5640,
       G5641,G5642,G5643,G5644,G5645,G5646,G5647,G5648,G5649,G5650,G5651,G5652,G5653,G5654,G5655,G5656,G5657,G5658,G5659,G5660,
       G5661,G5662,G5663,G5664,G5665,G5666,G5667,G5668,G5669,G5670,G5671,G5672,G5673,G5674,G5675,G5676,G5677,G5678,G5679,G5680,
       G5681,G5682,G5683,G5684,G5685,G5686,G5687,G5688,G5689,G5690,G5691,G5692,G5693,G5694,G5695,G5696,G5697,G5698,G5699,G5700,
       G5701,G5702,G5703,G5704,G5705,G5706,G5707,G5708,G5709,G5710,G5711,G5712,G5713,G5714,G5715,G5716,G5717,G5718,G5719,G5720,
       G5721,G5722,G5723,G5724,G5725,G5726,G5727,G5728,G5729,G5730,G5731,G5732,G5733,G5734,G5735,G5736,G5737,G5738,G5739,G5740,
       G5741,G5742,G5743,G5744,G5745,G5746,G5747,G5748,G5749,G5750,G5751,G5752,G5753,G5754,G5755,G5756,G5757,G5758,G5759,G5760,
       G5761,G5762,G5763,G5764,G5765,G5766,G5767,G5768,G5769,G5770,G5771,G5772,G5773,G5774,G5775,G5776,G5777,G5778,G5779,G5780,
       G5781,G5782,G5783,G5784,G5785,G5786,G5787,G5788,G5789,G5790,G5791,G5792,G5793,G5794,G5795,G5796,G5797,G5798,G5799,G5800,
       G5801,G5802,G5803,G5804,G5805,G5806,G5807,G5808,G5809,G5810,G5811,G5812,G5813,G5814,G5815,G5816,G5817,G5818,G5819,G5820,
       G5821,G5822,G5823,G5824,G5825,G5826,G5827,G5828,G5829,G5830,G5831,G5832,G5833,G5834,G5835,G5836,G5837,G5838,G5839,G5840,
       G5841,G5842,G5843,G5844,G5845,G5846,G5847,G5848,G5849,G5850,G5851,G5852,G5853,G5854,G5855,G5856,G5857,G5858,G5859,G5860,
       G5861,G5862,G5863,G5864,G5865,G5866,G5867,G5868,G5869,G5870,G5871,G5872,G5873,G5874,G5875,G5876,G5877,G5878,G5879,G5880,
       G5881,G5882,G5883,G5884,G5885,G5886,G5887,G5888,G5889,G5890,G5891,G5892,G5893,G5894,G5895,G5896,G5897,G5898,G5899,G5900,
       G5901,G5902,G5903,G5904,G5905,G5906,G5907,G5908,G5909,G5910,G5911,G5912,G5913,G5914,G5915,G5916,G5917,G5918,G5919,G5920,
       G5921,G5922,G5923,G5924,G5925,G5926,G5927,G5928,G5929,G5930,G5931,G5932,G5933,G5934,G5935,G5936,G5937,G5938,G5939,G5940,
       G5941,G5942,G5943,G5944,G5945,G5946,G5947,G5948,G5949,G5950,G5951,G5952,G5953,G5954,G5955,G5956,G5957,G5958,G5959,G5960,
       G5961,G5962,G5963,G5964,G5965,G5966,G5967,G5968,G5969,G5970,G5971,G5972,G5973,G5974,G5975,G5976,G5977,G5978,G5979,G5980,
       G5981,G5982,G5983,G5984,G5985,G5986,G5987,G5988,G5989,G5990,G5991,G5992,G5993,G5994,G5995,G5996,G5997,G5998,G5999,G6000,
       G6001,G6002,G6003,G6004,G6005,G6006,G6007,G6008,G6009,G6010,G6011,G6012,G6013,G6014,G6015,G6016,G6017,G6018,G6019,G6020,
       G6021,G6022,G6023,G6024,G6025,G6026,G6027,G6028,G6029,G6030,G6031,G6032,G6033,G6034,G6035,G6036,G6037,G6038,G6039,G6040,
       G6041,G6042,G6043,G6044,G6045,G6046,G6047,G6048,G6049,G6050,G6051,G6052,G6053,G6054,G6055,G6056,G6057,G6058,G6059,G6060,
       G6061,G6062,G6063,G6064,G6065,G6066,G6067,G6068,G6069,G6070,G6071,G6072,G6073,G6074,G6075,G6076,G6077,G6078,G6079,G6080,
       G6081,G6082,G6083,G6084,G6085,G6086,G6087,G6088,G6089,G6090,G6091,G6092,G6093,G6094,G6095,G6096,G6097,G6098,G6099,G6100,
       G6101,G6102,G6103,G6104,G6105,G6106,G6107,G6108,G6109,G6110,G6111,G6112,G6113,G6114,G6115,G6116,G6117,G6118,G6119,G6120,
       G6121,G6122,G6123,G6124,G6125,G6126,G6127,G6128,G6129,G6130,G6131,G6132,G6133,G6134,G6135,G6136,G6137,G6138,G6139,G6140,
       G6141,G6142,G6143,G6144,G6145,G6146,G6147,G6148,G6149,G6150,G6151,G6152,G6153,G6154,G6155,G6156,G6157,G6158,G6159,G6160,
       G6161,G6162,G6163,G6164,G6165,G6166,G6167,G6168,G6169,G6170,G6171,G6172,G6173,G6174,G6175,G6176,G6177,G6178,G6179,G6180,
       G6181,G6182,G6183,G6184,G6185,G6186,G6187,G6188,G6189,G6190,G6191,G6192,G6193,G6194,G6195,G6196,G6197,G6198,G6199,G6200,
       G6201,G6202,G6203,G6204,G6205,G6206,G6207,G6208,G6209,G6210,G6211,G6212,G6213,G6214,G6215,G6216,G6217,G6218,G6219,G6220,
       G6221,G6222,G6223,G6224,G6225,G6226,G6227,G6228,G6229,G6230,G6231,G6232,G6233,G6234,G6235,G6236,G6237,G6238,G6239,G6240,
       G6241,G6242,G6243,G6244,G6245,G6246,G6247,G6248,G6249,G6250,G6251,G6252,G6253,G6254,G6255,G6256,G6257,G6258,G6259,G6260,
       G6261,G6262,G6263,G6264,G6265,G6266,G6267,G6268,G6269,G6270,G6271,G6272,G6273,G6274,G6275,G6276,G6277,G6278,G6279,G6280,
       G6281,G6282,G6283,G6284,G6285,G6286,G6287,G6288,G6289,G6290,G6291,G6292,G6293,G6294,G6295,G6296,G6297,G6298,G6299,G6300,
       G6301,G6302,G6303,G6304,G6305,G6306,G6307,G6308,G6309,G6310,G6311,G6312,G6313,G6314,G6315,G6316,G6317,G6318,G6319,G6320,
       G6321,G6322,G6323,G6324,G6325,G6326,G6327,G6328,G6329,G6330,G6331,G6332,G6333,G6334,G6335,G6336,G6337,G6338,G6339,G6340,
       G6341,G6342,G6343,G6344,G6345,G6346,G6347,G6348,G6349,G6350,G6351,G6352,G6353,G6354,G6355,G6356,G6357,G6358,G6359,G6360,
       G6361,G6362,G6363,G6364,G6365,G6366,G6367,G6368,G6369,G6370,G6371,G6372,G6373,G6374,G6375,G6376,G6377,G6378,G6379,G6380,
       G6381,G6382,G6383,G6384,G6385,G6386,G6387,G6388,G6389,G6390,G6391,G6392,G6393,G6394,G6395,G6396,G6397,G6398,G6399,G6400,
       G6401,G6402,G6403,G6404,G6405,G6406,G6407,G6408,G6409,G6410,G6411,G6412,G6413,G6414,G6415,G6416,G6417,G6418,G6419,G6420,
       G6421,G6422,G6423,G6424,G6425,G6426,G6427,G6428,G6429,G6430,G6431,G6432,G6433,G6434,G6435,G6436,G6437,G6438,G6439,G6440,
       G6441,G6442,G6443,G6444,G6445,G6446,G6447,G6448,G6449,G6450,G6451,G6452,G6453,G6454,G6455,G6456,G6457,G6458,G6459,G6460,
       G6461,G6462,G6463,G6464,G6465,G6466,G6467,G6468,G6469,G6470,G6471,G6472,G6473,G6474,G6475,G6476,G6477,G6478,G6479,G6480,
       G6481,G6482,G6483,G6484,G6485,G6486,G6487,G6488,G6489,G6490,G6491,G6492,G6493,G6494,G6495,G6496,G6497,G6498,G6499,G6500,
       G6501,G6502,G6503,G6504,G6505,G6506,G6507,G6508,G6509,G6510,G6511,G6512,G6513,G6514,G6515,G6516,G6517,G6518,G6519,G6520,
       G6521,G6522,G6523,G6524,G6525,G6526,G6527,G6528,G6529,G6530,G6531,G6532,G6533,G6534,G6535,G6536,G6537,G6538,G6539,G6540,
       G6541,G6542,G6543,G6544,G6545,G6546,G6547,G6548,G6549,G6550,G6551,G6552,G6553,G6554,G6555,G6556,G6557,G6558,G6559,G6560,
       G6561,G6562,G6563,G6564,G6565,G6566,G6567,G6568,G6569,G6570,G6571,G6572,G6573,G6574,G6575,G6576,G6577,G6578,G6579,G6580,
       G6581,G6582,G6583,G6584,G6585,G6586,G6587,G6588,G6589,G6590,G6591,G6592,G6593,G6594,G6595,G6596,G6597,G6598,G6599,G6600,
       G6601,G6602,G6603,G6604,G6605,G6606,G6607,G6608,G6609,G6610,G6611,G6612,G6613,G6614,G6615,G6616,G6617,G6618,G6619,G6620,
       G6621,G6622,G6623,G6624,G6625,G6626,G6627,G6628,G6629,G6630,G6631,G6632,G6633,G6634,G6635,G6636,G6637,G6638,G6639,G6640,
       G6641,G6642,G6643,G6644,G6645,G6646,G6647,G6648,G6649,G6650,G6651,G6652,G6653,G6654,G6655,G6656,G6657,G6658,G6659,G6660,
       G6661,G6662,G6663,G6664,G6665,G6666,G6667,G6668,G6669,G6670,G6671,G6672,G6673,G6674,G6675,G6676,G6677,G6678,G6679,G6680,
       G6681,G6682,G6683,G6684,G6685,G6686,G6687,G6688,G6689,G6690,G6691,G6692,G6693,G6694,G6695,G6696,G6697,G6698,G6699,G6700,
       G6701,G6702,G6703,G6704,G6705,G6706,G6707,G6708,G6709,G6710,G6711,G6712,G6713,G6714,G6715,G6716,G6717,G6718,G6719,G6720,
       G6721,G6722,G6723,G6724,G6725,G6726,G6727,G6728,G6729,G6730,G6731,G6732,G6733,G6734,G6735,G6736,G6737,G6738,G6739,G6740,
       G6741,G6742,G6743,G6744,G6745,G6746,G6747,G6748,G6749,G6750,G6751,G6752,G6753,G6754,G6755,G6756,G6757,G6758,G6759,G6760,
       G6761,G6762,G6763,G6764,G6765,G6766,G6767,G6768,G6769,G6770,G6771,G6772,G6773,G6774,G6775,G6776,G6777,G6778,G6779,G6780,
       G6781,G6782,G6783,G6784,G6785,G6786,G6787,G6788,G6789,G6790,G6791,G6792,G6793,G6794,G6795,G6796,G6797,G6798,G6799,G6800,
       G6801,G6802,G6803,G6804,G6805,G6806,G6807,G6808,G6809,G6810,G6811,G6812,G6813,G6814,G6815,G6816,G6817,G6818,G6819,G6820,
       G6821,G6822,G6823,G6824,G6825,G6826,G6827,G6828,G6829,G6830,G6831,G6832,G6833,G6834,G6835,G6836,G6837,G6838,G6839,G6840,
       G6841,G6842,G6843,G6844,G6845,G6846,G6847,G6848,G6849,G6850,G6851,G6852,G6853,G6854,G6855,G6856,G6857,G6858,G6859,G6860,
       G6861,G6862,G6863,G6864,G6865,G6866,G6867,G6868,G6869,G6870,G6871,G6872,G6873,G6874,G6875,G6876,G6877,G6878,G6879,G6880,
       G6881,G6882,G6883,G6884,G6885,G6886,G6887,G6888,G6889,G6890,G6891,G6892,G6893,G6894,G6895,G6896,G6897,G6898,G6899,G6900,
       G6901,G6902,G6903,G6904,G6905,G6906,G6907,G6908,G6909,G6910,G6911,G6912,G6913,G6914,G6915,G6916,G6917,G6918,G6919,G6920,
       G6921,G6922,G6923,G6924,G6925,G6926,G6927,G6928,G6929,G6930,G6931,G6932,G6933,G6934,G6935,G6936,G6937,G6938,G6939,G6940,
       G6941,G6942,G6943,G6944,G6945,G6946,G6947,G6948,G6949,G6950,G6951,G6952,G6953,G6954,G6955,G6956,G6957,G6958,G6959,G6960,
       G6961,G6962,G6963,G6964,G6965,G6966,G6967,G6968,G6969,G6970,G6971,G6972,G6973,G6974,G6975,G6976,G6977,G6978,G6979,G6980,
       G6981,G6982,G6983,G6984,G6985,G6986,G6987,G6988,G6989,G6990,G6991,G6992,G6993,G6994,G6995,G6996,G6997,G6998,G6999,G7000,
       G7001,G7002,G7003,G7004,G7005,G7006,G7007,G7008,G7009,G7010,G7011,G7012,G7013,G7014,G7015,G7016,G7017,G7018,G7019,G7020,
       G7021,G7022,G7023,G7024,G7025,G7026,G7027,G7028,G7029,G7030,G7031,G7032,G7033,G7034,G7035,G7036,G7037,G7038,G7039,G7040,
       G7041,G7042,G7043,G7044,G7045,G7046,G7047,G7048,G7049,G7050,G7051,G7052,G7053,G7054,G7055,G7056,G7057,G7058,G7059,G7060,
       G7061,G7062,G7063,G7064,G7065,G7066,G7067,G7068,G7069,G7070,G7071,G7072,G7073,G7074,G7075,G7076,G7077,G7078,G7079,G7080,
       G7081,G7082,G7083,G7084,G7085,G7086,G7087,G7088,G7089,G7090,G7091,G7092,G7093,G7094,G7095,G7096,G7097,G7098,G7099,G7100,
       G7101,G7102,G7103,G7104,G7105,G7106,G7107,G7108,G7109,G7110,G7111,G7112,G7113,G7114,G7115,G7116,G7117,G7118,G7119,G7120,
       G7121,G7122,G7123,G7124,G7125,G7126,G7127,G7128,G7129,G7130,G7131,G7132,G7133,G7134,G7135,G7136,G7137,G7138,G7139,G7140,
       G7141,G7142,G7143,G7144,G7145,G7146,G7147,G7148,G7149,G7150,G7151,G7152,G7153,G7154,G7155,G7156,G7157,G7158,G7159,G7160,
       G7161,G7162,G7163,G7164,G7165,G7166,G7167,G7168,G7169,G7170,G7171,G7172,G7173,G7174,G7175,G7176,G7177,G7178,G7179,G7180,
       G7181,G7182,G7183,G7184,G7185,G7186,G7187,G7188,G7189,G7190,G7191,G7192,G7193,G7194,G7195,G7196,G7197,G7198,G7199,G7200,
       G7201,G7202,G7203,G7204,G7205,G7206,G7207,G7208,G7209,G7210,G7211,G7212,G7213,G7214,G7215,G7216,G7217,G7218,G7219,G7220,
       G7221,G7222,G7223,G7224,G7225,G7226,G7227,G7228,G7229,G7230,G7231,G7232,G7233,G7234,G7235,G7236,G7237,G7238,G7239,G7240,
       G7241,G7242,G7243,G7244,G7245,G7246,G7247,G7248,G7249,G7250,G7251,G7252,G7253,G7254,G7255,G7256,G7257,G7258,G7259,G7260,
       G7261,G7262,G7263,G7264,G7265,G7266,G7267,G7268,G7269,G7270,G7271,G7272,G7273,G7274,G7275,G7276,G7277,G7278,G7279,G7280,
       G7281,G7282,G7283,G7284,G7285,G7286,G7287,G7288,G7289,G7290,G7291,G7292,G7293,G7294,G7295,G7296,G7297,G7298,G7299,G7300,
       G7301,G7302,G7303,G7304,G7305,G7306,G7307,G7308,G7309,G7310,G7311,G7312,G7313,G7314,G7315,G7316,G7317,G7318,G7319,G7320,
       G7321,G7322,G7323,G7324,G7325,G7326,G7327,G7328,G7329,G7330,G7331,G7332,G7333,G7334,G7335,G7336,G7337,G7338,G7339,G7340,
       G7341,G7342,G7343,G7344,G7345,G7346,G7347,G7348,G7349,G7350,G7351,G7352,G7353,G7354,G7355,G7356,G7357,G7358,G7359,G7360,
       G7361,G7362,G7363,G7364,G7365,G7366,G7367,G7368,G7369,G7370,G7371,G7372,G7373,G7374,G7375,G7376,G7377,G7378,G7379,G7380,
       G7381,G7382,G7383,G7384,G7385,G7386,G7387,G7388,G7389,G7390,G7391,G7392,G7393,G7394,G7395,G7396,G7397,G7398,G7399,G7400,
       G7401,G7402,G7403,G7404,G7405,G7406,G7407,G7408,G7409,G7410,G7411,G7412,G7413,G7414,G7415,G7416,G7417,G7418,G7419,G7420,
       G7421,G7422,G7423,G7424,G7425,G7426,G7427,G7428,G7429,G7430,G7431,G7432,G7433,G7434,G7435,G7436,G7437,G7438,G7439,G7440,
       G7441,G7442,G7443,G7444,G7445,G7446,G7447,G7448,G7449,G7450,G7451,G7452,G7453,G7454,G7455,G7456,G7457,G7458,G7459,G7460,
       G7461,G7462,G7463,G7464,G7465,G7466,G7467,G7468,G7469,G7470,G7471,G7472,G7473,G7474,G7475,G7476,G7477,G7478,G7479,G7480,
       G7481,G7482,G7483,G7484,G7485,G7486,G7487,G7488,G7489,G7490,G7491,G7492,G7493,G7494,G7495,G7496,G7497,G7498,G7499,G7500,
       G7501,G7502,G7503,G7504,G7505,G7506,G7507,G7508,G7509,G7510,G7511,G7512,G7513,G7514,G7515,G7516,G7517,G7518,G7519,G7520,
       G7521,G7522,G7523,G7524,G7525,G7526,G7527,G7528,G7529,G7530,G7531,G7532,G7533,G7534,G7535,G7536,G7537,G7538,G7539,G7540,
       G7541,G7542,G7543,G7544,G7545,G7546,G7547,G7548,G7549,G7550,G7551,G7552,G7553,G7554,G7555,G7556,G7557,G7558,G7559,G7560,
       G7561,G7562,G7563,G7564,G7565,G7566,G7567,G7568,G7569,G7570,G7571,G7572,G7573,G7574,G7575,G7576,G7577,G7578,G7579,G7580,
       G7581,G7582,G7583,G7584,G7585,G7586,G7587,G7588,G7589,G7590,G7591,G7592,G7593,G7594,G7595,G7596,G7597,G7598,G7599,G7600,
       G7601,G7602,G7603,G7604,G7605,G7606,G7607,G7608,G7609,G7610,G7611,G7612,G7613,G7614,G7615,G7616,G7617,G7618,G7619,G7620,
       G7621,G7622,G7623,G7624,G7625,G7626,G7627,G7628,G7629,G7630,G7631,G7632,G7633,G7634,G7635,G7636,G7637,G7638,G7639,G7640,
       G7641,G7642,G7643,G7644,G7645,G7646,G7647,G7648,G7649,G7650,G7651,G7652,G7653,G7654,G7655,G7656,G7657,G7658,G7659,G7660,
       G7661,G7662,G7663,G7664,G7665,G7666,G7667,G7668,G7669,G7670,G7671,G7672,G7673,G7674,G7675,G7676,G7677,G7678,G7679,G7680,
       G7681,G7682,G7683,G7684,G7685,G7686,G7687,G7688,G7689,G7690,G7691,G7692,G7693,G7694,G7695,G7696,G7697,G7698,G7699,G7700,
       G7701,G7702,G7703,G7704,G7705,G7706,G7707,G7708,G7709,G7710,G7711,G7712,G7713,G7714,G7715,G7716,G7717,G7718,G7719,G7720,
       G7721,G7722,G7723,G7724,G7725,G7726,G7727,G7728,G7729,G7730,G7731,G7732,G7733,G7734,G7735,G7736,G7737,G7738,G7739,G7740,
       G7741,G7742,G7743,G7744,G7745,G7746,G7747,G7748,G7749,G7750,G7751,G7752,G7753,G7754,G7755,G7756,G7757,G7758,G7759,G7760,
       G7761,G7762,G7763,G7764,G7765,G7766,G7767,G7768,G7769,G7770,G7771,G7772,G7773,G7774,G7775,G7776,G7777,G7778,G7779,G7780,
       G7781,G7782,G7783,G7784,G7785,G7786,G7787,G7788,G7789,G7790,G7791,G7792,G7793,G7794,G7795,G7796,G7797,G7798,G7799,G7800,
       G7801,G7802,G7803,G7804,G7805,G7806,G7807,G7808,G7809,G7810,G7811,G7812,G7813,G7814,G7815,G7816,G7817,G7818,G7819,G7820,
       G7821,G7822,G7823,G7824,G7825,G7826,G7827,G7828,G7829,G7830,G7831,G7832,G7833,G7834,G7835,G7836,G7837,G7838,G7839,G7840,
       G7841,G7842,G7843,G7844,G7845,G7846,G7847,G7848,G7849,G7850,G7851,G7852,G7853,G7854,G7855,G7856,G7857,G7858,G7859,G7860,
       G7861,G7862,G7863,G7864,G7865,G7866,G7867,G7868,G7869,G7870,G7871,G7872,G7873,G7874,G7875,G7876,G7877,G7878,G7879,G7880,
       G7881,G7882,G7883,G7884,G7885,G7886,G7887,G7888,G7889,G7890,G7891,G7892,G7893,G7894,G7895,G7896,G7897,G7898,G7899,G7900,
       G7901,G7902,G7903,G7904,G7905,G7906,G7907,G7908,G7909,G7910,G7911,G7912,G7913,G7914,G7915,G7916,G7917,G7918,G7919,G7920,
       G7921,G7922,G7923,G7924,G7925,G7926,G7927,G7928,G7929,G7930,G7931,G7932,G7933,G7934,G7935,G7936,G7937,G7938,G7939,G7940,
       G7941,G7942,G7943,G7944,G7945,G7946,G7947,G7948,G7949,G7950,G7951,G7952,G7953,G7954,G7955,G7956,G7957,G7958,G7959,G7960,
       G7961,G7962,G7963,G7964,G7965,G7966,G7967,G7968,G7969,G7970,G7971,G7972,G7973,G7974,G7975,G7976,G7977,G7978,G7979,G7980,
       G7981,G7982,G7983,G7984,G7985,G7986,G7987,G7988,G7989,G7990,G7991,G7992,G7993,G7994,G7995,G7996,G7997,G7998,G7999,G8000,
       G8001,G8002,G8003,G8004,G8005,G8006,G8007,G8008,G8009,G8010,G8011,G8012,G8013,G8014,G8015,G8016,G8017,G8018,G8019,G8020,
       G8021,G8022,G8023,G8024,G8025,G8026,G8027,G8028,G8029,G8030,G8031,G8032,G8033,G8034,G8035,G8036,G8037,G8038,G8039,G8040,
       G8041,G8042,G8043,G8044,G8045,G8046,G8047,G8048,G8049,G8050,G8051,G8052,G8053,G8054,G8055,G8056,G8057,G8058,G8059,G8060,
       G8061,G8062,G8063,G8064,G8065,G8066,G8067,G8068,G8069,G8070,G8071,G8072,G8073,G8074,G8075,G8076,G8077,G8078,G8079,G8080,
       G8081,G8082,G8083,G8084,G8085,G8086,G8087,G8088,G8089,G8090,G8091,G8092,G8093,G8094,G8095,G8096,G8097,G8098,G8099,G8100,
       G8101,G8102,G8103,G8104,G8105,G8106,G8107,G8108,G8109,G8110,G8111,G8112,G8113,G8114,G8115,G8116,G8117,G8118,G8119,G8120,
       G8121,G8122,G8123,G8124,G8125,G8126,G8127,G8128,G8129,G8130,G8131,G8132,G8133,G8134,G8135,G8136,G8137,G8138,G8139,G8140,
       G8141,G8142,G8143,G8144,G8145,G8146,G8147,G8148,G8149,G8150,G8151,G8152,G8153,G8154,G8155,G8156,G8157,G8158,G8159,G8160,
       G8161,G8162,G8163,G8164,G8165,G8166,G8167,G8168,G8169,G8170,G8171,G8172,G8173,G8174,G8175,G8176,G8177,G8178,G8179,G8180,
       G8181,G8182,G8183,G8184,G8185,G8186,G8187,G8188,G8189,G8190,G8191,G8192,G8193,G8194,G8195,G8196,G8197,G8198,G8199,G8200,
       G8201,G8202,G8203,G8204,G8205,G8206,G8207,G8208,G8209,G8210,G8211,G8212,G8213,G8214,G8215,G8216,G8217,G8218,G8219,G8220,
       G8221,G8222,G8223,G8224,G8225,G8226,G8227,G8228,G8229,G8230,G8231,G8232,G8233,G8234,G8235,G8236,G8237,G8238,G8239,G8240,
       G8241,G8242,G8243,G8244,G8245,G8246,G8247,G8248,G8249,G8250,G8251,G8252,G8253,G8254,G8255,G8256,G8257,G8258,G8259,G8260,
       G8261,G8262,G8263,G8264,G8265,G8266,G8267,G8268,G8269,G8270,G8271,G8272,G8273,G8274,G8275,G8276,G8277,G8278,G8279,G8280,
       G8281,G8282,G8283,G8284,G8285,G8286,G8287,G8288,G8289,G8290,G8291,G8292,G8293,G8294,G8295,G8296,G8297,G8298,G8299,G8300,
       G8301,G8302,G8303,G8304,G8305,G8306,G8307,G8308,G8309,G8310,G8311,G8312,G8313,G8314,G8315,G8316,G8317,G8318,G8319,G8320,
       G8321,G8322,G8323,G8324,G8325,G8326,G8327,G8328,G8329,G8330,G8331,G8332,G8333,G8334,G8335,G8336,G8337,G8338,G8339,G8340,
       G8341,G8342,G8343,G8344,G8345,G8346,G8347,G8348,G8349,G8350,G8351,G8352,G8353,G8354,G8355,G8356,G8357,G8358,G8359,G8360,
       G8361,G8362,G8363,G8364,G8365,G8366,G8367,G8368,G8369,G8370,G8371,G8372,G8373,G8374,G8375,G8376,G8377,G8378,G8379,G8380,
       G8381,G8382,G8383,G8384,G8385,G8386,G8387,G8388,G8389,G8390,G8391,G8392,G8393,G8394,G8395,G8396,G8397,G8398,G8399,G8400,
       G8401,G8402,G8403,G8404,G8405,G8406,G8407,G8408,G8409,G8410,G8411,G8412,G8413,G8414,G8415,G8416,G8417,G8418,G8419,G8420,
       G8421,G8422,G8423,G8424,G8425,G8426,G8427,G8428,G8429,G8430,G8431,G8432,G8433,G8434,G8435,G8436,G8437,G8438,G8439,G8440,
       G8441,G8442,G8443,G8444,G8445,G8446,G8447,G8448,G8449,G8450,G8451,G8452,G8453,G8454,G8455,G8456,G8457,G8458,G8459,G8460,
       G8461,G8462,G8463,G8464,G8465,G8466,G8467,G8468,G8469,G8470,G8471,G8472,G8473,G8474,G8475,G8476,G8477,G8478,G8479,G8480,
       G8481,G8482,G8483,G8484,G8485,G8486,G8487,G8488,G8489,G8490,G8491,G8492,G8493,G8494,G8495,G8496,G8497,G8498,G8499,G8500,
       G8501,G8502,G8503,G8504,G8505,G8506,G8507,G8508,G8509,G8510,G8511,G8512,G8513,G8514,G8515,G8516,G8517,G8518,G8519,G8520,
       G8521,G8522,G8523,G8524,G8525,G8526,G8527,G8528,G8529,G8530,G8531,G8532,G8533,G8534,G8535,G8536,G8537,G8538,G8539,G8540,
       G8541,G8542,G8543,G8544,G8545,G8546,G8547,G8548,G8549,G8550,G8551,G8552,G8553,G8554,G8555,G8556,G8557,G8558,G8559,G8560,
       G8561,G8562,G8563,G8564,G8565,G8566,G8567,G8568,G8569,G8570,G8571,G8572,G8573,G8574,G8575,G8576,G8577,G8578,G8579,G8580,
       G8581,G8582,G8583,G8584,G8585,G8586,G8587,G8588,G8589,G8590,G8591,G8592,G8593,G8594,G8595,G8596,G8597,G8598,G8599,G8600,
       G8601,G8602,G8603,G8604,G8605,G8606,G8607,G8608,G8609,G8610,G8611,G8612,G8613,G8614,G8615,G8616,G8617,G8618,G8619,G8620,
       G8621,G8622,G8623,G8624,G8625,G8626,G8627,G8628,G8629,G8630,G8631,G8632,G8633,G8634,G8635,G8636,G8637,G8638,G8639,G8640,
       G8641,G8642,G8643,G8644,G8645,G8646,G8647,G8648,G8649,G8650,G8651,G8652,G8653,G8654,G8655,G8656,G8657,G8658,G8659,G8660,
       G8661,G8662,G8663,G8664,G8665,G8666,G8667,G8668,G8669,G8670,G8671,G8672,G8673,G8674,G8675,G8676,G8677,G8678,G8679,G8680,
       G8681,G8682,G8683,G8684,G8685,G8686,G8687,G8688,G8689,G8690,G8691,G8692,G8693,G8694,G8695,G8696,G8697,G8698,G8699,G8700,
       G8701,G8702,G8703,G8704,G8705,G8706,G8707,G8708,G8709,G8710,G8711,G8712,G8713,G8714,G8715,G8716,G8717,G8718,G8719,G8720,
       G8721,G8722,G8723,G8724,G8725,G8726,G8727,G8728,G8729,G8730,G8731,G8732,G8733,G8734,G8735,G8736,G8737,G8738,G8739,G8740,
       G8741,G8742,G8743,G8744,G8745,G8746,G8747,G8748,G8749,G8750,G8751,G8752,G8753,G8754,G8755,G8756,G8757,G8758,G8759,G8760,
       G8761,G8762,G8763,G8764,G8765,G8766,G8767,G8768,G8769,G8770,G8771,G8772,G8773,G8774,G8775,G8776,G8777,G8778,G8779,G8780,
       G8781,G8782,G8783,G8784,G8785,G8786,G8787,G8788,G8789,G8790,G8791,G8792,G8793,G8794,G8795,G8796,G8797,G8798,G8799,G8800,
       G8801,G8802,G8803,G8804,G8805,G8806,G8807,G8808,G8809,G8810,G8811,G8812,G8813,G8814,G8815,G8816,G8817,G8818,G8819,G8820,
       G8821,G8822,G8823,G8824,G8825,G8826,G8827,G8828,G8829,G8830,G8831,G8832,G8833,G8834,G8835,G8836,G8837,G8838,G8839,G8840,
       G8841,G8842,G8843,G8844,G8845,G8846,G8847,G8848,G8849,G8850,G8851,G8852,G8853,G8854,G8855,G8856,G8857,G8858,G8859,G8860,
       G8861,G8862,G8863,G8864,G8865,G8866,G8867,G8868,G8869,G8870,G8871,G8872,G8873,G8874,G8875,G8876,G8877,G8878,G8879,G8880,
       G8881,G8882,G8883,G8884,G8885,G8886,G8887,G8888,G8889,G8890,G8891,G8892,G8893,G8894,G8895,G8896,G8897,G8898,G8899,G8900,
       G8901,G8902,G8903,G8904,G8905,G8906,G8907,G8908,G8909,G8910,G8911,G8912,G8913,G8914,G8915,G8916,G8917,G8918,G8919,G8920,
       G8921,G8922,G8923,G8924,G8925,G8926,G8927,G8928,G8929,G8930,G8931,G8932,G8933,G8934,G8935,G8936,G8937,G8938,G8939,G8940,
       G8941,G8942,G8943,G8944,G8945,G8946,G8947,G8948,G8949,G8950,G8951,G8952,G8953,G8954,G8955,G8956,G8957,G8958,G8959,G8960,
       G8961,G8962,G8963,G8964,G8965,G8966,G8967,G8968,G8969,G8970,G8971,G8972,G8973,G8974,G8975,G8976,G8977,G8978,G8979,G8980,
       G8981,G8982,G8983,G8984,G8985,G8986,G8987,G8988,G8989,G8990,G8991,G8992,G8993,G8994,G8995,G8996,G8997,G8998,G8999,G9000,
       G9001,G9002,G9003,G9004,G9005,G9006,G9007,G9008,G9009,G9010,G9011,G9012,G9013,G9014,G9015,G9016,G9017,G9018,G9019,G9020,
       G9021,G9022,G9023,G9024,G9025,G9026,G9027,G9028,G9029,G9030,G9031,G9032,G9033,G9034,G9035,G9036,G9037,G9038,G9039,G9040,
       G9041,G9042,G9043,G9044,G9045,G9046,G9047,G9048,G9049,G9050,G9051,G9052,G9053,G9054,G9055,G9056,G9057,G9058,G9059,G9060,
       G9061,G9062,G9063,G9064,G9065,G9066,G9067,G9068,G9069,G9070,G9071,G9072,G9073,G9074,G9075,G9076,G9077,G9078,G9079,G9080,
       G9081,G9082,G9083,G9084,G9085,G9086,G9087,G9088,G9089,G9090,G9091,G9092,G9093,G9094,G9095,G9096,G9097,G9098,G9099,G9100,
       G9101,G9102,G9103,G9104,G9105,G9106,G9107,G9108,G9109,G9110,G9111,G9112,G9113,G9114,G9115,G9116,G9117,G9118,G9119,G9120,
       G9121,G9122,G9123,G9124,G9125,G9126,G9127,G9128,G9129,G9130,G9131,G9132,G9133,G9134,G9135,G9136,G9137,G9138,G9139,G9140,
       G9141,G9142,G9143,G9144,G9145,G9146,G9147,G9148,G9149,G9150,G9151,G9152,G9153,G9154,G9155,G9156,G9157,G9158,G9159,G9160,
       G9161,G9162,G9163,G9164,G9165,G9166,G9167,G9168,G9169,G9170,G9171,G9172,G9173,G9174,G9175,G9176,G9177,G9178,G9179,G9180,
       G9181,G9182,G9183,G9184,G9185,G9186,G9187,G9188,G9189,G9190,G9191,G9192,G9193,G9194,G9195,G9196,G9197,G9198,G9199,G9200,
       G9201,G9202,G9203,G9204,G9205,G9206,G9207,G9208,G9209,G9210,G9211,G9212,G9213,G9214,G9215,G9216,G9217,G9218,G9219,G9220,
       G9221,G9222,G9223,G9224,G9225,G9226,G9227,G9228,G9229,G9230,G9231,G9232,G9233,G9234,G9235,G9236,G9237,G9238,G9239,G9240,
       G9241,G9242,G9243,G9244,G9245,G9246,G9247,G9248,G9249,G9250,G9251,G9252,G9253,G9254,G9255,G9256,G9257,G9258,G9259,G9260,
       G9261,G9262,G9263,G9264,G9265,G9266,G9267,G9268,G9269,G9270,G9271,G9272,G9273,G9274,G9275,G9276,G9277,G9278,G9279,G9280,
       G9281,G9282,G9283,G9284,G9285,G9286,G9287,G9288,G9289,G9290,G9291,G9292,G9293,G9294,G9295,G9296,G9297,G9298,G9299,G9300,
       G9301,G9302,G9303,G9304,G9305,G9306,G9307,G9308,G9309,G9310,G9311,G9312,G9313,G9314,G9315,G9316,G9317,G9318,G9319,G9320,
       G9321,G9322,G9323,G9324,G9325,G9326,G9327,G9328,G9329,G9330,G9331,G9332,G9333,G9334,G9335,G9336,G9337,G9338,G9339,G9340,
       G9341,G9342,G9343,G9344,G9345,G9346,G9347,G9348,G9349,G9350,G9351,G9352,G9353,G9354,G9355,G9356,G9357,G9358,G9359,G9360,
       G9361,G9362,G9363,G9364,G9365,G9366,G9367,G9368,G9369,G9370,G9371,G9372,G9373,G9374,G9375,G9376,G9377,G9378,G9379,G9380,
       G9381,G9382,G9383,G9384,G9385,G9386,G9387,G9388,G9389,G9390,G9391,G9392,G9393,G9394,G9395,G9396,G9397,G9398,G9399,G9400,
       G9401,G9402,G9403,G9404,G9405,G9406,G9407,G9408,G9409,G9410,G9411,G9412,G9413,G9414,G9415,G9416,G9417,G9418,G9419,G9420,
       G9421,G9422,G9423,G9424,G9425,G9426,G9427,G9428,G9429,G9430,G9431,G9432,G9433,G9434,G9435,G9436,G9437,G9438,G9439,G9440,
       G9441,G9442,G9443,G9444,G9445,G9446,G9447,G9448,G9449,G9450,G9451,G9452,G9453,G9454,G9455,G9456,G9457,G9458,G9459,G9460,
       G9461,G9462,G9463,G9464,G9465,G9466,G9467,G9468,G9469,G9470,G9471,G9472,G9473,G9474,G9475,G9476,G9477,G9478,G9479,G9480,
       G9481,G9482,G9483,G9484,G9485,G9486,G9487,G9488,G9489,G9490,G9491,G9492,G9493,G9494,G9495,G9496,G9497,G9498,G9499,G9500,
       G9501,G9502,G9503,G9504,G9505,G9506,G9507,G9508,G9509,G9510,G9511,G9512,G9513,G9514,G9515,G9516,G9517,G9518,G9519,G9520,
       G9521,G9522,G9523,G9524,G9525,G9526,G9527,G9528,G9529,G9530,G9531,G9532,G9533,G9534,G9535,G9536,G9537,G9538,G9539,G9540,
       G9541,G9542,G9543,G9544,G9545,G9546,G9547,G9548,G9549,G9550,G9551,G9552,G9553,G9554,G9555,G9556,G9557,G9558,G9559,G9560,
       G9561,G9562,G9563,G9564,G9565,G9566,G9567,G9568,G9569,G9570,G9571,G9572,G9573,G9574,G9575,G9576,G9577,G9578,G9579,G9580,
       G9581,G9582,G9583,G9584,G9585,G9586,G9587,G9588,G9589,G9590,G9591,G9592,G9593,G9594,G9595,G9596,G9597,G9598,G9599,G9600,
       G9601,G9602,G9603,G9604,G9605,G9606,G9607,G9608,G9609,G9610,G9611,G9612,G9613,G9614,G9615,G9616,G9617,G9618,G9619,G9620,
       G9621,G9622,G9623,G9624,G9625,G9626,G9627,G9628,G9629,G9630,G9631,G9632,G9633,G9634,G9635,G9636,G9637,G9638,G9639,G9640,
       G9641,G9642,G9643,G9644,G9645,G9646,G9647,G9648,G9649,G9650,G9651,G9652,G9653,G9654,G9655,G9656,G9657,G9658,G9659,G9660,
       G9661,G9662,G9663,G9664,G9665,G9666,G9667,G9668,G9669,G9670,G9671,G9672,G9673,G9674,G9675,G9676,G9677,G9678,G9679,G9680,
       G9681,G9682,G9683,G9684,G9685,G9686,G9687,G9688,G9689,G9690,G9691,G9692,G9693,G9694,G9695,G9696,G9697,G9698,G9699,G9700,
       G9701,G9702,G9703,G9704,G9705,G9706,G9707,G9708,G9709,G9710,G9711,G9712,G9713,G9714,G9715,G9716,G9717,G9718,G9719,G9720,
       G9721,G9722,G9723,G9724,G9725,G9726,G9727,G9728,G9729,G9730,G9731,G9732,G9733,G9734,G9735,G9736,G9737,G9738,G9739,G9740,
       G9741,G9742,G9743,G9744,G9745,G9746,G9747,G9748,G9749,G9750,G9751,G9752,G9753,G9754,G9755,G9756,G9757,G9758,G9759,G9760,
       G9761,G9762,G9763,G9764,G9765,G9766,G9767,G9768,G9769,G9770,G9771,G9772,G9773,G9774,G9775,G9776,G9777,G9778,G9779,G9780,
       G9781,G9782,G9783,G9784,G9785,G9786,G9787,G9788,G9789,G9790,G9791,G9792,G9793,G9794,G9795,G9796,G9797,G9798,G9799,G9800,
       G9801,G9802,G9803,G9804,G9805,G9806,G9807,G9808,G9809,G9810,G9811,G9812,G9813,G9814,G9815,G9816,G9817,G9818,G9819,G9820,
       G9821,G9822,G9823,G9824,G9825,G9826,G9827,G9828,G9829,G9830,G9831,G9832,G9833,G9834,G9835,G9836,G9837,G9838,G9839,G9840,
       G9841,G9842,G9843,G9844,G9845,G9846,G9847,G9848,G9849,G9850,G9851,G9852,G9853,G9854,G9855,G9856,G9857,G9858,G9859,G9860,
       G9861,G9862,G9863,G9864,G9865,G9866,G9867,G9868,G9869,G9870,G9871,G9872,G9873,G9874,G9875,G9876,G9877,G9878,G9879,G9880,
       G9881,G9882,G9883,G9884,G9885,G9886,G9887,G9888,G9889,G9890,G9891,G9892,G9893,G9894,G9895,G9896,G9897,G9898,G9899,G9900,
       G9901,G9902,G9903,G9904,G9905,G9906,G9907,G9908,G9909,G9910,G9911,G9912,G9913,G9914,G9915,G9916,G9917,G9918,G9919,G9920,
       G9921,G9922,G9923,G9924,G9925,G9926,G9927,G9928,G9929,G9930,G9931,G9932,G9933,G9934,G9935,G9936,G9937,G9938,G9939,G9940,
       G9941,G9942,G9943,G9944,G9945,G9946,G9947,G9948,G9949,G9950,G9951,G9952,G9953,G9954,G9955,G9956,G9957,G9958,G9959,G9960,
       G9961,G9962,G9963,G9964,G9965,G9966,G9967,G9968,G9969,G9970,G9971,G9972,G9973,G9974,G9975,G9976,G9977,G9978,G9979,G9980,
       G9981,G9982,G9983,G9984,G9985,G9986,G9987,G9988,G9989,G9990,G9991,G9992,G9993,G9994,G9995,G9996,G9997,G9998,G9999,G10000,
       G10001,G10002,G10003,G10004,G10005,G10006,G10007,G10008,G10009,G10010,G10011,G10012,G10013,G10014,G10015,G10016,G10017,G10018,G10019,G10020,
       G10021,G10022,G10023,G10024,G10025,G10026,G10027,G10028,G10029,G10030,G10031,G10032,G10033,G10034,G10035,G10036,G10037,G10038,G10039,G10040,
       G10041,G10042,G10043,G10044,G10045,G10046,G10047,G10048,G10049,G10050,G10051,G10052,G10053,G10054,G10055,G10056,G10057,G10058,G10059,G10060,
       G10061,G10062,G10063,G10064,G10065,G10066,G10067,G10068,G10069,G10070,G10071,G10072,G10073,G10074,G10075,G10076,G10077,G10078,G10079,G10080,
       G10081,G10082,G10083,G10084,G10085,G10086,G10087,G10088,G10089,G10090,G10091,G10092,G10093,G10094,G10095,G10096,G10097,G10098,G10099,G10100,
       G10101,G10102,G10103,G10104,G10105,G10106,G10107,G10108,G10109,G10110,G10111,G10112,G10113,G10114,G10115,G10116,G10117,G10118,G10119,G10120,
       G10121,G10122,G10123,G10124,G10125,G10126,G10127,G10128,G10129,G10130,G10131,G10132,G10133,G10134,G10135,G10136,G10137,G10138,G10139,G10140,
       G10141,G10142,G10143,G10144,G10145,G10146,G10147,G10148,G10149,G10150,G10151,G10152,G10153,G10154,G10155,G10156,G10157,G10158,G10159,G10160,
       G10161,G10162,G10163,G10164,G10165,G10166,G10167,G10168,G10169,G10170,G10171,G10172,G10173,G10174,G10175,G10176,G10177,G10178,G10179,G10180,
       G10181,G10182,G10183,G10184,G10185,G10186,G10187,G10188,G10189,G10190,G10191,G10192,G10193,G10194,G10195,G10196,G10197,G10198,G10199,G10200,
       G10201,G10202,G10203,G10204,G10205,G10206,G10207,G10208,G10209,G10210,G10211,G10212,G10213,G10214,G10215,G10216,G10217,G10218,G10219,G10220,
       G10221,G10222,G10223,G10224,G10225,G10226,G10227,G10228,G10229,G10230,G10231,G10232,G10233,G10234,G10235,G10236,G10237,G10238,G10239,G10240,
       G10241,G10242,G10243,G10244,G10245,G10246,G10247,G10248,G10249,G10250,G10251,G10252,G10253,G10254,G10255,G10256,G10257,G10258,G10259,G10260,
       G10261,G10262,G10263,G10264,G10265,G10266,G10267,G10268,G10269,G10270,G10271,G10272,G10273,G10274,G10275,G10276,G10277,G10278,G10279,G10280,
       G10281,G10282,G10283,G10284,G10285,G10286,G10287,G10288,G10289,G10290,G10291,G10292,G10293,G10294,G10295,G10296,G10297,G10298,G10299,G10300,
       G10301,G10302,G10303,G10304,G10305,G10306,G10307,G10308,G10309,G10310,G10311,G10312,G10313,G10314,G10315,G10316,G10317,G10318,G10319,G10320,
       G10321,G10322,G10323,G10324,G10325,G10326,G10327,G10328,G10329,G10330,G10331,G10332,G10333,G10334,G10335,G10336,G10337,G10338,G10339,G10340,
       G10341,G10342,G10343,G10344,G10345,G10346,G10347,G10348,G10349,G10350,G10351,G10352,G10353,G10354,G10355,G10356,G10357,G10358,G10359,G10360,
       G10361,G10362,G10363,G10364,G10365,G10366,G10367,G10368,G10369,G10370,G10371,G10372,G10373,G10374,G10375,G10376,G10377,G10378,G10379,G10380,
       G10381,G10382,G10383,G10384,G10385,G10386,G10387,G10388,G10389,G10390,G10391,G10392,G10393,G10394,G10395,G10396,G10397,G10398,G10399,G10400,
       G10401,G10402,G10403,G10404,G10405,G10406,G10407,G10408,G10409,G10410,G10411,G10412,G10413,G10414,G10415,G10416,G10417,G10418,G10419,G10420,
       G10421,G10422,G10423,G10424,G10425,G10426,G10427,G10428,G10429,G10430,G10431,G10432,G10433,G10434,G10435,G10436,G10437,G10438,G10439,G10440,
       G10441,G10442,G10443,G10444,G10445,G10446,G10447,G10448,G10449,G10450,G10451,G10452,G10453,G10454,G10455,G10456,G10457,G10458,G10459,G10460,
       G10461,G10462,G10463,G10464,G10465,G10466,G10467,G10468,G10469,G10470,G10471,G10472,G10473,G10474,G10475,G10476,G10477,G10478,G10479,G10480,
       G10481,G10482,G10483,G10484,G10485,G10486,G10487,G10488,G10489,G10490,G10491,G10492,G10493,G10494,G10495,G10496,G10497,G10498,G10499,G10500,
       G10501,G10502,G10503,G10504,G10505,G10506,G10507,G10508,G10509,G10510,G10511,G10512,G10513,G10514,G10515,G10516,G10517,G10518,G10519,G10520,
       G10521,G10522,G10523,G10524,G10525,G10526,G10527,G10528,G10529,G10530,G10531,G10532,G10533,G10534,G10535,G10536,G10537,G10538,G10539,G10540,
       G10541,G10542,G10543,G10544,G10545,G10546,G10547,G10548,G10549,G10550,G10551,G10552,G10553,G10554,G10555,G10556,G10557,G10558,G10559,G10560,
       G10561,G10562,G10563,G10564,G10565,G10566,G10567,G10568,G10569,G10570,G10571,G10572,G10573,G10574,G10575,G10576,G10577,G10578,G10579,G10580,
       G10581,G10582,G10583,G10584,G10585,G10586,G10587,G10588,G10589,G10590,G10591,G10592,G10593,G10594,G10595,G10596,G10597,G10598,G10599,G10600,
       G10601,G10602,G10603,G10604,G10605,G10606,G10607,G10608,G10609,G10610,G10611,G10612,G10613,G10614,G10615,G10616,G10617,G10618,G10619,G10620,
       G10621,G10622,G10623,G10624,G10625,G10626,G10627,G10628,G10629,G10630,G10631,G10632,G10633,G10634,G10635,G10636,G10637,G10638,G10639,G10640,
       G10641,G10642,G10643,G10644,G10645,G10646,G10647,G10648,G10649,G10650,G10651,G10652,G10653,G10654,G10655,G10656,G10657,G10658,G10659,G10660,
       G10661,G10662,G10663,G10664,G10665,G10666,G10667,G10668,G10669,G10670,G10671,G10672,G10673,G10674,G10675,G10676,G10677,G10678,G10679,G10680,
       G10681,G10682,G10683,G10684,G10685,G10686,G10687,G10688,G10689,G10690,G10691,G10692,G10693,G10694,G10695,G10696,G10697,G10698,G10699,G10700,
       G10701,G10702,G10703,G10704,G10705,G10706,G10707,G10708,G10709,G10710,G10711,G10712,G10713,G10714,G10715,G10716,G10717,G10718,G10719,G10720,
       G10721,G10722,G10723,G10724,G10725,G10726,G10727,G10728,G10729,G10730,G10731,G10732,G10733,G10734,G10735,G10736,G10737,G10738,G10739,G10740,
       G10741,G10742,G10743,G10744,G10745,G10746,G10747,G10748,G10749,G10750,G10751,G10752,G10753,G10754,G10755,G10756,G10757,G10758,G10759,G10760,
       G10761,G10762,G10763,G10764,G10765,G10766,G10767,G10768,G10769,G10770,G10771,G10772,G10773,G10774,G10775,G10776,G10777,G10778,G10779,G10780,
       G10781,G10782,G10783,G10784,G10785,G10786,G10787,G10788,G10789,G10790,G10791,G10792,G10793,G10794,G10795,G10796,G10797,G10798,G10799,G10800,
       G10801,G10802,G10803,G10804,G10805,G10806,G10807,G10808,G10809,G10810,G10811,G10812,G10813,G10814,G10815,G10816,G10817,G10818,G10819,G10820,
       G10821,G10822,G10823,G10824,G10825,G10826,G10827,G10828,G10829,G10830,G10831,G10832,G10833,G10834,G10835,G10836,G10837,G10838,G10839,G10840,
       G10841,G10842,G10843,G10844,G10845,G10846,G10847,G10848,G10849,G10850,G10851,G10852,G10853,G10854,G10855,G10856,G10857,G10858,G10859,G10860,
       G10861,G10862,G10863,G10864,G10865,G10866,G10867,G10868,G10869,G10870,G10871,G10872,G10873,G10874,G10875,G10876,G10877,G10878,G10879,G10880,
       G10881,G10882,G10883,G10884,G10885,G10886,G10887,G10888,G10889,G10890,G10891,G10892,G10893,G10894,G10895,G10896,G10897,G10898,G10899,G10900,
       G10901,G10902,G10903,G10904,G10905,G10906,G10907,G10908,G10909,G10910,G10911,G10912,G10913,G10914,G10915,G10916,G10917,G10918,G10919,G10920,
       G10921,G10922,G10923,G10924,G10925,G10926,G10927,G10928,G10929,G10930,G10931,G10932,G10933,G10934,G10935,G10936,G10937,G10938,G10939,G10940,
       G10941,G10942,G10943,G10944,G10945,G10946,G10947,G10948,G10949,G10950,G10951,G10952,G10953,G10954,G10955,G10956,G10957,G10958,G10959,G10960,
       G10961,G10962,G10963,G10964,G10965,G10966,G10967,G10968,G10969,G10970,G10971,G10972,G10973,G10974,G10975,G10976,G10977,G10978,G10979,G10980,
       G10981,G10982,G10983,G10984,G10985,G10986,G10987,G10988,G10989,G10990,G10991,G10992,G10993,G10994,G10995,G10996,G10997,G10998,G10999,G11000,
       G11001,G11002,G11003,G11004,G11005,G11006,G11007,G11008,G11009,G11010,G11011,G11012,G11013,G11014,G11015,G11016,G11017,G11018,G11019,G11020,
       G11021,G11022,G11023,G11024,G11025,G11026,G11027,G11028,G11029,G11030,G11031,G11032,G11033,G11034,G11035,G11036,G11037,G11038,G11039,G11040,
       G11041,G11042,G11043,G11044,G11045,G11046,G11047,G11048,G11049,G11050,G11051,G11052,G11053,G11054,G11055,G11056,G11057,G11058,G11059,G11060,
       G11061,G11062,G11063,G11064,G11065,G11066,G11067,G11068,G11069,G11070,G11071,G11072,G11073,G11074,G11075,G11076,G11077,G11078,G11079,G11080,
       G11081,G11082,G11083,G11084,G11085,G11086,G11087,G11088,G11089,G11090,G11091,G11092,G11093,G11094,G11095,G11096,G11097,G11098,G11099,G11100,
       G11101,G11102,G11103,G11104,G11105,G11106,G11107,G11108,G11109,G11110,G11111,G11112,G11113,G11114,G11115,G11116,G11117,G11118,G11119,G11120,
       G11121,G11122,G11123,G11124,G11125,G11126,G11127,G11128,G11129,G11130,G11131,G11132,G11133,G11134,G11135,G11136,G11137,G11138,G11139,G11140,
       G11141,G11142,G11143,G11144,G11145,G11146,G11147,G11148,G11149,G11150,G11151,G11152,G11153,G11154,G11155,G11156,G11157,G11158,G11159,G11160,
       G11161,G11162,G11163,G11164,G11165,G11166,G11167,G11168,G11169,G11170,G11171,G11172,G11173,G11174,G11175,G11176,G11177,G11178,G11179,G11180,
       G11181,G11182,G11183,G11184,G11185,G11186,G11187,G11188,G11189,G11190,G11191,G11192,G11193,G11194,G11195,G11196,G11197,G11198,G11199,G11200,
       G11201,G11202,G11203,G11204,G11205,G11206,G11207,G11208,G11209,G11210,G11211,G11212,G11213,G11214,G11215,G11216,G11217,G11218,G11219,G11220,
       G11221,G11222,G11223,G11224,G11225,G11226,G11227,G11228,G11229,G11230,G11231,G11232,G11233,G11234,G11235,G11236,G11237,G11238,G11239,G11240,
       G11241,G11242,G11243,G11244,G11245,G11246,G11247,G11248,G11249,G11250,G11251,G11252,G11253,G11254,G11255,G11256,G11257,G11258,G11259,G11260,
       G11261,G11262,G11263,G11264,G11265,G11266,G11267,G11268,G11269,G11270,G11271,G11272,G11273,G11274,G11275,G11276,G11277,G11278,G11279,G11280,
       G11281,G11282,G11283,G11284,G11285,G11286,G11287,G11288,G11289,G11290,G11291,G11292,G11293,G11294,G11295,G11296,G11297,G11298,G11299,G11300,
       G11301,G11302,G11303,G11304,G11305,G11306,G11307,G11308,G11309,G11310,G11311,G11312,G11313,G11314,G11315,G11316,G11317,G11318,G11319,G11320,
       G11321,G11322,G11323,G11324,G11325,G11326,G11327,G11328,G11329,G11330,G11331,G11332,G11333,G11334,G11335,G11336,G11337,G11338,G11339,G11340,
       G11341,G11342,G11343,G11344,G11345,G11346,G11347,G11348,G11349,G11350,G11351,G11352,G11353,G11354,G11355,G11356,G11357,G11358,G11359,G11360,
       G11361,G11362,G11363,G11364,G11365,G11366,G11367,G11368,G11369,G11370,G11371,G11372,G11373,G11374,G11375,G11376,G11377,G11378,G11379,G11380,
       G11381,G11382,G11383,G11384,G11385,G11386,G11387,G11388,G11389,G11390,G11391,G11392,G11393,G11394,G11395,G11396,G11397,G11398,G11399,G11400,
       G11401,G11402,G11403,G11404,G11405,G11406,G11407,G11408,G11409,G11410,G11411,G11412,G11413,G11414,G11415,G11416,G11417,G11418,G11419,G11420,
       G11421,G11422,G11423,G11424,G11425,G11426,G11427,G11428,G11429,G11430,G11431,G11432,G11433,G11434,G11435,G11436,G11437,G11438,G11439,G11440,
       G11441,G11442,G11443,G11444,G11445,G11446,G11447,G11448,G11449,G11450,G11451,G11452,G11453,G11454,G11455,G11456,G11457,G11458,G11459,G11460,
       G11461,G11462,G11463,G11464,G11465,G11466,G11467,G11468,G11469,G11470,G11471,G11472,G11473,G11474,G11475,G11476,G11477,G11478,G11479,G11480,
       G11481,G11482,G11483,G11484,G11485,G11486,G11487,G11488,G11489,G11490,G11491,G11492,G11493,G11494,G11495,G11496,G11497,G11498,G11499,G11500,
       G11501,G11502,G11503,G11504,G11505,G11506,G11507,G11508,G11509,G11510,G11511,G11512,G11513,G11514,G11515,G11516,G11517,G11518,G11519,G11520,
       G11521,G11522,G11523,G11524,G11525,G11526,G11527,G11528,G11529,G11530,G11531,G11532,G11533,G11534,G11535,G11536,G11537,G11538,G11539,G11540,
       G11541,G11542,G11543,G11544,G11545,G11546,G11547,G11548,G11549,G11550,G11551,G11552,G11553,G11554,G11555,G11556,G11557,G11558,G11559,G11560,
       G11561,G11562,G11563,G11564,G11565,G11566,G11567,G11568,G11569,G11570,G11571,G11572,G11573,G11574,G11575,G11576,G11577,G11578,G11579,G11580,
       G11581,G11582,G11583,G11584,G11585,G11586,G11587,G11588,G11589,G11590,G11591,G11592,G11593,G11594,G11595,G11596,G11597,G11598,G11599,G11600,
       G11601,G11602,G11603,G11604,G11605,G11606,G11607,G11608,G11609,G11610,G11611,G11612,G11613,G11614,G11615,G11616,G11617,G11618,G11619,G11620,
       G11621,G11622,G11623,G11624,G11625,G11626,G11627,G11628,G11629,G11630,G11631,G11632,G11633,G11634,G11635,G11636,G11637,G11638,G11639,G11640,
       G11641,G11642,G11643,G11644,G11645,G11646,G11647,G11648,G11649,G11650,G11651,G11652,G11653,G11654,G11655,G11656,G11657,G11658,G11659,G11660,
       G11661,G11662,G11663,G11664,G11665,G11666,G11667,G11668,G11669,G11670,G11671,G11672,G11673,G11674,G11675,G11676,G11677,G11678,G11679,G11680,
       G11681,G11682,G11683,G11684,G11685,G11686,G11687,G11688,G11689,G11690,G11691,G11692,G11693,G11694,G11695,G11696,G11697,G11698,G11699,G11700,
       G11701,G11702,G11703,G11704,G11705,G11706,G11707,G11708,G11709,G11710,G11711,G11712,G11713,G11714,G11715,G11716,G11717,G11718,G11719,G11720,
       G11721,G11722,G11723,G11724,G11725,G11726,G11727,G11728,G11729,G11730,G11731,G11732,G11733,G11734,G11735,G11736,G11737,G11738,G11739,G11740,
       G11741,G11742,G11743,G11744,G11745,G11746,G11747,G11748,G11749,G11750,G11751,G11752,G11753,G11754,G11755,G11756,G11757,G11758,G11759,G11760,
       G11761,G11762,G11763,G11764,G11765,G11766,G11767,G11768,G11769,G11770,G11771,G11772,G11773,G11774,G11775,G11776,G11777,G11778,G11779,G11780,
       G11781,G11782,G11783,G11784,G11785,G11786,G11787,G11788,G11789,G11790,G11791,G11792,G11793,G11794,G11795,G11796,G11797,G11798,G11799,G11800,
       G11801,G11802,G11803,G11804,G11805,G11806,G11807,G11808,G11809,G11810,G11811,G11812,G11813,G11814,G11815,G11816,G11817,G11818,G11819,G11820,
       G11821,G11822,G11823,G11824,G11825,G11826,G11827,G11828,G11829,G11830,G11831,G11832,G11833,G11834,G11835,G11836,G11837,G11838,G11839,G11840,
       G11841,G11842,G11843,G11844,G11845,G11846,G11847,G11848,G11849,G11850,G11851,G11852,G11853,G11854,G11855,G11856,G11857,G11858,G11859,G11860,
       G11861,G11862,G11863,G11864,G11865,G11866,G11867,G11868,G11869,G11870,G11871,G11872,G11873,G11874,G11875,G11876,G11877,G11878,G11879,G11880,
       G11881,G11882,G11883,G11884,G11885,G11886,G11887,G11888,G11889,G11890,G11891,G11892,G11893,G11894,G11895,G11896,G11897,G11898,G11899,G11900,
       G11901,G11902,G11903,G11904,G11905,G11906,G11907,G11908,G11909,G11910,G11911,G11912,G11913,G11914,G11915,G11916,G11917,G11918,G11919,G11920,
       G11921,G11922,G11923,G11924,G11925,G11926,G11927,G11928,G11929,G11930,G11931,G11932,G11933,G11934,G11935,G11936,G11937,G11938,G11939,G11940,
       G11941,G11942,G11943,G11944,G11945,G11946,G11947,G11948,G11949,G11950,G11951,G11952,G11953,G11954,G11955,G11956,G11957,G11958,G11959,G11960,
       G11961,G11962,G11963,G11964,G11965,G11966,G11967,G11968,G11969,G11970,G11971,G11972,G11973,G11974,G11975,G11976,G11977,G11978,G11979,G11980,
       G11981,G11982,G11983,G11984,G11985,G11986,G11987,G11988,G11989,G11990,G11991,G11992,G11993,G11994,G11995,G11996,G11997,G11998,G11999,G12000,
       G12001,G12002,G12003,G12004,G12005,G12006,G12007,G12008,G12009,G12010,G12011,G12012,G12013,G12014,G12015,G12016,G12017,G12018,G12019,G12020,
       G12021,G12022,G12023,G12024,G12025,G12026,G12027,G12028,G12029,G12030,G12031,G12032,G12033,G12034,G12035,G12036,G12037,G12038,G12039,G12040,
       G12041,G12042,G12043,G12044,G12045,G12046,G12047,G12048,G12049,G12050,G12051,G12052,G12053,G12054,G12055,G12056,G12057,G12058,G12059,G12060,
       G12061,G12062,G12063,G12064,G12065,G12066,G12067,G12068,G12069,G12070,G12071,G12072,G12073,G12074,G12075,G12076,G12077,G12078,G12079,G12080,
       G12081,G12082,G12083,G12084,G12085,G12086,G12087,G12088,G12089,G12090,G12091,G12092,G12093,G12094,G12095,G12096,G12097,G12098,G12099,G12100,
       G12101,G12102,G12103,G12104,G12105,G12106,G12107,G12108,G12109,G12110,G12111,G12112,G12113,G12114,G12115,G12116,G12117,G12118,G12119,G12120,
       G12121,G12122,G12123,G12124,G12125,G12126,G12127,G12128,G12129,G12130,G12131,G12132,G12133,G12134,G12135,G12136,G12137,G12138,G12139,G12140,
       G12141,G12142,G12143,G12144,G12145,G12146,G12147,G12148,G12149,G12150,G12151,G12152,G12153,G12154,G12155,G12156,G12157,G12158,G12159,G12160,
       G12161,G12162,G12163,G12164,G12165,G12166,G12167,G12168,G12169,G12170,G12171,G12172,G12173,G12174,G12175,G12176,G12177,G12178,G12179,G12180,
       G12181,G12182,G12183,G12184,G12185,G12186,G12187,G12188,G12189,G12190,G12191,G12192,G12193,G12194,G12195,G12196,G12197,G12198,G12199,G12200,
       G12201,G12202,G12203,G12204,G12205,G12206,G12207,G12208,G12209,G12210,G12211,G12212,G12213,G12214,G12215,G12216,G12217,G12218,G12219,G12220,
       G12221,G12222,G12223,G12224,G12225,G12226,G12227,G12228,G12229,G12230,G12231,G12232,G12233,G12234,G12235,G12236,G12237,G12238,G12239,G12240,
       G12241,G12242,G12243,G12244,G12245,G12246,G12247,G12248,G12249,G12250,G12251,G12252,G12253,G12254,G12255,G12256,G12257,G12258,G12259,G12260,
       G12261,G12262,G12263,G12264,G12265,G12266,G12267,G12268,G12269,G12270,G12271,G12272,G12273,G12274,G12275,G12276,G12277,G12278,G12279,G12280,
       G12281,G12282,G12283,G12284,G12285,G12286,G12287,G12288,G12289,G12290,G12291,G12292,G12293,G12294,G12295,G12296,G12297,G12298,G12299,G12300,
       G12301,G12302,G12303,G12304,G12305,G12306,G12307,G12308,G12309,G12310,G12311,G12312,G12313,G12314,G12315,G12316,G12317,G12318,G12319,G12320,
       G12321,G12322,G12323,G12324,G12325,G12326,G12327,G12328,G12329,G12330,G12331,G12332,G12333,G12334,G12335,G12336,G12337,G12338,G12339,G12340,
       G12341,G12342,G12343,G12344,G12345,G12346,G12347,G12348,G12349,G12350,G12351,G12352,G12353,G12354,G12355,G12356,G12357,G12358,G12359,G12360,
       G12361,G12362,G12363,G12364,G12365,G12366,G12367,G12368,G12369,G12370,G12371,G12372,G12373,G12374,G12375,G12376,G12377,G12378,G12379,G12380,
       G12381,G12382,G12383,G12384,G12385,G12386,G12387,G12388,G12389,G12390,G12391,G12392,G12393,G12394,G12395,G12396,G12397,G12398,G12399,G12400,
       G12401,G12402,G12403,G12404,G12405,G12406,G12407,G12408,G12409,G12410,G12411,G12412,G12413,G12414,G12415,G12416,G12417,G12418,G12419,G12420,
       G12421,G12422,G12423,G12424,G12425,G12426,G12427,G12428,G12429,G12430,G12431,G12432,G12433,G12434,G12435,G12436,G12437,G12438,G12439,G12440,
       G12441,G12442,G12443,G12444,G12445,G12446,G12447,G12448,G12449,G12450,G12451,G12452,G12453,G12454,G12455,G12456,G12457,G12458,G12459,G12460,
       G12461,G12462,G12463,G12464,G12465,G12466,G12467,G12468,G12469,G12470,G12471,G12472,G12473,G12474,G12475,G12476,G12477,G12478,G12479,G12480,
       G12481,G12482,G12483,G12484,G12485,G12486,G12487,G12488,G12489,G12490,G12491,G12492,G12493,G12494,G12495,G12496,G12497,G12498,G12499,G12500,
       G12501,G12502,G12503,G12504,G12505,G12506,G12507,G12508,G12509,G12510,G12511,G12512,G12513,G12514,G12515,G12516,G12517,G12518,G12519,G12520,
       G12521,G12522,G12523,G12524,G12525,G12526,G12527,G12528,G12529,G12530,G12531,G12532,G12533,G12534,G12535,G12536,G12537,G12538,G12539,G12540,
       G12541,G12542,G12543,G12544,G12545,G12546,G12547,G12548,G12549,G12550,G12551,G12552,G12553,G12554,G12555,G12556,G12557,G12558,G12559,G12560,
       G12561,G12562,G12563,G12564,G12565,G12566,G12567,G12568,G12569,G12570,G12571,G12572,G12573,G12574,G12575,G12576,G12577,G12578,G12579,G12580,
       G12581,G12582,G12583,G12584,G12585,G12586,G12587,G12588,G12589,G12590,G12591,G12592,G12593,G12594,G12595,G12596,G12597,G12598,G12599,G12600,
       G12601,G12602,G12603,G12604,G12605,G12606,G12607,G12608,G12609,G12610,G12611,G12612,G12613,G12614,G12615,G12616,G12617,G12618,G12619,G12620,
       G12621,G12622,G12623,G12624,G12625,G12626,G12627,G12628,G12629,G12630,G12631,G12632,G12633,G12634,G12635,G12636,G12637,G12638,G12639,G12640,
       G12641,G12642,G12643,G12644,G12645,G12646,G12647,G12648,G12649,G12650,G12651,G12652,G12653,G12654,G12655,G12656,G12657,G12658,G12659,G12660,
       G12661,G12662,G12663,G12664,G12665,G12666,G12667,G12668,G12669,G12670,G12671,G12672,G12673,G12674,G12675,G12676,G12677,G12678,G12679,G12680,
       G12681,G12682,G12683,G12684,G12685,G12686,G12687,G12688,G12689,G12690,G12691,G12692,G12693,G12694,G12695,G12696,G12697,G12698,G12699,G12700,
       G12701,G12702,G12703,G12704,G12705,G12706,G12707,G12708,G12709,G12710,G12711,G12712,G12713,G12714,G12715,G12716,G12717,G12718,G12719,G12720,
       G12721,G12722,G12723,G12724,G12725,G12726,G12727,G12728,G12729,G12730,G12731,G12732,G12733,G12734,G12735,G12736,G12737,G12738,G12739,G12740,
       G12741,G12742,G12743,G12744,G12745,G12746,G12747,G12748,G12749,G12750,G12751,G12752,G12753,G12754,G12755,G12756,G12757,G12758,G12759,G12760,
       G12761,G12762,G12763,G12764,G12765,G12766,G12767,G12768,G12769,G12770,G12771,G12772,G12773,G12774,G12775,G12776,G12777,G12778,G12779,G12780,
       G12781,G12782,G12783,G12784,G12785,G12786,G12787,G12788,G12789,G12790,G12791,G12792,G12793,G12794,G12795,G12796,G12797,G12798,G12799,G12800,
       G12801,G12802,G12803,G12804,G12805,G12806,G12807,G12808,G12809,G12810,G12811,G12812,G12813,G12814,G12815,G12816,G12817,G12818,G12819,G12820,
       G12821,G12822,G12823,G12824,G12825,G12826,G12827,G12828,G12829,G12830,G12831,G12832,G12833,G12834,G12835,G12836,G12837,G12838,G12839,G12840,
       G12841,G12842,G12843,G12844,G12845,G12846,G12847,G12848,G12849,G12850,G12851,G12852,G12853,G12854,G12855,G12856,G12857,G12858,G12859,G12860,
       G12861,G12862,G12863,G12864,G12865,G12866,G12867,G12868,G12869,G12870,G12871,G12872,G12873,G12874,G12875,G12876,G12877,G12878,G12879,G12880,
       G12881,G12882,G12883,G12884,G12885,G12886,G12887,G12888,G12889,G12890,G12891,G12892,G12893,G12894,G12895,G12896,G12897,G12898,G12899,G12900,
       G12901,G12902,G12903,G12904,G12905,G12906,G12907,G12908,G12909,G12910,G12911,G12912,G12913,G12914,G12915,G12916,G12917,G12918,G12919,G12920,
       G12921,G12922,G12923,G12924,G12925,G12926,G12927,G12928,G12929,G12930,G12931,G12932,G12933,G12934,G12935,G12936,G12937,G12938,G12939,G12940,
       G12941,G12942,G12943,G12944,G12945,G12946,G12947,G12948,G12949,G12950,G12951,G12952,G12953,G12954,G12955,G12956,G12957,G12958,G12959,G12960,
       G12961,G12962,G12963,G12964,G12965,G12966,G12967,G12968,G12969,G12970,G12971,G12972,G12973,G12974,G12975,G12976,G12977,G12978,G12979,G12980,
       G12981,G12982,G12983,G12984,G12985,G12986,G12987,G12988,G12989,G12990,G12991,G12992,G12993,G12994,G12995,G12996,G12997,G12998,G12999,G13000,
       G13001,G13002,G13003,G13004,G13005,G13006,G13007,G13008,G13009,G13010,G13011,G13012,G13013,G13014,G13015,G13016,G13017,G13018,G13019,G13020,
       G13021,G13022,G13023,G13024,G13025,G13026,G13027,G13028,G13029,G13030,G13031,G13032,G13033,G13034,G13035,G13036,G13037,G13038,G13039,G13040,
       G13041,G13042,G13043,G13044,G13045,G13046,G13047,G13048,G13049,G13050,G13051,G13052,G13053,G13054,G13055,G13056,G13057,G13058,G13059,G13060,
       G13061,G13062,G13063,G13064,G13065,G13066,G13067,G13068,G13069,G13070,G13071,G13072,G13073,G13074,G13075,G13076,G13077,G13078,G13079,G13080,
       G13081,G13082,G13083,G13084,G13085,G13086,G13087,G13088,G13089,G13090,G13091,G13092,G13093,G13094,G13095,G13096,G13097,G13098,G13099,G13100,
       G13101,G13102,G13103,G13104,G13105,G13106,G13107,G13108,G13109,G13110,G13111,G13112,G13113,G13114,G13115,G13116,G13117,G13118,G13119,G13120,
       G13121,G13122,G13123,G13124,G13125,G13126,G13127,G13128,G13129,G13130,G13131,G13132,G13133,G13134,G13135,G13136,G13137,G13138,G13139,G13140,
       G13141,G13142,G13143,G13144,G13145,G13146,G13147,G13148,G13149,G13150,G13151,G13152,G13153,G13154,G13155,G13156,G13157,G13158,G13159,G13160,
       G13161,G13162,G13163,G13164,G13165,G13166,G13167,G13168,G13169,G13170,G13171,G13172,G13173,G13174,G13175,G13176,G13177,G13178,G13179,G13180,
       G13181,G13182,G13183,G13184,G13185,G13186,G13187,G13188,G13189,G13190,G13191,G13192,G13193,G13194,G13195,G13196,G13197,G13198,G13199,G13200,
       G13201,G13202,G13203,G13204,G13205,G13206,G13207,G13208,G13209,G13210,G13211,G13212,G13213,G13214,G13215,G13216,G13217,G13218,G13219,G13220,
       G13221,G13222,G13223,G13224,G13225,G13226,G13227,G13228,G13229,G13230,G13231,G13232,G13233,G13234,G13235,G13236,G13237,G13238,G13239,G13240,
       G13241,G13242,G13243,G13244,G13245,G13246,G13247,G13248,G13249,G13250,G13251,G13252,G13253,G13254,G13255,G13256,G13257,G13258,G13259,G13260,
       G13261,G13262,G13263,G13264,G13265,G13266,G13267,G13268,G13269,G13270,G13271,G13272,G13273,G13274,G13275,G13276,G13277,G13278,G13279,G13280,
       G13281,G13282,G13283,G13284,G13285,G13286,G13287,G13288,G13289,G13290,G13291,G13292,G13293,G13294,G13295,G13296,G13297,G13298,G13299,G13300,
       G13301,G13302,G13303,G13304,G13305,G13306,G13307,G13308,G13309,G13310,G13311,G13312,G13313,G13314,G13315,G13316,G13317,G13318,G13319,G13320,
       G13321,G13322,G13323,G13324,G13325,G13326,G13327,G13328,G13329,G13330,G13331,G13332,G13333,G13334,G13335,G13336,G13337,G13338,G13339,G13340,
       G13341,G13342,G13343,G13344,G13345,G13346,G13347,G13348,G13349,G13350,G13351,G13352,G13353,G13354,G13355,G13356,G13357,G13358,G13359,G13360,
       G13361,G13362,G13363,G13364,G13365,G13366,G13367,G13368,G13369,G13370,G13371,G13372,G13373,G13374,G13375,G13376,G13377,G13378,G13379,G13380,
       G13381,G13382,G13383,G13384,G13385,G13386,G13387,G13388,G13389,G13390,G13391,G13392,G13393,G13394,G13395,G13396,G13397,G13398,G13399,G13400,
       G13401,G13402,G13403,G13404,G13405,G13406,G13407,G13408,G13409,G13410,G13411,G13412,G13413,G13414,G13415,G13416,G13417,G13418,G13419,G13420,
       G13421,G13422,G13423,G13424,G13425,G13426,G13427,G13428,G13429,G13430,G13431,G13432,G13433,G13434,G13435,G13436,G13437,G13438,G13439,G13440,
       G13441,G13442,G13443,G13444,G13445,G13446,G13447,G13448,G13449,G13450,G13451,G13452,G13453,G13454,G13455,G13456,G13457,G13458,G13459,G13460,
       G13461,G13462,G13463,G13464,G13465,G13466,G13467,G13468,G13469,G13470,G13471,G13472,G13473,G13474,G13475,G13476,G13477,G13478,G13479,G13480,
       G13481,G13482,G13483,G13484,G13485,G13486,G13487,G13488,G13489,G13490,G13491,G13492,G13493,G13494,G13495,G13496,G13497,G13498,G13499,G13500,
       G13501,G13502,G13503,G13504,G13505,G13506,G13507,G13508,G13509,G13510,G13511,G13512,G13513,G13514,G13515,G13516,G13517,G13518,G13519,G13520,
       G13521,G13522,G13523,G13524,G13525,G13526,G13527,G13528,G13529,G13530,G13531,G13532,G13533,G13534,G13535,G13536,G13537,G13538,G13539,G13540,
       G13541,G13542,G13543,G13544,G13545,G13546,G13547,G13548,G13549,G13550,G13551,G13552,G13553,G13554,G13555,G13556,G13557,G13558,G13559,G13560,
       G13561,G13562,G13563,G13564,G13565,G13566,G13567,G13568,G13569,G13570,G13571,G13572,G13573,G13574,G13575,G13576,G13577,G13578,G13579,G13580,
       G13581,G13582,G13583,G13584,G13585,G13586,G13587,G13588,G13589,G13590,G13591,G13592,G13593,G13594,G13595,G13596,G13597,G13598,G13599,G13600,
       G13601,G13602,G13603,G13604,G13605,G13606,G13607,G13608,G13609,G13610,G13611,G13612,G13613,G13614,G13615,G13616,G13617,G13618,G13619,G13620,
       G13621,G13622,G13623,G13624,G13625,G13626,G13627,G13628,G13629,G13630,G13631,G13632,G13633,G13634,G13635,G13636,G13637,G13638,G13639,G13640,
       G13641,G13642,G13643,G13644,G13645,G13646,G13647,G13648,G13649,G13650,G13651,G13652,G13653,G13654,G13655,G13656,G13657,G13658,G13659,G13660,
       G13661,G13662,G13663,G13664,G13665,G13666,G13667,G13668,G13669,G13670,G13671,G13672,G13673,G13674,G13675,G13676,G13677,G13678,G13679,G13680,
       G13681,G13682,G13683,G13684,G13685,G13686,G13687,G13688,G13689,G13690,G13691,G13692,G13693,G13694,G13695,G13696,G13697,G13698,G13699,G13700,
       G13701,G13702,G13703,G13704,G13705,G13706,G13707,G13708,G13709,G13710,G13711,G13712,G13713,G13714,G13715,G13716,G13717,G13718,G13719,G13720,
       G13721,G13722,G13723,G13724,G13725,G13726,G13727,G13728,G13729,G13730,G13731,G13732,G13733,G13734,G13735,G13736,G13737,G13738,G13739,G13740,
       G13741,G13742,G13743,G13744,G13745,G13746,G13747,G13748,G13749,G13750,G13751,G13752,G13753,G13754,G13755,G13756,G13757,G13758,G13759,G13760,
       G13761,G13762,G13763,G13764,G13765,G13766,G13767,G13768,G13769,G13770,G13771,G13772,G13773,G13774,G13775,G13776,G13777,G13778,G13779,G13780,
       G13781,G13782,G13783,G13784,G13785,G13786,G13787,G13788,G13789,G13790,G13791,G13792,G13793,G13794,G13795,G13796,G13797,G13798,G13799,G13800,
       G13801,G13802,G13803,G13804,G13805,G13806,G13807,G13808,G13809,G13810,G13811,G13812,G13813,G13814,G13815,G13816,G13817,G13818,G13819,G13820,
       G13821,G13822,G13823,G13824,G13825,G13826,G13827,G13828,G13829,G13830,G13831,G13832,G13833,G13834,G13835,G13836,G13837,G13838,G13839,G13840,
       G13841,G13842,G13843,G13844,G13845,G13846,G13847,G13848,G13849,G13850,G13851,G13852,G13853,G13854,G13855,G13856,G13857,G13858,G13859,G13860,
       G13861,G13862,G13863,G13864,G13865,G13866,G13867,G13868,G13869,G13870,G13871,G13872,G13873,G13874,G13875,G13876,G13877,G13878,G13879,G13880,
       G13881,G13882,G13883,G13884,G13885,G13886,G13887,G13888,G13889,G13890,G13891,G13892,G13893,G13894,G13895,G13896,G13897,G13898,G13899,G13900,
       G13901,G13902,G13903,G13904,G13905,G13906,G13907,G13908,G13909,G13910,G13911,G13912,G13913,G13914,G13915,G13916,G13917,G13918,G13919,G13920,
       G13921,G13922,G13923,G13924,G13925,G13926,G13927,G13928,G13929,G13930,G13931,G13932,G13933,G13934,G13935,G13936,G13937,G13938,G13939,G13940,
       G13941,G13942,G13943,G13944,G13945,G13946,G13947,G13948,G13949,G13950,G13951,G13952,G13953,G13954,G13955,G13956,G13957,G13958,G13959,G13960,
       G13961,G13962,G13963,G13964,G13965,G13966,G13967,G13968,G13969,G13970,G13971,G13972,G13973,G13974,G13975,G13976,G13977,G13978,G13979,G13980,
       G13981,G13982,G13983,G13984,G13985,G13986,G13987,G13988,G13989,G13990,G13991,G13992,G13993,G13994,G13995,G13996,G13997,G13998,G13999,G14000,
       G14001,G14002,G14003,G14004,G14005,G14006,G14007,G14008,G14009,G14010,G14011,G14012,G14013,G14014,G14015,G14016,G14017,G14018,G14019,G14020,
       G14021,G14022,G14023,G14024,G14025,G14026,G14027,G14028,G14029,G14030,G14031,G14032,G14033,G14034,G14035,G14036,G14037,G14038,G14039,G14040,
       G14041,G14042,G14043,G14044,G14045,G14046,G14047,G14048,G14049,G14050,G14051,G14052,G14053,G14054,G14055,G14056,G14057,G14058,G14059,G14060,
       G14061,G14062,G14063,G14064,G14065,G14066,G14067,G14068,G14069,G14070,G14071,G14072,G14073,G14074,G14075,G14076,G14077,G14078,G14079,G14080,
       G14081,G14082,G14083,G14084,G14085,G14086,G14087,G14088,G14089,G14090,G14091,G14092,G14093,G14094,G14095,G14096,G14097,G14098,G14099,G14100,
       G14101,G14102,G14103,G14104,G14105,G14106,G14107,G14108,G14109,G14110,G14111,G14112,G14113,G14114,G14115,G14116,G14117,G14118,G14119,G14120,
       G14121,G14122,G14123,G14124,G14125,G14126,G14127,G14128,G14129,G14130,G14131,G14132,G14133,G14134,G14135,G14136,G14137,G14138,G14139,G14140,
       G14141,G14142,G14143,G14144,G14145,G14146,G14147,G14148,G14149,G14150,G14151,G14152,G14153,G14154,G14155,G14156,G14157,G14158,G14159,G14160,
       G14161,G14162,G14163,G14164,G14165,G14166,G14167,G14168,G14169,G14170,G14171,G14172,G14173,G14174,G14175,G14176,G14177,G14178,G14179,G14180,
       G14181,G14182,G14183,G14184,G14185,G14186,G14187,G14188,G14189,G14190,G14191,G14192,G14193,G14194,G14195,G14196,G14197,G14198,G14199,G14200,
       G14201,G14202,G14203,G14204,G14205,G14206,G14207,G14208,G14209,G14210,G14211,G14212,G14213,G14214,G14215,G14216,G14217,G14218,G14219,G14220,
       G14221,G14222,G14223,G14224,G14225,G14226,G14227,G14228,G14229,G14230,G14231,G14232,G14233,G14234,G14235,G14236,G14237,G14238,G14239,G14240,
       G14241,G14242,G14243,G14244,G14245,G14246,G14247,G14248,G14249,G14250,G14251,G14252,G14253,G14254,G14255,G14256,G14257,G14258,G14259,G14260,
       G14261,G14262,G14263,G14264,G14265,G14266,G14267,G14268,G14269,G14270,G14271,G14272,G14273,G14274,G14275,G14276,G14277,G14278,G14279,G14280,
       G14281,G14282,G14283,G14284,G14285,G14286,G14287,G14288,G14289,G14290,G14291,G14292,G14293,G14294,G14295,G14296,G14297,G14298,G14299,G14300,
       G14301,G14302,G14303,G14304,G14305,G14306,G14307,G14308,G14309,G14310,G14311,G14312,G14313,G14314,G14315,G14316,G14317,G14318,G14319,G14320,
       G14321,G14322,G14323,G14324,G14325,G14326,G14327,G14328,G14329,G14330,G14331,G14332,G14333,G14334,G14335,G14336,G14337,G14338,G14339,G14340,
       G14341,G14342,G14343,G14344,G14345,G14346,G14347,G14348,G14349,G14350,G14351,G14352,G14353,G14354,G14355,G14356,G14357,G14358,G14359,G14360,
       G14361,G14362,G14363,G14364,G14365,G14366,G14367,G14368,G14369,G14370,G14371,G14372,G14373,G14374,G14375,G14376,G14377,G14378,G14379,G14380,
       G14381,G14382,G14383,G14384,G14385,G14386,G14387,G14388,G14389,G14390,G14391,G14392,G14393,G14394,G14395,G14396,G14397,G14398,G14399,G14400,
       G14401,G14402,G14403,G14404,G14405,G14406,G14407,G14408,G14409,G14410,G14411,G14412,G14413,G14414,G14415,G14416,G14417,G14418,G14419,G14420,
       G14421,G14422,G14423,G14424,G14425,G14426,G14427,G14428,G14429,G14430,G14431,G14432,G14433,G14434,G14435,G14436,G14437,G14438,G14439,G14440,
       G14441,G14442,G14443,G14444,G14445,G14446,G14447,G14448,G14449,G14450,G14451,G14452,G14453,G14454,G14455,G14456,G14457,G14458,G14459,G14460,
       G14461,G14462,G14463,G14464,G14465,G14466,G14467,G14468,G14469,G14470,G14471,G14472,G14473,G14474,G14475,G14476,G14477,G14478,G14479,G14480,
       G14481,G14482,G14483,G14484,G14485,G14486,G14487,G14488,G14489,G14490,G14491,G14492,G14493,G14494,G14495,G14496,G14497,G14498,G14499,G14500,
       G14501,G14502,G14503,G14504,G14505,G14506,G14507,G14508,G14509,G14510,G14511,G14512,G14513,G14514,G14515,G14516,G14517,G14518,G14519,G14520,
       G14521,G14522,G14523,G14524,G14525,G14526,G14527,G14528,G14529,G14530,G14531,G14532,G14533,G14534,G14535,G14536,G14537,G14538,G14539,G14540,
       G14541,G14542,G14543,G14544,G14545,G14546,G14547,G14548,G14549,G14550,G14551,G14552,G14553,G14554,G14555,G14556,G14557,G14558,G14559,G14560,
       G14561,G14562,G14563,G14564,G14565,G14566,G14567,G14568,G14569,G14570,G14571,G14572,G14573,G14574,G14575,G14576,G14577,G14578,G14579,G14580,
       G14581,G14582,G14583,G14584,G14585,G14586,G14587,G14588,G14589,G14590,G14591,G14592,G14593,G14594,G14595,G14596,G14597,G14598,G14599,G14600,
       G14601,G14602,G14603,G14604,G14605,G14606,G14607,G14608,G14609,G14610,G14611,G14612,G14613,G14614,G14615,G14616,G14617,G14618,G14619,G14620,
       G14621,G14622,G14623,G14624,G14625,G14626,G14627,G14628,G14629,G14630,G14631,G14632,G14633,G14634,G14635,G14636,G14637,G14638,G14639,G14640,
       G14641,G14642,G14643,G14644,G14645,G14646,G14647,G14648,G14649,G14650,G14651,G14652,G14653,G14654,G14655,G14656,G14657,G14658,G14659,G14660,
       G14661,G14662,G14663,G14664,G14665,G14666,G14667,G14668,G14669,G14670,G14671,G14672,G14673,G14674,G14675,G14676,G14677,G14678,G14679,G14680,
       G14681,G14682,G14683,G14684,G14685,G14686,G14687,G14688,G14689,G14690,G14691,G14692,G14693,G14694,G14695,G14696,G14697,G14698,G14699,G14700,
       G14701,G14702,G14703,G14704,G14705,G14706,G14707,G14708,G14709,G14710,G14711,G14712,G14713,G14714,G14715,G14716,G14717,G14718,G14719,G14720,
       G14721,G14722,G14723,G14724,G14725,G14726,G14727,G14728,G14729,G14730,G14731,G14732,G14733,G14734,G14735,G14736,G14737,G14738,G14739,G14740,
       G14741,G14742,G14743,G14744,G14745,G14746,G14747,G14748,G14749,G14750,G14751,G14752,G14753,G14754,G14755,G14756,G14757,G14758,G14759,G14760,
       G14761,G14762,G14763,G14764,G14765,G14766,G14767,G14768,G14769,G14770,G14771,G14772,G14773,G14774,G14775,G14776,G14777,G14778,G14779,G14780,
       G14781,G14782,G14783,G14784,G14785,G14786,G14787,G14788,G14789,G14790,G14791,G14792,G14793,G14794,G14795,G14796,G14797,G14798,G14799,G14800,
       G14801,G14802,G14803,G14804,G14805,G14806,G14807,G14808,G14809,G14810,G14811,G14812,G14813,G14814,G14815,G14816,G14817,G14818,G14819,G14820,
       G14821,G14822,G14823,G14824,G14825,G14826,G14827,G14828,G14829,G14830,G14831,G14832,G14833,G14834,G14835,G14836,G14837,G14838,G14839,G14840,
       G14841,G14842,G14843,G14844,G14845,G14846,G14847,G14848,G14849,G14850,G14851,G14852,G14853,G14854,G14855,G14856,G14857,G14858,G14859,G14860,
       G14861,G14862,G14863,G14864,G14865,G14866,G14867,G14868,G14869,G14870,G14871,G14872,G14873,G14874,G14875,G14876,G14877,G14878,G14879,G14880,
       G14881,G14882,G14883,G14884,G14885,G14886,G14887,G14888,G14889,G14890,G14891,G14892,G14893,G14894,G14895,G14896,G14897,G14898,G14899,G14900,
       G14901,G14902,G14903,G14904,G14905,G14906,G14907,G14908,G14909,G14910,G14911,G14912,G14913,G14914,G14915,G14916,G14917,G14918,G14919,G14920,
       G14921,G14922,G14923,G14924,G14925,G14926,G14927,G14928,G14929,G14930,G14931,G14932,G14933,G14934,G14935,G14936,G14937,G14938,G14939,G14940,
       G14941,G14942,G14943,G14944,G14945,G14946,G14947,G14948,G14949,G14950,G14951,G14952,G14953,G14954,G14955,G14956,G14957,G14958,G14959,G14960,
       G14961,G14962,G14963,G14964,G14965,G14966,G14967,G14968,G14969,G14970,G14971,G14972,G14973,G14974,G14975,G14976,G14977,G14978,G14979,G14980,
       G14981,G14982,G14983,G14984,G14985,G14986,G14987,G14988,G14989,G14990,G14991,G14992,G14993,G14994,G14995,G14996,G14997,G14998,G14999,G15000,
       G15001,G15002,G15003,G15004,G15005,G15006,G15007,G15008,G15009,G15010,G15011,G15012,G15013,G15014,G15015,G15016,G15017,G15018,G15019,G15020,
       G15021,G15022,G15023,G15024,G15025,G15026,G15027,G15028,G15029,G15030,G15031,G15032,G15033,G15034,G15035,G15036,G15037,G15038,G15039,G15040,
       G15041,G15042,G15043,G15044,G15045,G15046,G15047,G15048,G15049,G15050,G15051,G15052,G15053,G15054,G15055,G15056,G15057,G15058,G15059,G15060,
       G15061,G15062,G15063,G15064,G15065,G15066,G15067,G15068,G15069,G15070,G15071,G15072,G15073,G15074,G15075,G15076,G15077,G15078,G15079,G15080,
       G15081,G15082,G15083,G15084,G15085,G15086,G15087,G15088,G15089,G15090,G15091,G15092,G15093,G15094,G15095,G15096,G15097,G15098,G15099,G15100,
       G15101,G15102,G15103,G15104,G15105,G15106,G15107,G15108,G15109,G15110,G15111,G15112,G15113,G15114,G15115,G15116,G15117,G15118,G15119,G15120,
       G15121,G15122,G15123,G15124,G15125,G15126,G15127,G15128,G15129,G15130,G15131,G15132,G15133,G15134,G15135,G15136,G15137,G15138,G15139,G15140,
       G15141,G15142,G15143,G15144,G15145,G15146,G15147,G15148,G15149,G15150,G15151,G15152,G15153,G15154,G15155,G15156,G15157,G15158,G15159,G15160,
       G15161,G15162,G15163,G15164,G15165,G15166,G15167,G15168,G15169,G15170,G15171,G15172,G15173,G15174,G15175,G15176,G15177,G15178,G15179,G15180,
       G15181,G15182,G15183,G15184,G15185,G15186,G15187,G15188,G15189,G15190,G15191,G15192,G15193,G15194,G15195,G15196,G15197,G15198,G15199,G15200,
       G15201,G15202,G15203,G15204,G15205,G15206,G15207,G15208,G15209,G15210,G15211,G15212,G15213,G15214,G15215,G15216,G15217,G15218,G15219,G15220,
       G15221,G15222,G15223,G15224,G15225,G15226,G15227,G15228,G15229,G15230,G15231,G15232,G15233,G15234,G15235,G15236,G15237,G15238,G15239,G15240,
       G15241,G15242,G15243,G15244,G15245,G15246,G15247,G15248,G15249,G15250,G15251,G15252,G15253,G15254,G15255,G15256,G15257,G15258,G15259,G15260,
       G15261,G15262,G15263,G15264,G15265,G15266,G15267,G15268,G15269,G15270,G15271,G15272,G15273,G15274,G15275,G15276,G15277,G15278,G15279,G15280,
       G15281,G15282,G15283,G15284,G15285,G15286,G15287,G15288,G15289,G15290,G15291,G15292,G15293,G15294,G15295,G15296,G15297,G15298,G15299,G15300,
       G15301,G15302,G15303,G15304,G15305,G15306,G15307,G15308,G15309,G15310,G15311,G15312,G15313,G15314,G15315,G15316,G15317,G15318,G15319,G15320,
       G15321,G15322,G15323,G15324,G15325,G15326,G15327,G15328,G15329,G15330,G15331,G15332,G15333,G15334,G15335,G15336,G15337,G15338,G15339,G15340,
       G15341,G15342,G15343,G15344,G15345,G15346,G15347,G15348,G15349,G15350,G15351,G15352,G15353,G15354,G15355,G15356,G15357,G15358,G15359,G15360,
       G15361,G15362,G15363,G15364,G15365,G15366,G15367,G15368,G15369,G15370,G15371,G15372,G15373,G15374,G15375,G15376,G15377,G15378,G15379,G15380,
       G15381,G15382,G15383,G15384,G15385,G15386,G15387,G15388,G15389,G15390,G15391,G15392,G15393,G15394,G15395,G15396,G15397,G15398,G15399,G15400,
       G15401,G15402,G15403,G15404,G15405,G15406,G15407,G15408,G15409,G15410,G15411,G15412,G15413,G15414,G15415,G15416,G15417,G15418,G15419,G15420,
       G15421,G15422,G15423,G15424,G15425,G15426,G15427,G15428,G15429,G15430,G15431,G15432,G15433,G15434,G15435,G15436,G15437,G15438,G15439,G15440,
       G15441,G15442,G15443,G15444,G15445,G15446,G15447,G15448,G15449,G15450,G15451,G15452,G15453,G15454,G15455,G15456,G15457,G15458,G15459,G15460,
       G15461,G15462,G15463,G15464,G15465,G15466,G15467,G15468,G15469,G15470,G15471,G15472,G15473,G15474,G15475,G15476,G15477,G15478,G15479,G15480,
       G15481,G15482,G15483,G15484,G15485,G15486,G15487,G15488,G15489,G15490,G15491,G15492,G15493,G15494,G15495,G15496,G15497,G15498,G15499,G15500,
       G15501,G15502,G15503,G15504,G15505,G15506,G15507,G15508,G15509,G15510,G15511,G15512,G15513,G15514,G15515,G15516,G15517,G15518,G15519,G15520,
       G15521,G15522,G15523,G15524,G15525,G15526,G15527,G15528,G15529,G15530,G15531,G15532,G15533,G15534,G15535,G15536,G15537,G15538,G15539,G15540,
       G15541,G15542,G15543,G15544,G15545,G15546,G15547,G15548,G15549,G15550,G15551,G15552,G15553,G15554,G15555,G15556,G15557,G15558,G15559,G15560,
       G15561,G15562,G15563,G15564,G15565,G15566,G15567,G15568,G15569,G15570,G15571,G15572,G15573,G15574,G15575,G15576,G15577,G15578,G15579,G15580,
       G15581,G15582,G15583,G15584,G15585,G15586,G15587,G15588,G15589,G15590,G15591,G15592,G15593,G15594,G15595,G15596,G15597,G15598,G15599,G15600,
       G15601,G15602,G15603,G15604,G15605,G15606,G15607,G15608,G15609,G15610,G15611,G15612,G15613,G15614,G15615,G15616,G15617,G15618,G15619,G15620,
       G15621,G15622,G15623,G15624,G15625,G15626,G15627,G15628,G15629,G15630,G15631,G15632,G15633,G15634,G15635,G15636,G15637,G15638,G15639,G15640,
       G15641,G15642,G15643,G15644,G15645,G15646,G15647,G15648,G15649,G15650,G15651,G15652,G15653,G15654,G15655,G15656,G15657,G15658,G15659,G15660,
       G15661,G15662,G15663,G15664,G15665,G15666,G15667,G15668,G15669,G15670,G15671,G15672,G15673,G15674,G15675,G15676,G15677,G15678,G15679,G15680,
       G15681,G15682,G15683,G15684,G15685,G15686,G15687,G15688,G15689,G15690,G15691,G15692,G15693,G15694,G15695,G15696,G15697,G15698,G15699,G15700,
       G15701,G15702,G15703,G15704,G15705,G15706,G15707,G15708,G15709,G15710,G15711,G15712,G15713,G15714,G15715,G15716,G15717,G15718,G15719,G15720,
       G15721,G15722,G15723,G15724,G15725,G15726,G15727,G15728,G15729,G15730,G15731,G15732,G15733,G15734,G15735,G15736,G15737,G15738,G15739,G15740,
       G15741,G15742,G15743,G15744,G15745,G15746,G15747,G15748,G15749,G15750,G15751,G15752,G15753,G15754,G15755,G15756,G15757,G15758,G15759,G15760,
       G15761,G15762,G15763,G15764,G15765,G15766,G15767,G15768,G15769,G15770,G15771,G15772,G15773,G15774,G15775,G15776,G15777,G15778,G15779,G15780,
       G15781,G15782,G15783,G15784,G15785,G15786,G15787,G15788,G15789,G15790,G15791,G15792,G15793,G15794,G15795,G15796,G15797,G15798,G15799,G15800,
       G15801,G15802,G15803,G15804,G15805,G15806,G15807,G15808,G15809,G15810,G15811,G15812,G15813,G15814,G15815,G15816,G15817,G15818,G15819,G15820,
       G15821,G15822,G15823,G15824,G15825,G15826,G15827,G15828,G15829,G15830,G15831,G15832,G15833,G15834,G15835,G15836,G15837,G15838,G15839,G15840,
       G15841,G15842,G15843,G15844,G15845,G15846,G15847,G15848,G15849,G15850,G15851,G15852,G15853,G15854,G15855,G15856,G15857,G15858,G15859,G15860,
       G15861,G15862,G15863,G15864,G15865,G15866,G15867,G15868,G15869,G15870,G15871,G15872,G15873,G15874,G15875,G15876,G15877,G15878,G15879,G15880,
       G15881,G15882,G15883,G15884,G15885,G15886,G15887,G15888,G15889,G15890,G15891,G15892,G15893,G15894,G15895,G15896,G15897,G15898,G15899,G15900,
       G15901,G15902,G15903,G15904,G15905,G15906,G15907,G15908,G15909,G15910,G15911,G15912,G15913,G15914,G15915,G15916,G15917,G15918,G15919,G15920,
       G15921,G15922,G15923,G15924,G15925,G15926,G15927,G15928,G15929,G15930,G15931,G15932,G15933,G15934,G15935,G15936,G15937,G15938,G15939,G15940,
       G15941,G15942,G15943,G15944,G15945,G15946,G15947,G15948,G15949,G15950,G15951,G15952,G15953,G15954,G15955,G15956,G15957,G15958,G15959,G15960,
       G15961,G15962,G15963,G15964,G15965,G15966,G15967,G15968,G15969,G15970,G15971,G15972,G15973,G15974,G15975,G15976,G15977,G15978,G15979,G15980,
       G15981,G15982,G15983,G15984,G15985,G15986,G15987,G15988,G15989,G15990,G15991,G15992,G15993,G15994,G15995,G15996,G15997,G15998,G15999,G16000,
       G16001,G16002,G16003,G16004,G16005,G16006,G16007,G16008,G16009,G16010,G16011,G16012,G16013,G16014,G16015,G16016,G16017,G16018,G16019,G16020,
       G16021,G16022,G16023,G16024,G16025,G16026,G16027,G16028,G16029,G16030,G16031,G16032,G16033,G16034,G16035,G16036,G16037,G16038,G16039,G16040,
       G16041,G16042,G16043,G16044,G16045,G16046,G16047,G16048,G16049,G16050,G16051,G16052,G16053,G16054,G16055,G16056,G16057,G16058,G16059,G16060,
       G16061,G16062,G16063,G16064,G16065,G16066,G16067,G16068,G16069,G16070,G16071,G16072,G16073,G16074,G16075,G16076,G16077,G16078,G16079,G16080,
       G16081,G16082,G16083,G16084,G16085,G16086,G16087,G16088,G16089,G16090,G16091,G16092,G16093,G16094,G16095,G16096,G16097,G16098,G16099,G16100,
       G16101,G16102,G16103,G16104,G16105,G16106,G16107,G16108,G16109,G16110,G16111,G16112,G16113,G16114,G16115,G16116,G16117,G16118,G16119,G16120,
       G16121,G16122,G16123,G16124,G16125,G16126,G16127,G16128,G16129,G16130,G16131,G16132,G16133,G16134,G16135,G16136,G16137,G16138,G16139,G16140,
       G16141,G16142,G16143,G16144,G16145,G16146,G16147,G16148,G16149,G16150,G16151,G16152,G16153,G16154,G16155,G16156,G16157,G16158,G16159,G16160,
       G16161,G16162,G16163,G16164,G16165,G16166,G16167,G16168,G16169,G16170,G16171,G16172,G16173,G16174,G16175,G16176,G16177,G16178,G16179,G16180,
       G16181,G16182,G16183,G16184,G16185,G16186,G16187,G16188,G16189,G16190,G16191,G16192,G16193,G16194,G16195,G16196,G16197,G16198,G16199,G16200,
       G16201,G16202,G16203,G16204,G16205,G16206,G16207,G16208,G16209,G16210,G16211,G16212,G16213,G16214,G16215,G16216,G16217,G16218,G16219,G16220,
       G16221,G16222,G16223,G16224,G16225,G16226,G16227,G16228,G16229,G16230,G16231,G16232,G16233,G16234,G16235,G16236,G16237,G16238,G16239,G16240,
       G16241,G16242,G16243,G16244,G16245,G16246,G16247,G16248,G16249,G16250,G16251,G16252,G16253,G16254,G16255,G16256,G16257,G16258,G16259,G16260,
       G16261,G16262,G16263,G16264,G16265,G16266,G16267,G16268,G16269,G16270,G16271,G16272,G16273,G16274,G16275,G16276,G16277,G16278,G16279,G16280,
       G16281,G16282,G16283,G16284,G16285,G16286,G16287,G16288,G16289,G16290,G16291,G16292,G16293,G16294,G16295,G16296,G16297,G16298,G16299,G16300,
       G16301,G16302,G16303,G16304,G16305,G16306,G16307,G16308,G16309,G16310,G16311,G16312,G16313,G16314,G16315,G16316,G16317,G16318,G16319,G16320,
       G16321,G16322,G16323,G16324,G16325,G16326,G16327,G16328,G16329,G16330,G16331,G16332,G16333,G16334,G16335,G16336,G16337,G16338,G16339,G16340,
       G16341,G16342,G16343,G16344,G16345,G16346,G16347,G16348,G16349,G16350,G16351,G16352,G16353,G16354,G16355,G16356,G16357,G16358,G16359,G16360,
       G16361,G16362,G16363,G16364,G16365,G16366,G16367,G16368,G16369,G16370,G16371,G16372,G16373,G16374,G16375,G16376,G16377,G16378,G16379,G16380,
       G16381,G16382,G16383,G16384,G16385,G16386,G16387,G16388,G16389,G16390,G16391,G16392,G16393,G16394,G16395,G16396,G16397,G16398,G16399,G16400,
       G16401,G16402,G16403,G16404,G16405,G16406,G16407,G16408,G16409,G16410,G16411,G16412,G16413,G16414,G16415,G16416,G16417,G16418,G16419,G16420,
       G16421,G16422,G16423,G16424,G16425,G16426,G16427,G16428,G16429,G16430,G16431,G16432,G16433,G16434,G16435,G16436,G16437,G16438,G16439,G16440,
       G16441,G16442,G16443,G16444,G16445,G16446,G16447,G16448,G16449,G16450,G16451,G16452,G16453,G16454,G16455,G16456,G16457,G16458,G16459,G16460,
       G16461,G16462,G16463,G16464,G16465,G16466,G16467,G16468,G16469,G16470,G16471,G16472,G16473,G16474,G16475,G16476,G16477,G16478,G16479,G16480,
       G16481,G16482,G16483,G16484,G16485,G16486,G16487,G16488,G16489,G16490,G16491,G16492,G16493,G16494,G16495,G16496,G16497,G16498,G16499,G16500,
       G16501,G16502,G16503,G16504,G16505,G16506,G16507,G16508,G16509,G16510,G16511,G16512,G16513,G16514,G16515,G16516,G16517,G16518,G16519,G16520,
       G16521,G16522,G16523,G16524,G16525,G16526,G16527,G16528,G16529,G16530,G16531,G16532,G16533,G16534,G16535,G16536,G16537,G16538,G16539,G16540,
       G16541,G16542,G16543,G16544,G16545,G16546,G16547,G16548,G16549,G16550,G16551,G16552,G16553,G16554,G16555,G16556,G16557,G16558,G16559,G16560,
       G16561,G16562,G16563,G16564,G16565,G16566,G16567,G16568,G16569,G16570,G16571,G16572,G16573,G16574,G16575,G16576,G16577,G16578,G16579,G16580,
       G16581,G16582,G16583,G16584,G16585,G16586,G16587,G16588,G16589,G16590,G16591,G16592,G16593,G16594,G16595,G16596,G16597,G16598,G16599,G16600,
       G16601,G16602,G16603,G16604,G16605,G16606,G16607,G16608,G16609,G16610,G16611,G16612,G16613,G16614,G16615,G16616,G16617,G16618,G16619,G16620,
       G16621,G16622,G16623,G16624,G16625,G16626,G16627,G16628,G16629,G16630,G16631,G16632,G16633,G16634,G16635,G16636,G16637,G16638,G16639,G16640,
       G16641,G16642,G16643,G16644,G16645,G16646,G16647,G16648,G16649,G16650,G16651,G16652,G16653,G16654,G16655,G16656,G16657,G16658,G16659,G16660,
       G16661,G16662,G16663,G16664,G16665,G16666,G16667,G16668,G16669,G16670,G16671,G16672,G16673,G16674,G16675,G16676,G16677,G16678,G16679,G16680,
       G16681,G16682,G16683,G16684,G16685,G16686,G16687,G16688,G16689,G16690,G16691,G16692,G16693,G16694,G16695,G16696,G16697,G16698,G16699,G16700,
       G16701,G16702,G16703,G16704,G16705,G16706,G16707,G16708,G16709,G16710,G16711,G16712,G16713,G16714,G16715,G16716,G16717,G16718,G16719,G16720,
       G16721,G16722,G16723,G16724,G16725,G16726,G16727,G16728,G16729,G16730,G16731,G16732,G16733,G16734,G16735,G16736,G16737,G16738,G16739,G16740,
       G16741,G16742,G16743,G16744,G16745,G16746,G16747,G16748,G16749,G16750,G16751,G16752,G16753,G16754,G16755,G16756,G16757,G16758,G16759,G16760,
       G16761,G16762,G16763,G16764,G16765,G16766,G16767,G16768,G16769,G16770,G16771,G16772,G16773,G16774,G16775,G16776,G16777,G16778,G16779,G16780,
       G16781,G16782,G16783,G16784,G16785,G16786,G16787,G16788,G16789,G16790,G16791,G16792,G16793,G16794,G16795,G16796,G16797,G16798,G16799,G16800,
       G16801,G16802,G16803,G16804,G16805,G16806,G16807,G16808,G16809,G16810,G16811,G16812,G16813,G16814,G16815,G16816,G16817,G16818,G16819,G16820,
       G16821,G16822,G16823,G16824,G16825,G16826,G16827,G16828,G16829,G16830,G16831,G16832,G16833,G16834,G16835,G16836,G16837,G16838,G16839,G16840,
       G16841,G16842,G16843,G16844,G16845,G16846,G16847,G16848,G16849,G16850,G16851,G16852,G16853,G16854,G16855,G16856,G16857,G16858,G16859,G16860,
       G16861,G16862,G16863,G16864,G16865,G16866,G16867,G16868,G16869,G16870,G16871,G16872,G16873,G16874,G16875,G16876,G16877,G16878,G16879,G16880,
       G16881,G16882,G16883,G16884,G16885,G16886,G16887,G16888,G16889,G16890,G16891,G16892,G16893,G16894,G16895,G16896,G16897,G16898,G16899,G16900,
       G16901,G16902,G16903,G16904,G16905,G16906,G16907,G16908,G16909,G16910,G16911,G16912,G16913,G16914,G16915,G16916,G16917,G16918,G16919,G16920,
       G16921,G16922,G16923,G16924,G16925,G16926,G16927,G16928,G16929,G16930,G16931,G16932,G16933,G16934,G16935,G16936,G16937,G16938,G16939,G16940,
       G16941,G16942,G16943,G16944,G16945,G16946,G16947,G16948,G16949,G16950,G16951,G16952,G16953,G16954,G16955,G16956,G16957,G16958,G16959,G16960,
       G16961,G16962,G16963,G16964,G16965,G16966,G16967,G16968,G16969,G16970,G16971,G16972,G16973,G16974,G16975,G16976,G16977,G16978,G16979,G16980,
       G16981,G16982,G16983,G16984,G16985,G16986,G16987,G16988,G16989,G16990,G16991,G16992,G16993,G16994,G16995,G16996,G16997,G16998,G16999,G17000,
       G17001,G17002,G17003,G17004,G17005,G17006,G17007,G17008,G17009,G17010,G17011,G17012,G17013,G17014,G17015,G17016,G17017,G17018,G17019,G17020,
       G17021,G17022,G17023,G17024,G17025,G17026,G17027,G17028,G17029,G17030,G17031,G17032,G17033,G17034,G17035,G17036,G17037,G17038,G17039,G17040,
       G17041,G17042,G17043,G17044,G17045,G17046,G17047,G17048,G17049,G17050,G17051,G17052,G17053,G17054,G17055,G17056,G17057,G17058,G17059,G17060,
       G17061,G17062,G17063,G17064,G17065,G17066,G17067,G17068,G17069,G17070,G17071,G17072,G17073,G17074,G17075,G17076,G17077,G17078,G17079,G17080,
       G17081,G17082,G17083,G17084,G17085,G17086,G17087,G17088,G17089,G17090,G17091,G17092,G17093,G17094,G17095,G17096,G17097,G17098,G17099,G17100,
       G17101,G17102,G17103,G17104,G17105,G17106,G17107,G17108,G17109,G17110,G17111,G17112,G17113,G17114,G17115,G17116,G17117,G17118,G17119,G17120,
       G17121,G17122,G17123,G17124,G17125,G17126,G17127,G17128,G17129,G17130,G17131,G17132,G17133,G17134,G17135,G17136,G17137,G17138,G17139,G17140,
       G17141,G17142,G17143,G17144,G17145,G17146,G17147,G17148,G17149,G17150,G17151,G17152,G17153,G17154,G17155,G17156,G17157,G17158,G17159,G17160,
       G17161,G17162,G17163,G17164,G17165,G17166,G17167,G17168,G17169,G17170,G17171,G17172,G17173,G17174,G17175,G17176,G17177,G17178,G17179,G17180,
       G17181,G17182,G17183,G17184,G17185,G17186,G17187,G17188,G17189,G17190,G17191,G17192,G17193,G17194,G17195,G17196,G17197,G17198,G17199,G17200,
       G17201,G17202,G17203,G17204,G17205,G17206,G17207,G17208,G17209,G17210,G17211,G17212,G17213,G17214,G17215,G17216,G17217,G17218,G17219,G17220,
       G17221,G17222,G17223,G17224,G17225,G17226,G17227,G17228,G17229,G17230,G17231,G17232,G17233,G17234,G17235,G17236,G17237,G17238,G17239,G17240,
       G17241,G17242,G17243,G17244,G17245,G17246,G17247,G17248,G17249,G17250,G17251,G17252,G17253,G17254,G17255,G17256,G17257,G17258,G17259,G17260,
       G17261,G17262,G17263,G17264,G17265,G17266,G17267,G17268,G17269,G17270,G17271,G17272,G17273,G17274,G17275,G17276,G17277,G17278,G17279,G17280,
       G17281,G17282,G17283,G17284,G17285,G17286,G17287,G17288,G17289,G17290,G17291,G17292,G17293,G17294,G17295,G17296,G17297,G17298,G17299,G17300,
       G17301,G17302,G17303,G17304,G17305,G17306,G17307,G17308,G17309,G17310,G17311,G17312,G17313,G17314,G17315,G17316,G17317,G17318,G17319,G17320,
       G17321,G17322,G17323,G17324,G17325,G17326,G17327,G17328,G17329,G17330,G17331,G17332,G17333,G17334,G17335,G17336,G17337,G17338,G17339,G17340,
       G17341,G17342,G17343,G17344,G17345,G17346,G17347,G17348,G17349,G17350,G17351,G17352,G17353,G17354,G17355,G17356,G17357,G17358,G17359,G17360,
       G17361,G17362,G17363,G17364,G17365,G17366,G17367,G17368,G17369,G17370,G17371,G17372,G17373,G17374,G17375,G17376,G17377,G17378,G17379,G17380,
       G17381,G17382,G17383,G17384,G17385,G17386,G17387,G17388,G17389,G17390,G17391,G17392,G17393,G17394,G17395,G17396,G17397,G17398,G17399,G17400,
       G17401,G17402,G17403,G17404,G17405,G17406,G17407,G17408,G17409,G17410,G17411,G17412,G17413,G17414,G17415,G17416,G17417,G17418,G17419,G17420,
       G17421,G17422,G17423,G17424,G17425,G17426,G17427,G17428,G17429,G17430,G17431,G17432,G17433,G17434,G17435,G17436,G17437,G17438,G17439,G17440,
       G17441,G17442,G17443,G17444,G17445,G17446,G17447,G17448,G17449,G17450,G17451,G17452,G17453,G17454,G17455,G17456,G17457,G17458,G17459,G17460,
       G17461,G17462,G17463,G17464,G17465,G17466,G17467,G17468,G17469,G17470,G17471,G17472,G17473,G17474,G17475,G17476,G17477,G17478,G17479,G17480,
       G17481,G17482,G17483,G17484,G17485,G17486,G17487,G17488,G17489,G17490,G17491,G17492,G17493,G17494,G17495,G17496,G17497,G17498,G17499,G17500,
       G17501,G17502,G17503,G17504,G17505,G17506,G17507,G17508,G17509,G17510,G17511,G17512,G17513,G17514,G17515,G17516,G17517,G17518,G17519,G17520,
       G17521,G17522,G17523,G17524,G17525,G17526,G17527,G17528,G17529,G17530,G17531,G17532,G17533,G17534,G17535,G17536,G17537,G17538,G17539,G17540,
       G17541,G17542,G17543,G17544,G17545,G17546,G17547,G17548,G17549,G17550,G17551,G17552,G17553,G17554,G17555,G17556,G17557,G17558,G17559,G17560,
       G17561,G17562,G17563,G17564,G17565,G17566,G17567,G17568,G17569,G17570,G17571,G17572,G17573,G17574,G17575,G17576,G17577,G17578,G17579,G17580,
       G17581,G17582,G17583,G17584,G17585,G17586,G17587,G17588,G17589,G17590,G17591,G17592,G17593,G17594,G17595,G17596,G17597,G17598,G17599,G17600,
       G17601,G17602,G17603,G17604,G17605,G17606,G17607,G17608,G17609,G17610,G17611,G17612,G17613,G17614,G17615,G17616,G17617,G17618,G17619,G17620,
       G17621,G17622,G17623,G17624,G17625,G17626,G17627,G17628,G17629,G17630,G17631,G17632,G17633,G17634,G17635,G17636,G17637,G17638,G17639,G17640,
       G17641,G17642,G17643,G17644,G17645,G17646,G17647,G17648,G17649,G17650,G17651,G17652,G17653,G17654,G17655,G17656,G17657,G17658,G17659,G17660,
       G17661,G17662,G17663,G17664,G17665,G17666,G17667,G17668,G17669,G17670,G17671,G17672,G17673,G17674,G17675,G17676,G17677,G17678,G17679,G17680,
       G17681,G17682,G17683,G17684,G17685,G17686,G17687,G17688,G17689,G17690,G17691,G17692,G17693,G17694,G17695,G17696,G17697,G17698,G17699,G17700,
       G17701,G17702,G17703,G17704,G17705,G17706,G17707,G17708,G17709,G17710,G17711,G17712,G17713,G17714,G17715,G17716,G17717,G17718,G17719,G17720,
       G17721,G17722,G17723,G17724,G17725,G17726,G17727,G17728,G17729,G17730,G17731,G17732,G17733,G17734,G17735,G17736,G17737,G17738,G17739,G17740,
       G17741,G17742,G17743,G17744,G17745,G17746,G17747,G17748,G17749,G17750,G17751,G17752,G17753,G17754,G17755,G17756,G17757,G17758,G17759,G17760,
       G17761,G17762,G17763,G17764,G17765,G17766,G17767,G17768,G17769,G17770,G17771,G17772,G17773,G17774,G17775,G17776,G17777,G17778,G17779,G17780,
       G17781,G17782,G17783,G17784,G17785,G17786,G17787,G17788,G17789,G17790,G17791,G17792,G17793,G17794,G17795,G17796,G17797,G17798,G17799,G17800,
       G17801,G17802,G17803,G17804,G17805,G17806,G17807,G17808,G17809,G17810,G17811,G17812,G17813,G17814,G17815,G17816,G17817,G17818,G17819,G17820,
       G17821,G17822,G17823,G17824,G17825,G17826,G17827,G17828,G17829,G17830,G17831,G17832,G17833,G17834,G17835,G17836,G17837,G17838,G17839,G17840,
       G17841,G17842,G17843,G17844,G17845,G17846,G17847,G17848,G17849,G17850,G17851,G17852,G17853,G17854,G17855,G17856,G17857,G17858,G17859,G17860,
       G17861,G17862,G17863,G17864,G17865,G17866,G17867,G17868,G17869,G17870,G17871,G17872,G17873,G17874,G17875,G17876,G17877,G17878,G17879,G17880,
       G17881,G17882,G17883,G17884,G17885,G17886,G17887,G17888,G17889,G17890,G17891,G17892,G17893,G17894,G17895,G17896,G17897,G17898,G17899,G17900,
       G17901,G17902,G17903,G17904,G17905,G17906,G17907,G17908,G17909,G17910,G17911,G17912,G17913,G17914,G17915,G17916,G17917,G17918,G17919,G17920,
       G17921,G17922,G17923,G17924,G17925,G17926,G17927,G17928,G17929,G17930,G17931,G17932,G17933,G17934,G17935,G17936,G17937,G17938,G17939,G17940,
       G17941,G17942,G17943,G17944,G17945,G17946,G17947,G17948,G17949,G17950,G17951,G17952,G17953,G17954,G17955,G17956,G17957,G17958,G17959,G17960,
       G17961,G17962,G17963,G17964,G17965,G17966,G17967,G17968,G17969,G17970,G17971,G17972,G17973,G17974,G17975,G17976,G17977,G17978,G17979,G17980,
       G17981,G17982,G17983,G17984,G17985,G17986,G17987,G17988,G17989,G17990,G17991,G17992,G17993,G17994,G17995,G17996,G17997,G17998,G17999,G18000,
       G18001,G18002,G18003,G18004,G18005,G18006,G18007,G18008,G18009,G18010,G18011,G18012,G18013,G18014,G18015,G18016,G18017,G18018,G18019,G18020,
       G18021,G18022,G18023,G18024,G18025,G18026,G18027,G18028,G18029,G18030,G18031,G18032,G18033,G18034,G18035,G18036,G18037,G18038,G18039,G18040,
       G18041,G18042,G18043,G18044,G18045,G18046,G18047,G18048,G18049,G18050,G18051,G18052,G18053,G18054,G18055,G18056,G18057,G18058,G18059,G18060,
       G18061,G18062,G18063,G18064,G18065,G18066,G18067,G18068,G18069,G18070,G18071,G18072,G18073,G18074,G18075,G18076,G18077,G18078,G18079,G18080,
       G18081,G18082,G18083,G18084,G18085,G18086,G18087,G18088,G18089,G18090,G18091,G18092,G18093,G18094,G18095,G18096,G18097,G18098,G18099,G18100,
       G18101,G18102,G18103,G18104,G18105,G18106,G18107,G18108,G18109,G18110,G18111,G18112,G18113,G18114,G18115,G18116,G18117,G18118,G18119,G18120,
       G18121,G18122,G18123,G18124,G18125,G18126,G18127,G18128,G18129,G18130,G18131,G18132,G18133,G18134,G18135,G18136,G18137,G18138,G18139,G18140,
       G18141,G18142,G18143,G18144,G18145,G18146,G18147,G18148,G18149,G18150,G18151,G18152,G18153,G18154,G18155,G18156,G18157,G18158,G18159,G18160,
       G18161,G18162,G18163,G18164,G18165,G18166,G18167,G18168,G18169,G18170,G18171,G18172,G18173,G18174,G18175,G18176,G18177,G18178,G18179,G18180,
       G18181,G18182,G18183,G18184,G18185,G18186,G18187,G18188,G18189,G18190,G18191,G18192,G18193,G18194,G18195,G18196,G18197,G18198,G18199,G18200,
       G18201,G18202,G18203,G18204,G18205,G18206,G18207,G18208,G18209,G18210,G18211,G18212,G18213,G18214,G18215,G18216,G18217,G18218,G18219,G18220,
       G18221,G18222,G18223,G18224,G18225,G18226,G18227,G18228,G18229,G18230,G18231,G18232,G18233,G18234,G18235,G18236,G18237,G18238,G18239,G18240,
       G18241,G18242,G18243,G18244,G18245,G18246,G18247,G18248,G18249,G18250,G18251,G18252,G18253,G18254,G18255,G18256,G18257,G18258,G18259,G18260,
       G18261,G18262,G18263,G18264,G18265,G18266,G18267,G18268,G18269,G18270,G18271,G18272,G18273,G18274,G18275,G18276,G18277,G18278,G18279,G18280,
       G18281,G18282,G18283,G18284,G18285,G18286,G18287,G18288,G18289,G18290,G18291,G18292,G18293,G18294,G18295,G18296,G18297,G18298,G18299,G18300,
       G18301,G18302,G18303,G18304,G18305,G18306,G18307,G18308,G18309,G18310,G18311,G18312,G18313,G18314,G18315,G18316,G18317,G18318,G18319,G18320,
       G18321,G18322,G18323,G18324,G18325,G18326,G18327,G18328,G18329,G18330,G18331,G18332,G18333,G18334,G18335,G18336,G18337,G18338,G18339,G18340,
       G18341,G18342,G18343,G18344,G18345,G18346,G18347,G18348,G18349,G18350,G18351,G18352,G18353,G18354,G18355,G18356,G18357,G18358,G18359,G18360,
       G18361,G18362,G18363,G18364,G18365,G18366,G18367,G18368,G18369,G18370,G18371,G18372,G18373,G18374,G18375,G18376,G18377,G18378,G18379,G18380,
       G18381,G18382,G18383,G18384,G18385,G18386,G18387,G18388,G18389,G18390,G18391,G18392,G18393,G18394,G18395,G18396,G18397,G18398,G18399,G18400,
       G18401,G18402,G18403,G18404,G18405,G18406,G18407,G18408,G18409,G18410,G18411,G18412,G18413,G18414,G18415,G18416,G18417,G18418,G18419,G18420,
       G18421,G18422,G18423,G18424,G18425,G18426,G18427,G18428,G18429,G18430,G18431,G18432,G18433,G18434,G18435,G18436,G18437,G18438,G18439,G18440,
       G18441,G18442,G18443,G18444,G18445,G18446,G18447,G18448,G18449,G18450,G18451,G18452,G18453,G18454,G18455,G18456,G18457,G18458,G18459,G18460,
       G18461,G18462,G18463,G18464,G18465,G18466,G18467,G18468,G18469,G18470,G18471,G18472,G18473,G18474,G18475,G18476,G18477,G18478,G18479,G18480,
       G18481,G18482,G18483,G18484,G18485,G18486,G18487,G18488,G18489,G18490,G18491,G18492,G18493,G18494,G18495,G18496,G18497,G18498,G18499,G18500,
       G18501,G18502,G18503,G18504,G18505,G18506,G18507,G18508,G18509,G18510,G18511,G18512,G18513,G18514,G18515,G18516,G18517,G18518,G18519,G18520,
       G18521,G18522,G18523,G18524,G18525,G18526,G18527,G18528,G18529,G18530,G18531,G18532,G18533,G18534,G18535,G18536,G18537,G18538,G18539,G18540,
       G18541,G18542,G18543,G18544,G18545,G18546,G18547,G18548,G18549,G18550,G18551,G18552,G18553,G18554,G18555,G18556,G18557,G18558,G18559,G18560,
       G18561,G18562,G18563,G18564,G18565,G18566,G18567,G18568,G18569,G18570,G18571,G18572,G18573,G18574,G18575,G18576,G18577,G18578,G18579,G18580,
       G18581,G18582,G18583,G18584,G18585,G18586,G18587,G18588,G18589,G18590,G18591,G18592,G18593,G18594,G18595,G18596,G18597,G18598,G18599,G18600,
       G18601,G18602,G18603,G18604,G18605,G18606,G18607,G18608,G18609,G18610,G18611,G18612,G18613,G18614,G18615,G18616,G18617,G18618,G18619,G18620,
       G18621,G18622,G18623,G18624,G18625,G18626,G18627,G18628,G18629,G18630,G18631,G18632,G18633,G18634,G18635,G18636,G18637,G18638,G18639,G18640,
       G18641,G18642,G18643,G18644,G18645,G18646,G18647,G18648,G18649,G18650,G18651,G18652,G18653,G18654,G18655,G18656,G18657,G18658,G18659,G18660,
       G18661,G18662,G18663,G18664,G18665,G18666,G18667,G18668,G18669,G18670,G18671,G18672,G18673,G18674,G18675,G18676,G18677,G18678,G18679,G18680,
       G18681,G18682,G18683,G18684,G18685,G18686,G18687,G18688,G18689,G18690,G18691,G18692,G18693,G18694,G18695,G18696,G18697,G18698,G18699,G18700,
       G18701,G18702,G18703,G18704,G18705,G18706,G18707,G18708,G18709,G18710,G18711,G18712,G18713,G18714,G18715,G18716,G18717,G18718,G18719,G18720,
       G18721,G18722,G18723,G18724,G18725,G18726,G18727,G18728,G18729,G18730,G18731,G18732,G18733,G18734,G18735,G18736,G18737,G18738,G18739,G18740,
       G18741,G18742,G18743,G18744,G18745,G18746,G18747,G18748,G18749,G18750,G18751,G18752,G18753,G18754,G18755,G18756,G18757,G18758,G18759,G18760,
       G18761,G18762,G18763,G18764,G18765,G18766,G18767,G18768,G18769,G18770,G18771,G18772,G18773,G18774,G18775,G18776,G18777,G18778,G18779,G18780,
       G18781,G18782,G18783,G18784,G18785,G18786,G18787,G18788,G18789,G18790,G18791,G18792,G18793,G18794,G18795,G18796,G18797,G18798,G18799,G18800,
       G18801,G18802,G18803,G18804,G18805,G18806,G18807,G18808,G18809,G18810,G18811,G18812,G18813,G18814,G18815,G18816,G18817,G18818,G18819,G18820,
       G18821,G18822,G18823,G18824,G18825,G18826,G18827,G18828,G18829,G18830,G18831,G18832,G18833,G18834,G18835,G18836,G18837,G18838,G18839,G18840,
       G18841,G18842,G18843,G18844,G18845,G18846,G18847,G18848,G18849,G18850,G18851,G18852,G18853,G18854,G18855,G18856,G18857,G18858,G18859,G18860,
       G18861,G18862,G18863,G18864,G18865,G18866,G18867,G18868,G18869,G18870,G18871,G18872,G18873,G18874,G18875,G18876,G18877,G18878,G18879,G18880,
       G18881,G18882,G18883,G18884,G18885,G18886,G18887,G18888,G18889,G18890,G18891,G18892,G18893,G18894,G18895,G18896,G18897,G18898,G18899,G18900,
       G18901,G18902,G18903,G18904,G18905,G18906,G18907,G18908,G18909,G18910,G18911,G18912,G18913,G18914,G18915,G18916,G18917,G18918,G18919,G18920,
       G18921,G18922,G18923,G18924,G18925,G18926,G18927,G18928,G18929,G18930,G18931,G18932,G18933,G18934,G18935,G18936,G18937,G18938,G18939,G18940,
       G18941,G18942,G18943,G18944,G18945,G18946,G18947,G18948,G18949,G18950,G18951,G18952,G18953,G18954,G18955,G18956,G18957,G18958,G18959,G18960,
       G18961,G18962,G18963,G18964,G18965,G18966,G18967,G18968,G18969,G18970,G18971,G18972,G18973,G18974,G18975,G18976,G18977,G18978,G18979,G18980,
       G18981,G18982,G18983,G18984,G18985,G18986,G18987,G18988,G18989,G18990,G18991,G18992,G18993,G18994,G18995,G18996,G18997,G18998,G18999,G19000,
       G19001,G19002,G19003,G19004,G19005,G19006,G19007,G19008,G19009,G19010,G19011,G19012,G19013,G19014,G19015,G19016,G19017,G19018,G19019,G19020,
       G19021,G19022,G19023,G19024,G19025,G19026,G19027,G19028,G19029,G19030,G19031,G19032,G19033,G19034,G19035,G19036,G19037,G19038,G19039,G19040,
       G19041,G19042,G19043,G19044,G19045,G19046,G19047,G19048,G19049,G19050,G19051,G19052,G19053,G19054,G19055,G19056,G19057,G19058,G19059,G19060,
       G19061,G19062,G19063,G19064,G19065,G19066,G19067,G19068,G19069,G19070,G19071,G19072,G19073,G19074,G19075,G19076,G19077,G19078,G19079,G19080,
       G19081,G19082,G19083,G19084,G19085,G19086,G19087,G19088,G19089,G19090,G19091,G19092,G19093,G19094,G19095,G19096,G19097,G19098,G19099,G19100,
       G19101,G19102,G19103,G19104,G19105,G19106,G19107,G19108,G19109,G19110,G19111,G19112,G19113,G19114,G19115,G19116,G19117,G19118,G19119,G19120,
       G19121,G19122,G19123,G19124,G19125,G19126,G19127,G19128,G19129,G19130,G19131,G19132,G19133,G19134,G19135,G19136,G19137,G19138,G19139,G19140,
       G19141,G19142,G19143,G19144,G19145,G19146,G19147,G19148,G19149,G19150,G19151,G19152,G19153,G19154,G19155,G19156,G19157,G19158,G19159,G19160,
       G19161,G19162,G19163,G19164,G19165,G19166,G19167,G19168,G19169,G19170,G19171,G19172,G19173,G19174,G19175,G19176,G19177,G19178,G19179,G19180,
       G19181,G19182,G19183,G19184,G19185,G19186,G19187,G19188,G19189,G19190,G19191,G19192,G19193,G19194,G19195,G19196,G19197,G19198,G19199,G19200,
       G19201,G19202,G19203,G19204,G19205,G19206,G19207,G19208,G19209,G19210,G19211,G19212,G19213,G19214,G19215,G19216,G19217,G19218,G19219,G19220,
       G19221,G19222,G19223,G19224,G19225,G19226,G19227,G19228,G19229,G19230,G19231,G19232,G19233,G19234,G19235,G19236,G19237,G19238,G19239,G19240,
       G19241,G19242,G19243,G19244,G19245,G19246,G19247,G19248,G19249,G19250,G19251,G19252,G19253,G19254,G19255,G19256,G19257,G19258,G19259,G19260,
       G19261,G19262,G19263,G19264,G19265,G19266,G19267,G19268,G19269,G19270,G19271,G19272,G19273,G19274,G19275,G19276,G19277,G19278,G19279,G19280,
       G19281,G19282,G19283,G19284,G19285,G19286,G19287,G19288,G19289,G19290,G19291,G19292,G19293,G19294,G19295,G19296,G19297,G19298,G19299,G19300,
       G19301,G19302,G19303,G19304,G19305,G19306,G19307,G19308,G19309,G19310,G19311,G19312,G19313,G19314,G19315,G19316,G19317,G19318,G19319,G19320,
       G19321,G19322,G19323,G19324,G19325,G19326,G19327,G19328,G19329,G19330,G19331,G19332,G19333,G19334,G19335,G19336,G19337,G19338,G19339,G19340,
       G19341,G19342,G19343,G19344,G19345,G19346,G19347,G19348,G19349,G19350,G19351,G19352,G19353,G19354,G19355,G19356,G19357,G19358,G19359,G19360,
       G19361,G19362,G19363,G19364,G19365,G19366,G19367,G19368,G19369,G19370,G19371,G19372,G19373,G19374,G19375,G19376,G19377,G19378,G19379,G19380,
       G19381,G19382,G19383,G19384,G19385,G19386,G19387,G19388,G19389,G19390,G19391,G19392,G19393,G19394,G19395,G19396,G19397,G19398,G19399,G19400,
       G19401,G19402,G19403,G19404,G19405,G19406,G19407,G19408,G19409,G19410,G19411,G19412,G19413,G19414,G19415,G19416,G19417,G19418,G19419,G19420,
       G19421,G19422,G19423,G19424,G19425,G19426,G19427,G19428,G19429,G19430,G19431,G19432,G19433,G19434,G19435,G19436,G19437,G19438,G19439,G19440,
       G19441,G19442,G19443,G19444,G19445,G19446,G19447,G19448,G19449,G19450,G19451,G19452,G19453,G19454,G19455,G19456,G19457,G19458,G19459,G19460,
       G19461,G19462,G19463,G19464,G19465,G19466,G19467,G19468,G19469,G19470,G19471,G19472,G19473,G19474,G19475,G19476,G19477,G19478,G19479,G19480,
       G19481,G19482,G19483,G19484,G19485,G19486,G19487,G19488,G19489,G19490,G19491,G19492,G19493,G19494,G19495,G19496,G19497,G19498,G19499,G19500,
       G19501,G19502,G19503,G19504,G19505,G19506,G19507,G19508,G19509,G19510,G19511,G19512,G19513,G19514,G19515,G19516,G19517,G19518,G19519,G19520,
       G19521,G19522,G19523,G19524,G19525,G19526,G19527,G19528,G19529,G19530,G19531,G19532,G19533,G19534,G19535,G19536,G19537,G19538,G19539,G19540,
       G19541,G19542,G19543,G19544,G19545,G19546,G19547,G19548,G19549,G19550,G19551,G19552,G19553,G19554,G19555,G19556,G19557,G19558,G19559,G19560,
       G19561,G19562,G19563,G19564,G19565,G19566,G19567,G19568,G19569,G19570,G19571,G19572,G19573,G19574,G19575,G19576,G19577,G19578,G19579,G19580,
       G19581,G19582,G19583,G19584,G19585,G19586,G19587,G19588,G19589,G19590,G19591,G19592,G19593,G19594,G19595,G19596,G19597,G19598,G19599,G19600,
       G19601,G19602,G19603,G19604,G19605,G19606,G19607,G19608,G19609,G19610,G19611,G19612,G19613,G19614,G19615,G19616,G19617,G19618,G19619,G19620,
       G19621,G19622,G19623,G19624,G19625,G19626,G19627,G19628,G19629,G19630,G19631,G19632,G19633,G19634,G19635,G19636,G19637,G19638,G19639,G19640,
       G19641,G19642,G19643,G19644,G19645,G19646,G19647,G19648,G19649,G19650,G19651,G19652,G19653,G19654,G19655,G19656,G19657,G19658,G19659,G19660,
       G19661,G19662,G19663,G19664,G19665,G19666,G19667,G19668,G19669,G19670,G19671,G19672,G19673,G19674,G19675,G19676,G19677,G19678,G19679,G19680,
       G19681,G19682,G19683,G19684,G19685,G19686,G19687,G19688,G19689,G19690,G19691,G19692,G19693,G19694,G19695,G19696,G19697,G19698,G19699,G19700,
       G19701,G19702,G19703,G19704,G19705,G19706,G19707,G19708,G19709,G19710,G19711,G19712,G19713,G19714,G19715,G19716,G19717,G19718,G19719,G19720,
       G19721,G19722,G19723,G19724,G19725,G19726,G19727,G19728,G19729,G19730,G19731,G19732,G19733,G19734,G19735,G19736,G19737,G19738,G19739,G19740,
       G19741,G19742,G19743,G19744,G19745,G19746,G19747,G19748,G19749,G19750,G19751,G19752,G19753,G19754,G19755,G19756,G19757,G19758,G19759,G19760,
       G19761,G19762,G19763,G19764,G19765,G19766,G19767,G19768,G19769,G19770,G19771,G19772,G19773,G19774,G19775,G19776,G19777,G19778,G19779,G19780,
       G19781,G19782,G19783,G19784,G19785,G19786,G19787,G19788,G19789,G19790,G19791,G19792,G19793,G19794,G19795,G19796,G19797,G19798,G19799,G19800,
       G19801,G19802,G19803,G19804,G19805,G19806,G19807,G19808,G19809,G19810,G19811,G19812,G19813,G19814,G19815,G19816,G19817,G19818,G19819,G19820,
       G19821,G19822,G19823,G19824,G19825,G19826,G19827,G19828,G19829,G19830,G19831,G19832,G19833,G19834,G19835,G19836,G19837,G19838,G19839,G19840,
       G19841,G19842,G19843,G19844,G19845,G19846,G19847,G19848,G19849,G19850,G19851,G19852,G19853,G19854,G19855,G19856,G19857,G19858,G19859,G19860,
       G19861,G19862,G19863,G19864,G19865,G19866,G19867,G19868,G19869,G19870,G19871,G19872,G19873,G19874,G19875,G19876,G19877,G19878,G19879,G19880,
       G19881,G19882,G19883,G19884,G19885,G19886,G19887,G19888,G19889,G19890,G19891,G19892,G19893,G19894,G19895,G19896,G19897,G19898,G19899,G19900,
       G19901,G19902,G19903,G19904,G19905,G19906,G19907,G19908,G19909,G19910,G19911,G19912,G19913,G19914,G19915,G19916,G19917,G19918,G19919,G19920,
       G19921,G19922,G19923,G19924,G19925,G19926,G19927,G19928,G19929,G19930,G19931,G19932,G19933,G19934,G19935,G19936,G19937,G19938,G19939,G19940,
       G19941,G19942,G19943,G19944,G19945,G19946,G19947,G19948,G19949,G19950,G19951,G19952,G19953,G19954,G19955,G19956,G19957,G19958,G19959,G19960,
       G19961,G19962,G19963,G19964,G19965,G19966,G19967,G19968,G19969,G19970,G19971,G19972,G19973,G19974,G19975,G19976,G19977,G19978,G19979,G19980,
       G19981,G19982,G19983,G19984,G19985,G19986,G19987,G19988,G19989,G19990,G19991,G19992,G19993,G19994,G19995,G19996,G19997,G19998,G19999,G20000,
       G20001,G20002,G20003,G20004,G20005,G20006,G20007,G20008,G20009,G20010,G20011,G20012,G20013,G20014,G20015,G20016,G20017,G20018,G20019,G20020,
       G20021,G20022,G20023,G20024,G20025,G20026,G20027,G20028,G20029,G20030,G20031,G20032,G20033,G20034,G20035,G20036,G20037,G20038,G20039,G20040,
       G20041,G20042,G20043,G20044,G20045,G20046,G20047,G20048,G20049,G20050,G20051,G20052,G20053,G20054,G20055,G20056,G20057,G20058,G20059,G20060,
       G20061,G20062,G20063,G20064,G20065,G20066,G20067,G20068,G20069,G20070,G20071,G20072,G20073,G20074,G20075,G20076,G20077,G20078,G20079,G20080,
       G20081,G20082,G20083,G20084,G20085,G20086,G20087,G20088,G20089,G20090,G20091,G20092,G20093,G20094,G20095,G20096,G20097,G20098,G20099,G20100,
       G20101,G20102,G20103,G20104,G20105,G20106,G20107,G20108,G20109,G20110,G20111,G20112,G20113,G20114,G20115,G20116,G20117,G20118,G20119,G20120,
       G20121,G20122,G20123,G20124,G20125,G20126,G20127,G20128,G20129,G20130,G20131,G20132,G20133,G20134,G20135,G20136,G20137,G20138,G20139,G20140,
       G20141,G20142,G20143,G20144,G20145,G20146,G20147,G20148,G20149,G20150,G20151,G20152,G20153,G20154,G20155,G20156,G20157,G20158,G20159,G20160,
       G20161,G20162,G20163,G20164,G20165,G20166,G20167,G20168,G20169,G20170,G20171,G20172,G20173,G20174,G20175,G20176,G20177,G20178,G20179,G20180,
       G20181,G20182,G20183,G20184,G20185,G20186,G20187,G20188,G20189,G20190,G20191,G20192,G20193,G20194,G20195,G20196,G20197,G20198,G20199,G20200,
       G20201,G20202,G20203,G20204,G20205,G20206,G20207,G20208,G20209,G20210,G20211,G20212,G20213,G20214,G20215,G20216,G20217,G20218,G20219,G20220,
       G20221,G20222,G20223,G20224,G20225,G20226,G20227,G20228,G20229,G20230,G20231,G20232,G20233,G20234,G20235,G20236,G20237,G20238,G20239,G20240,
       G20241,G20242,G20243,G20244,G20245,G20246,G20247,G20248,G20249,G20250,G20251,G20252,G20253,G20254,G20255,G20256,G20257,G20258,G20259,G20260,
       G20261,G20262,G20263,G20264,G20265,G20266,G20267,G20268,G20269,G20270,G20271,G20272,G20273,G20274,G20275,G20276,G20277,G20278,G20279,G20280,
       G20281,G20282,G20283,G20284,G20285,G20286,G20287,G20288,G20289,G20290,G20291,G20292,G20293,G20294,G20295,G20296,G20297,G20298,G20299,G20300,
       G20301,G20302,G20303,G20304,G20305,G20306,G20307,G20308,G20309,G20310,G20311,G20312,G20313,G20314,G20315,G20316,G20317,G20318,G20319,G20320,
       G20321,G20322,G20323,G20324,G20325,G20326,G20327,G20328,G20329,G20330,G20331,G20332,G20333,G20334,G20335,G20336,G20337,G20338,G20339,G20340,
       G20341,G20342,G20343,G20344,G20345,G20346,G20347,G20348,G20349,G20350,G20351,G20352,G20353,G20354,G20355,G20356,G20357,G20358,G20359,G20360,
       G20361,G20362,G20363,G20364,G20365,G20366,G20367,G20368,G20369,G20370,G20371,G20372,G20373,G20374,G20375,G20376,G20377,G20378,G20379,G20380,
       G20381,G20382,G20383,G20384,G20385,G20386,G20387,G20388,G20389,G20390,G20391,G20392,G20393,G20394,G20395,G20396,G20397,G20398,G20399,G20400,
       G20401,G20402,G20403,G20404,G20405,G20406,G20407,G20408,G20409,G20410,G20411,G20412,G20413,G20414,G20415,G20416,G20417,G20418,G20419,G20420,
       G20421,G20422,G20423,G20424,G20425,G20426,G20427,G20428,G20429,G20430,G20431,G20432,G20433,G20434,G20435,G20436,G20437,G20438,G20439,G20440,
       G20441,G20442,G20443,G20444,G20445,G20446,G20447,G20448,G20449,G20450,G20451,G20452,G20453,G20454,G20455,G20456,G20457,G20458,G20459,G20460,
       G20461,G20462,G20463,G20464,G20465,G20466,G20467,G20468,G20469,G20470,G20471,G20472,G20473,G20474,G20475,G20476,G20477,G20478,G20479,G20480,
       G20481,G20482,G20483,G20484,G20485,G20486,G20487,G20488,G20489,G20490,G20491,G20492,G20493,G20494,G20495,G20496,G20497,G20498,G20499,G20500,
       G20501,G20502,G20503,G20504,G20505,G20506,G20507,G20508,G20509,G20510,G20511,G20512,G20513,G20514,G20515,G20516,G20517,G20518,G20519,G20520,
       G20521,G20522,G20523,G20524,G20525,G20526,G20527,G20528,G20529,G20530,G20531,G20532,G20533,G20534,G20535,G20536,G20537,G20538,G20539,G20540,
       G20541,G20542,G20543,G20544,G20545,G20546,G20547,G20548,G20549,G20550,G20551,G20552,G20553,G20554,G20555,G20556,G20557,G20558,G20559,G20560,
       G20561,G20562,G20563,G20564,G20565,G20566,G20567,G20568,G20569,G20570,G20571,G20572,G20573,G20574,G20575,G20576,G20577,G20578,G20579,G20580,
       G20581,G20582,G20583,G20584,G20585,G20586,G20587,G20588,G20589,G20590,G20591,G20592,G20593,G20594,G20595,G20596,G20597,G20598,G20599,G20600,
       G20601,G20602,G20603,G20604,G20605,G20606,G20607,G20608,G20609,G20610,G20611,G20612,G20613,G20614,G20615,G20616,G20617,G20618,G20619,G20620,
       G20621,G20622,G20623,G20624,G20625,G20626,G20627,G20628,G20629,G20630,G20631,G20632,G20633,G20634,G20635,G20636,G20637,G20638,G20639,G20640,
       G20641,G20642,G20643,G20644,G20645,G20646,G20647,G20648,G20649,G20650,G20651,G20652,G20653,G20654,G20655,G20656,G20657,G20658,G20659,G20660,
       G20661,G20662,G20663,G20664,G20665,G20666,G20667,G20668,G20669,G20670,G20671,G20672,G20673,G20674,G20675,G20676,G20677,G20678,G20679,G20680,
       G20681,G20682,G20683,G20684,G20685,G20686,G20687,G20688,G20689,G20690,G20691,G20692,G20693,G20694,G20695,G20696,G20697,G20698,G20699,G20700,
       G20701,G20702,G20703,G20704,G20705,G20706,G20707,G20708,G20709,G20710,G20711,G20712,G20713,G20714,G20715,G20716,G20717,G20718,G20719,G20720,
       G20721,G20722,G20723,G20724,G20725,G20726,G20727,G20728,G20729,G20730,G20731,G20732,G20733,G20734,G20735,G20736,G20737,G20738,G20739,G20740,
       G20741,G20742,G20743,G20744,G20745,G20746,G20747,G20748,G20749,G20750,G20751,G20752,G20753,G20754,G20755,G20756,G20757,G20758,G20759,G20760,
       G20761,G20762,G20763,G20764,G20765,G20766,G20767,G20768,G20769,G20770,G20771,G20772,G20773,G20774,G20775,G20776,G20777,G20778,G20779,G20780,
       G20781,G20782,G20783,G20784,G20785,G20786,G20787,G20788,G20789,G20790,G20791,G20792,G20793,G20794,G20795,G20796,G20797,G20798,G20799,G20800,
       G20801,G20802,G20803,G20804,G20805,G20806,G20807,G20808,G20809,G20810,G20811,G20812,G20813,G20814,G20815,G20816,G20817,G20818,G20819,G20820,
       G20821,G20822,G20823,G20824,G20825,G20826,G20827,G20828,G20829,G20830,G20831,G20832,G20833,G20834,G20835,G20836,G20837,G20838,G20839,G20840,
       G20841,G20842,G20843,G20844,G20845,G20846,G20847,G20848,G20849,G20850,G20851,G20852,G20853,G20854,G20855,G20856,G20857,G20858,G20859,G20860,
       G20861,G20862,G20863,G20864,G20865,G20866,G20867,G20868,G20869,G20870,G20871,G20872,G20873,G20874,G20875,G20876,G20877,G20878,G20879,G20880,
       G20881,G20882,G20883,G20884,G20885,G20886,G20887,G20888,G20889,G20890,G20891,G20892,G20893,G20894,G20895,G20896,G20897,G20898,G20899,G20900,
       G20901,G20902,G20903,G20904,G20905,G20906,G20907,G20908,G20909,G20910,G20911,G20912,G20913,G20914,G20915,G20916,G20917,G20918,G20919,G20920,
       G20921,G20922,G20923,G20924,G20925,G20926,G20927,G20928,G20929,G20930,G20931,G20932,G20933,G20934,G20935,G20936,G20937,G20938,G20939,G20940,
       G20941,G20942,G20943,G20944,G20945,G20946,G20947,G20948,G20949,G20950,G20951,G20952,G20953,G20954,G20955,G20956,G20957,G20958,G20959,G20960,
       G20961,G20962,G20963,G20964,G20965,G20966,G20967,G20968,G20969,G20970,G20971,G20972,G20973,G20974,G20975,G20976,G20977,G20978,G20979,G20980,
       G20981,G20982,G20983,G20984,G20985,G20986,G20987,G20988,G20989,G20990,G20991,G20992,G20993,G20994,G20995,G20996,G20997,G20998,G20999,G21000,
       G21001,G21002,G21003,G21004,G21005,G21006,G21007,G21008,G21009,G21010,G21011,G21012,G21013,G21014,G21015,G21016,G21017,G21018,G21019,G21020,
       G21021,G21022,G21023,G21024,G21025,G21026,G21027,G21028,G21029,G21030,G21031,G21032,G21033,G21034,G21035,G21036,G21037,G21038,G21039,G21040,
       G21041,G21042,G21043,G21044,G21045,G21046,G21047,G21048,G21049,G21050,G21051,G21052,G21053,G21054,G21055,G21056,G21057,G21058,G21059,G21060,
       G21061,G21062,G21063,G21064,G21065,G21066,G21067,G21068,G21069,G21070,G21071,G21072,G21073,G21074,G21075,G21076,G21077,G21078,G21079,G21080,
       G21081,G21082,G21083,G21084,G21085,G21086,G21087,G21088,G21089,G21090,G21091,G21092,G21093,G21094,G21095,G21096,G21097,G21098,G21099,G21100,
       G21101,G21102,G21103,G21104,G21105,G21106,G21107,G21108,G21109,G21110,G21111,G21112,G21113,G21114,G21115,G21116,G21117,G21118,G21119,G21120,
       G21121,G21122,G21123,G21124,G21125,G21126,G21127,G21128,G21129,G21130,G21131,G21132,G21133,G21134,G21135,G21136,G21137,G21138,G21139,G21140,
       G21141,G21142,G21143,G21144,G21145,G21146,G21147,G21148,G21149,G21150,G21151,G21152,G21153,G21154,G21155,G21156,G21157,G21158,G21159,G21160,
       G21161,G21162,G21163,G21164,G21165,G21166,G21167,G21168,G21169,G21170,G21171,G21172,G21173,G21174,G21175,G21176,G21177,G21178,G21179,G21180,
       G21181,G21182,G21183,G21184,G21185,G21186,G21187,G21188,G21189,G21190,G21191,G21192,G21193,G21194,G21195,G21196,G21197,G21198,G21199,G21200,
       G21201,G21202,G21203,G21204,G21205,G21206,G21207,G21208,G21209,G21210,G21211,G21212,G21213,G21214,G21215,G21216,G21217,G21218,G21219,G21220,
       G21221,G21222,G21223,G21224,G21225,G21226,G21227,G21228,G21229,G21230,G21231,G21232,G21233,G21234,G21235,G21236,G21237,G21238,G21239,G21240,
       G21241,G21242,G21243,G21244,G21245,G21246,G21247,G21248,G21249,G21250,G21251,G21252,G21253,G21254,G21255,G21256,G21257,G21258,G21259,G21260,
       G21261,G21262,G21263,G21264,G21265,G21266,G21267,G21268,G21269,G21270,G21271,G21272,G21273,G21274,G21275,G21276,G21277,G21278,G21279,G21280,
       G21281,G21282,G21283,G21284,G21285,G21286,G21287,G21288,G21289,G21290,G21291,G21292,G21293,G21294,G21295,G21296,G21297,G21298,G21299,G21300,
       G21301,G21302,G21303,G21304,G21305,G21306,G21307,G21308,G21309,G21310,G21311,G21312,G21313,G21314,G21315,G21316,G21317,G21318,G21319,G21320,
       G21321,G21322,G21323,G21324,G21325,G21326,G21327,G21328,G21329,G21330,G21331,G21332,G21333,G21334,G21335,G21336,G21337,G21338,G21339,G21340,
       G21341,G21342,G21343,G21344,G21345,G21346,G21347,G21348,G21349,G21350,G21351,G21352,G21353,G21354,G21355,G21356,G21357,G21358,G21359,G21360,
       G21361,G21362,G21363,G21364,G21365,G21366,G21367,G21368,G21369,G21370,G21371,G21372,G21373,G21374,G21375,G21376,G21377,G21378,G21379,G21380,
       G21381,G21382,G21383,G21384,G21385,G21386,G21387,G21388,G21389,G21390,G21391,G21392,G21393,G21394,G21395,G21396,G21397,G21398,G21399,G21400,
       G21401,G21402,G21403,G21404,G21405,G21406,G21407,G21408,G21409,G21410,G21411,G21412,G21413,G21414,G21415,G21416,G21417,G21418,G21419,G21420,
       G21421,G21422,G21423,G21424,G21425,G21426,G21427,G21428,G21429,G21430,G21431,G21432,G21433,G21434,G21435,G21436,G21437,G21438,G21439,G21440,
       G21441,G21442,G21443,G21444,G21445,G21446,G21447,G21448,G21449,G21450,G21451,G21452,G21453,G21454,G21455,G21456,G21457,G21458,G21459,G21460,
       G21461,G21462,G21463,G21464,G21465,G21466,G21467,G21468,G21469,G21470,G21471,G21472,G21473,G21474,G21475,G21476,G21477,G21478,G21479,G21480,
       G21481,G21482,G21483,G21484,G21485,G21486,G21487,G21488,G21489,G21490,G21491,G21492,G21493,G21494,G21495,G21496,G21497,G21498,G21499,G21500,
       G21501,G21502,G21503,G21504,G21505,G21506,G21507,G21508,G21509,G21510,G21511,G21512,G21513,G21514,G21515,G21516,G21517,G21518,G21519,G21520,
       G21521,G21522,G21523,G21524,G21525,G21526,G21527,G21528,G21529,G21530,G21531,G21532,G21533,G21534,G21535,G21536,G21537,G21538,G21539,G21540,
       G21541,G21542,G21543,G21544,G21545,G21546,G21547,G21548,G21549,G21550,G21551,G21552,G21553,G21554,G21555,G21556,G21557,G21558,G21559,G21560,
       G21561,G21562,G21563,G21564,G21565,G21566,G21567,G21568,G21569,G21570,G21571,G21572,G21573,G21574,G21575,G21576,G21577,G21578,G21579,G21580,
       G21581,G21582,G21583,G21584,G21585,G21586,G21587,G21588,G21589,G21590,G21591,G21592,G21593,G21594,G21595,G21596,G21597,G21598,G21599,G21600,
       G21601,G21602,G21603,G21604,G21605,G21606,G21607,G21608,G21609,G21610,G21611,G21612,G21613,G21614,G21615,G21616,G21617,G21618,G21619,G21620,
       G21621,G21622,G21623,G21624,G21625,G21626,G21627,G21628,G21629,G21630,G21631,G21632,G21633,G21634,G21635,G21636,G21637,G21638,G21639,G21640,
       G21641,G21642,G21643,G21644,G21645,G21646,G21647,G21648,G21649,G21650,G21651,G21652,G21653,G21654,G21655,G21656,G21657,G21658,G21659,G21660,
       G21661,G21662,G21663,G21664,G21665,G21666,G21667,G21668,G21669,G21670,G21671,G21672,G21673,G21674,G21675,G21676,G21677,G21678,G21679,G21680,
       G21681,G21682,G21683,G21684,G21685,G21686,G21687,G21688,G21689,G21690,G21691,G21692,G21693,G21694,G21695,G21696,G21697,G21698,G21699,G21700,
       G21701,G21702,G21703,G21704,G21705,G21706,G21707,G21708,G21709,G21710,G21711,G21712,G21713,G21714,G21715,G21716,G21717,G21718,G21719,G21720,
       G21721,G21722,G21723,G21724,G21725,G21726,G21727,G21728,G21729,G21730,G21731,G21732,G21733,G21734,G21735,G21736,G21737,G21738,G21739,G21740,
       G21741,G21742,G21743,G21744,G21745,G21746,G21747,G21748,G21749,G21750,G21751,G21752,G21753,G21754,G21755,G21756,G21757,G21758,G21759,G21760,
       G21761,G21762,G21763,G21764,G21765,G21766,G21767,G21768,G21769,G21770,G21771,G21772,G21773,G21774,G21775,G21776,G21777,G21778,G21779,G21780,
       G21781,G21782,G21783,G21784,G21785,G21786,G21787,G21788,G21789,G21790,G21791,G21792,G21793,G21794,G21795,G21796,G21797,G21798,G21799,G21800,
       G21801,G21802,G21803,G21804,G21805,G21806,G21807,G21808,G21809,G21810,G21811,G21812,G21813,G21814,G21815,G21816,G21817,G21818,G21819,G21820,
       G21821,G21822,G21823,G21824,G21825,G21826,G21827,G21828,G21829,G21830,G21831,G21832,G21833,G21834,G21835,G21836,G21837,G21838,G21839,G21840,
       G21841,G21842,G21843,G21844,G21845,G21846,G21847,G21848,G21849,G21850,G21851,G21852,G21853,G21854,G21855,G21856,G21857,G21858,G21859,G21860,
       G21861,G21862,G21863,G21864,G21865,G21866,G21867,G21868,G21869,G21870,G21871,G21872,G21873,G21874,G21875,G21876,G21877,G21878,G21879,G21880,
       G21881,G21882,G21883,G21884,G21885,G21886,G21887,G21888,G21889,G21890,G21891,G21892,G21893,G21894,G21895,G21896,G21897,G21898,G21899,G21900,
       G21901,G21902,G21903,G21904,G21905,G21906,G21907,G21908,G21909,G21910,G21911,G21912,G21913,G21914,G21915,G21916,G21917,G21918,G21919,G21920,
       G21921,G21922,G21923,G21924,G21925,G21926,G21927,G21928,G21929,G21930,G21931,G21932,G21933,G21934,G21935,G21936,G21937,G21938,G21939,G21940,
       G21941,G21942,G21943,G21944,G21945,G21946,G21947,G21948,G21949,G21950,G21951,G21952,G21953,G21954,G21955,G21956,G21957,G21958,G21959,G21960,
       G21961,G21962,G21963,G21964,G21965,G21966,G21967,G21968,G21969,G21970,G21971,G21972,G21973,G21974,G21975,G21976,G21977,G21978,G21979,G21980,
       G21981,G21982,G21983,G21984,G21985,G21986,G21987,G21988,G21989,G21990,G21991,G21992,G21993,G21994,G21995,G21996,G21997,G21998,G21999,G22000,
       G22001,G22002,G22003,G22004,G22005,G22006,G22007,G22008,G22009,G22010,G22011,G22012,G22013,G22014,G22015,G22016,G22017,G22018,G22019,G22020,
       G22021,G22022,G22023,G22024,G22025,G22026,G22027,G22028,G22029,G22030,G22031,G22032,G22033,G22034,G22035,G22036,G22037,G22038,G22039,G22040,
       G22041,G22042,G22043,G22044,G22045,G22046,G22047,G22048,G22049,G22050,G22051,G22052,G22053,G22054,G22055,G22056,G22057,G22058,G22059,G22060,
       G22061,G22062,G22063,G22064,G22065,G22066,G22067,G22068,G22069,G22070,G22071,G22072,G22073,G22074,G22075,G22076,G22077,G22078,G22079,G22080,
       G22081,G22082,G22083,G22084,G22085,G22086,G22087,G22088,G22089,G22090,G22091,G22092,G22093,G22094,G22095,G22096,G22097,G22098,G22099,G22100,
       G22101,G22102,G22103,G22104,G22105,G22106,G22107,G22108,G22109,G22110,G22111,G22112,G22113,G22114,G22115,G22116,G22117,G22118,G22119,G22120,
       G22121,G22122,G22123,G22124,G22125,G22126,G22127,G22128,G22129,G22130,G22131,G22132,G22133,G22134,G22135,G22136,G22137,G22138,G22139,G22140,
       G22141,G22142,G22143,G22144,G22145,G22146,G22147,G22148,G22149,G22150,G22151,G22152,G22153,G22154,G22155,G22156,G22157,G22158,G22159,G22160,
       G22161,G22162,G22163,G22164,G22165,G22166,G22167,G22168,G22169,G22170,G22171,G22172,G22173,G22174,G22175,G22176,G22177,G22178,G22179,G22180,
       G22181,G22182,G22183,G22184,G22185,G22186,G22187,G22188,G22189,G22190,G22191,G22192,G22193,G22194,G22195,G22196,G22197,G22198,G22199,G22200,
       G22201,G22202,G22203,G22204,G22205,G22206,G22207,G22208,G22209,G22210,G22211,G22212,G22213,G22214,G22215,G22216,G22217,G22218,G22219,G22220,
       G22221,G22222,G22223,G22224,G22225,G22226,G22227,G22228,G22229,G22230,G22231,G22232,G22233,G22234,G22235,G22236,G22237,G22238,G22239,G22240,
       G22241,G22242,G22243,G22244,G22245,G22246,G22247,G22248,G22249,G22250,G22251,G22252,G22253,G22254,G22255,G22256,G22257,G22258,G22259,G22260,
       G22261,G22262,G22263,G22264,G22265,G22266,G22267,G22268,G22269,G22270,G22271,G22272,G22273,G22274,G22275,G22276,G22277,G22278,G22279,G22280,
       G22281,G22282,G22283,G22284,G22285,G22286,G22287,G22288,G22289,G22290,G22291,G22292,G22293,G22294,G22295,G22296,G22297,G22298,G22299,G22300,
       G22301,G22302,G22303,G22304,G22305,G22306,G22307,G22308,G22309,G22310,G22311,G22312,G22313,G22314,G22315,G22316,G22317,G22318,G22319,G22320,
       G22321,G22322,G22323,G22324,G22325,G22326,G22327,G22328,G22329,G22330,G22331,G22332,G22333,G22334,G22335,G22336,G22337,G22338,G22339,G22340,
       G22341,G22342,G22343,G22344,G22345,G22346,G22347,G22348,G22349,G22350,G22351,G22352,G22353,G22354,G22355,G22356,G22357,G22358,G22359,G22360,
       G22361,G22362,G22363,G22364,G22365,G22366,G22367,G22368,G22369,G22370,G22371,G22372,G22373,G22374,G22375,G22376,G22377,G22378,G22379,G22380,
       G22381,G22382,G22383,G22384,G22385,G22386,G22387,G22388,G22389,G22390,G22391,G22392,G22393,G22394,G22395,G22396,G22397,G22398,G22399,G22400,
       G22401,G22402,G22403,G22404,G22405,G22406,G22407,G22408,G22409,G22410,G22411,G22412,G22413,G22414,G22415,G22416,G22417,G22418,G22419,G22420,
       G22421,G22422,G22423,G22424,G22425,G22426,G22427,G22428,G22429,G22430,G22431,G22432,G22433,G22434,G22435,G22436,G22437,G22438,G22439,G22440,
       G22441,G22442,G22443,G22444,G22445,G22446,G22447,G22448,G22449,G22450,G22451,G22452,G22453,G22454,G22455,G22456,G22457,G22458,G22459,G22460,
       G22461,G22462,G22463,G22464,G22465,G22466,G22467,G22468,G22469,G22470,G22471,G22472,G22473,G22474,G22475,G22476,G22477,G22478,G22479,G22480,
       G22481,G22482,G22483,G22484,G22485,G22486,G22487,G22488,G22489,G22490,G22491,G22492,G22493,G22494,G22495,G22496,G22497,G22498,G22499,G22500,
       G22501,G22502,G22503,G22504,G22505,G22506,G22507,G22508,G22509,G22510,G22511,G22512,G22513,G22514,G22515,G22516,G22517,G22518,G22519,G22520,
       G22521,G22522,G22523,G22524,G22525,G22526,G22527,G22528,G22529,G22530,G22531,G22532,G22533,G22534,G22535,G22536,G22537,G22538,G22539,G22540,
       G22541,G22542,G22543,G22544,G22545,G22546,G22547,G22548,G22549,G22550,G22551,G22552,G22553,G22554,G22555,G22556,G22557,G22558,G22559,G22560,
       G22561,G22562,G22563,G22564,G22565,G22566,G22567,G22568,G22569,G22570,G22571,G22572,G22573,G22574,G22575,G22576,G22577,G22578,G22579,G22580,
       G22581,G22582,G22583,G22584,G22585,G22586,G22587,G22588,G22589,G22590,G22591,G22592,G22593,G22594,G22595,G22596,G22597,G22598,G22599,G22600,
       G22601,G22602,G22603,G22604,G22605,G22606,G22607,G22608,G22609,G22610,G22611,G22612,G22613,G22614,G22615,G22616,G22617,G22618,G22619,G22620,
       G22621,G22622,G22623,G22624,G22625,G22626,G22627,G22628,G22629,G22630,G22631,G22632,G22633,G22634,G22635,G22636,G22637,G22638,G22639,G22640,
       G22641,G22642,G22643,G22644,G22645,G22646,G22647,G22648,G22649,G22650,G22651,G22652,G22653,G22654,G22655,G22656,G22657,G22658,G22659,G22660,
       G22661,G22662,G22663,G22664,G22665,G22666,G22667,G22668,G22669,G22670,G22671,G22672,G22673,G22674,G22675,G22676,G22677,G22678,G22679,G22680,
       G22681,G22682,G22683,G22684,G22685,G22686,G22687,G22688,G22689,G22690,G22691,G22692,G22693,G22694,G22695,G22696,G22697,G22698,G22699,G22700,
       G22701,G22702,G22703,G22704,G22705,G22706,G22707,G22708,G22709,G22710,G22711,G22712,G22713,G22714,G22715,G22716,G22717,G22718,G22719,G22720,
       G22721,G22722,G22723,G22724,G22725,G22726,G22727,G22728,G22729,G22730,G22731,G22732,G22733,G22734,G22735,G22736,G22737,G22738,G22739,G22740,
       G22741,G22742,G22743,G22744,G22745,G22746,G22747,G22748,G22749,G22750,G22751,G22752,G22753,G22754,G22755,G22756,G22757,G22758,G22759,G22760,
       G22761,G22762,G22763,G22764,G22765,G22766,G22767,G22768,G22769,G22770,G22771,G22772,G22773,G22774,G22775,G22776,G22777,G22778,G22779,G22780,
       G22781,G22782,G22783,G22784,G22785,G22786,G22787,G22788,G22789,G22790,G22791,G22792,G22793,G22794,G22795,G22796,G22797,G22798,G22799,G22800,
       G22801,G22802,G22803,G22804,G22805,G22806,G22807,G22808,G22809,G22810,G22811,G22812,G22813,G22814,G22815,G22816,G22817,G22818,G22819,G22820,
       G22821,G22822,G22823,G22824,G22825,G22826,G22827,G22828,G22829,G22830,G22831,G22832,G22833,G22834,G22835,G22836,G22837,G22838,G22839,G22840,
       G22841,G22842,G22843,G22844,G22845,G22846,G22847,G22848,G22849,G22850,G22851,G22852,G22853,G22854,G22855,G22856,G22857,G22858,G22859,G22860,
       G22861,G22862,G22863,G22864,G22865,G22866,G22867,G22868,G22869,G22870,G22871,G22872,G22873,G22874,G22875,G22876,G22877,G22878,G22879,G22880,
       G22881,G22882,G22883,G22884,G22885,G22886,G22887,G22888,G22889,G22890,G22891,G22892,G22893,G22894,G22895,G22896,G22897,G22898,G22899,G22900,
       G22901,G22902,G22903,G22904,G22905,G22906,G22907,G22908,G22909,G22910,G22911,G22912,G22913,G22914,G22915,G22916,G22917,G22918,G22919,G22920,
       G22921,G22922,G22923,G22924,G22925,G22926,G22927,G22928,G22929,G22930,G22931,G22932,G22933,G22934,G22935,G22936,G22937,G22938,G22939,G22940,
       G22941,G22942,G22943,G22944,G22945,G22946,G22947,G22948,G22949,G22950,G22951,G22952,G22953,G22954,G22955,G22956,G22957,G22958,G22959,G22960,
       G22961,G22962,G22963,G22964,G22965,G22966,G22967,G22968,G22969,G22970,G22971,G22972,G22973,G22974,G22975,G22976,G22977,G22978,G22979,G22980,
       G22981,G22982,G22983,G22984,G22985,G22986,G22987,G22988,G22989,G22990,G22991,G22992,G22993,G22994,G22995,G22996,G22997,G22998,G22999,G23000,
       G23001,G23002,G23003,G23004,G23005,G23006,G23007,G23008,G23009,G23010,G23011,G23012,G23013,G23014,G23015,G23016,G23017,G23018,G23019,G23020,
       G23021,G23022,G23023,G23024,G23025,G23026,G23027,G23028,G23029,G23030,G23031,G23032,G23033,G23034,G23035,G23036,G23037,G23038,G23039,G23040,
       G23041,G23042,G23043,G23044,G23045,G23046,G23047,G23048,G23049,G23050,G23051,G23052,G23053,G23054,G23055,G23056,G23057,G23058,G23059,G23060,
       G23061,G23062,G23063,G23064,G23065,G23066,G23067,G23068,G23069,G23070,G23071,G23072,G23073,G23074,G23075,G23076,G23077,G23078,G23079,G23080,
       G23081,G23082,G23083,G23084,G23085,G23086,G23087,G23088,G23089,G23090,G23091,G23092,G23093,G23094,G23095,G23096,G23097,G23098,G23099,G23100,
       G23101,G23102,G23103,G23104,G23105,G23106,G23107,G23108,G23109,G23110,G23111,G23112,G23113,G23114,G23115,G23116,G23117,G23118,G23119,G23120,
       G23121,G23122,G23123,G23124,G23125,G23126,G23127,G23128,G23129,G23130,G23131,G23132,G23133,G23134,G23135,G23136,G23137,G23138,G23139,G23140,
       G23141,G23142,G23143,G23144,G23145,G23146,G23147,G23148,G23149,G23150,G23151,G23152,G23153,G23154,G23155,G23156,G23157,G23158,G23159,G23160,
       G23161,G23162,G23163,G23164,G23165,G23166,G23167,G23168,G23169,G23170,G23171,G23172,G23173,G23174,G23175,G23176,G23177,G23178,G23179,G23180,
       G23181,G23182,G23183,G23184,G23185,G23186,G23187,G23188,G23189,G23190,G23191,G23192,G23193,G23194,G23195,G23196,G23197,G23198,G23199,G23200,
       G23201,G23202,G23203,G23204,G23205,G23206,G23207,G23208,G23209,G23210,G23211,G23212,G23213,G23214,G23215,G23216,G23217,G23218,G23219,G23220,
       G23221,G23222,G23223,G23224,G23225,G23226,G23227,G23228,G23229,G23230,G23231,G23232,G23233,G23234,G23235,G23236,G23237,G23238,G23239,G23240,
       G23241,G23242,G23243,G23244,G23245,G23246,G23247,G23248,G23249,G23250,G23251,G23252,G23253,G23254,G23255,G23256,G23257,G23258,G23259,G23260,
       G23261,G23262,G23263,G23264,G23265,G23266,G23267,G23268,G23269,G23270,G23271,G23272,G23273,G23274,G23275,G23276,G23277,G23278,G23279,G23280,
       G23281,G23282,G23283,G23284,G23285,G23286,G23287,G23288,G23289,G23290,G23291,G23292,G23293,G23294,G23295,G23296,G23297,G23298,G23299,G23300,
       G23301,G23302,G23303,G23304,G23305,G23306,G23307,G23308,G23309,G23310,G23311,G23312,G23313,G23314,G23315,G23316,G23317,G23318,G23319,G23320,
       G23321,G23322,G23323,G23324,G23325,G23326,G23327,G23328,G23329,G23330,G23331,G23332,G23333,G23334,G23335,G23336,G23337,G23338,G23339,G23340,
       G23341,G23342,G23343,G23344,G23345,G23346,G23347,G23348,G23349,G23350,G23351,G23352,G23353,G23354,G23355,G23356,G23357,G23358,G23359,G23360,
       G23361,G23362,G23363,G23364,G23365,G23366,G23367,G23368,G23369,G23370,G23371,G23372,G23373,G23374,G23375,G23376,G23377,G23378,G23379,G23380,
       G23381,G23382,G23383,G23384,G23385,G23386,G23387,G23388,G23389,G23390,G23391,G23392,G23393,G23394,G23395,G23396,G23397,G23398,G23399,G23400,
       G23401,G23402,G23403,G23404,G23405,G23406,G23407,G23408,G23409,G23410,G23411,G23412,G23413,G23414,G23415,G23416,G23417,G23418,G23419,G23420,
       G23421,G23422,G23423,G23424,G23425,G23426,G23427,G23428,G23429,G23430,G23431,G23432,G23433,G23434,G23435,G23436,G23437,G23438,G23439,G23440,
       G23441,G23442,G23443,G23444,G23445,G23446,G23447,G23448,G23449,G23450,G23451,G23452,G23453,G23454,G23455,G23456,G23457,G23458,G23459,G23460,
       G23461,G23462,G23463,G23464,G23465,G23466,G23467,G23468,G23469,G23470,G23471,G23472,G23473,G23474,G23475,G23476,G23477,G23478,G23479,G23480,
       G23481,G23482,G23483,G23484,G23485,G23486,G23487,G23488,G23489,G23490,G23491,G23492,G23493,G23494,G23495,G23496,G23497,G23498,G23499,G23500,
       G23501,G23502,G23503,G23504,G23505,G23506,G23507,G23508,G23509,G23510,G23511,G23512,G23513,G23514,G23515,G23516,G23517,G23518,G23519,G23520,
       G23521,G23522,G23523,G23524,G23525,G23526,G23527,G23528,G23529,G23530,G23531,G23532,G23533,G23534,G23535,G23536,G23537,G23538,G23539,G23540,
       G23541,G23542,G23543,G23544,G23545,G23546,G23547,G23548,G23549,G23550,G23551,G23552,G23553,G23554,G23555,G23556,G23557,G23558,G23559,G23560,
       G23561,G23562,G23563,G23564,G23565,G23566,G23567,G23568,G23569,G23570,G23571,G23572,G23573,G23574,G23575,G23576,G23577,G23578,G23579,G23580,
       G23581,G23582,G23583,G23584,G23585,G23586,G23587,G23588,G23589,G23590,G23591,G23592,G23593,G23594,G23595,G23596,G23597,G23598,G23599,G23600,
       G23601,G23602,G23603,G23604,G23605,G23606,G23607,G23608,G23609,G23610,G23611,G23612,G23613,G23614,G23615,G23616,G23617,G23618,G23619,G23620,
       G23621,G23622,G23623,G23624,G23625,G23626,G23627,G23628,G23629,G23630,G23631,G23632,G23633,G23634,G23635,G23636,G23637,G23638,G23639,G23640,
       G23641,G23642,G23643,G23644,G23645,G23646,G23647,G23648,G23649,G23650,G23651,G23652,G23653,G23654,G23655,G23656,G23657,G23658,G23659,G23660,
       G23661,G23662,G23663,G23664,G23665,G23666,G23667,G23668,G23669,G23670,G23671,G23672,G23673,G23674,G23675,G23676,G23677,G23678,G23679,G23680,
       G23681,G23682,G23683,G23684,G23685,G23686,G23687,G23688,G23689,G23690,G23691,G23692,G23693,G23694,G23695,G23696,G23697,G23698,G23699,G23700,
       G23701,G23702,G23703,G23704,G23705,G23706,G23707,G23708,G23709,G23710,G23711,G23712,G23713,G23714,G23715,G23716,G23717,G23718,G23719,G23720,
       G23721,G23722,G23723,G23724,G23725,G23726,G23727,G23728,G23729,G23730,G23731,G23732,G23733,G23734,G23735,G23736,G23737,G23738,G23739,G23740,
       G23741,G23742,G23743,G23744,G23745,G23746,G23747,G23748,G23749,G23750,G23751,G23752,G23753,G23754,G23755,G23756,G23757,G23758,G23759,G23760,
       G23761,G23762,G23763,G23764,G23765,G23766,G23767,G23768,G23769,G23770,G23771,G23772,G23773,G23774,G23775,G23776,G23777,G23778,G23779,G23780,
       G23781,G23782,G23783,G23784,G23785,G23786,G23787,G23788,G23789,G23790,G23791,G23792,G23793,G23794,G23795,G23796,G23797,G23798,G23799,G23800,
       G23801,G23802,G23803,G23804,G23805,G23806,G23807,G23808,G23809,G23810,G23811,G23812,G23813,G23814,G23815,G23816,G23817,G23818,G23819,G23820,
       G23821,G23822,G23823,G23824,G23825,G23826,G23827,G23828,G23829,G23830,G23831,G23832,G23833,G23834,G23835,G23836,G23837,G23838,G23839,G23840,
       G23841,G23842,G23843,G23844,G23845,G23846,G23847,G23848,G23849,G23850,G23851,G23852,G23853,G23854,G23855,G23856,G23857,G23858,G23859,G23860,
       G23861,G23862,G23863,G23864,G23865,G23866,G23867,G23868,G23869,G23870,G23871,G23872,G23873,G23874,G23875,G23876,G23877,G23878,G23879,G23880,
       G23881,G23882,G23883,G23884,G23885,G23886,G23887,G23888,G23889,G23890,G23891,G23892,G23893,G23894,G23895,G23896,G23897,G23898,G23899,G23900,
       G23901,G23902,G23903,G23904,G23905,G23906,G23907,G23908,G23909,G23910,G23911,G23912,G23913,G23914,G23915,G23916,G23917,G23918,G23919,G23920,
       G23921,G23922,G23923,G23924,G23925,G23926,G23927,G23928,G23929,G23930,G23931,G23932,G23933,G23934,G23935,G23936,G23937,G23938,G23939,G23940,
       G23941,G23942,G23943,G23944,G23945,G23946,G23947,G23948,G23949,G23950,G23951,G23952,G23953,G23954,G23955,G23956,G23957,G23958,G23959,G23960,
       G23961,G23962,G23963,G23964,G23965,G23966,G23967,G23968,G23969,G23970,G23971,G23972,G23973,G23974,G23975,G23976,G23977,G23978,G23979,G23980,
       G23981,G23982,G23983,G23984,G23985,G23986,G23987,G23988,G23989,G23990,G23991,G23992,G23993,G23994,G23995,G23996,G23997,G23998,G23999,G24000,
       G24001,G24002,G24003,G24004,G24005,G24006,G24007,G24008,G24009,G24010,G24011,G24012,G24013,G24014,G24015,G24016,G24017,G24018,G24019,G24020,
       G24021,G24022,G24023,G24024,G24025,G24026,G24027,G24028,G24029,G24030,G24031,G24032,G24033,G24034,G24035,G24036,G24037,G24038,G24039,G24040,
       G24041,G24042,G24043,G24044,G24045,G24046,G24047,G24048,G24049,G24050,G24051,G24052,G24053,G24054,G24055,G24056,G24057,G24058,G24059,G24060,
       G24061,G24062,G24063,G24064,G24065,G24066,G24067,G24068,G24069,G24070,G24071,G24072,G24073,G24074,G24075,G24076,G24077,G24078,G24079,G24080,
       G24081,G24082,G24083,G24084,G24085,G24086,G24087,G24088,G24089,G24090,G24091,G24092,G24093,G24094,G24095,G24096,G24097,G24098,G24099,G24100,
       G24101,G24102,G24103,G24104,G24105,G24106,G24107,G24108,G24109,G24110,G24111,G24112,G24113,G24114,G24115,G24116,G24117,G24118,G24119,G24120,
       G24121,G24122,G24123,G24124,G24125,G24126,G24127,G24128,G24129,G24130,G24131,G24132,G24133,G24134,G24135,G24136,G24137,G24138,G24139,G24140,
       G24141,G24142,G24143,G24144,G24145,G24146,G24147,G24148,G24149,G24150,G24151,G24152,G24153,G24154,G24155,G24156,G24157,G24158,G24159,G24160,
       G24161,G24162,G24163,G24164,G24165,G24166,G24167,G24168,G24169,G24170,G24171,G24172,G24173,G24174,G24175,G24176,G24177,G24178,G24179,G24180,
       G24181,G24182,G24183,G24184,G24185,G24186,G24187,G24188,G24189,G24190,G24191,G24192,G24193,G24194,G24195,G24196,G24197,G24198,G24199,G24200,
       G24201,G24202,G24203,G24204,G24205,G24206,G24207,G24208,G24209,G24210,G24211,G24212,G24213,G24214,G24215,G24216,G24217,G24218,G24219,G24220,
       G24221,G24222,G24223,G24224,G24225,G24226,G24227,G24228,G24229,G24230,G24231,G24232,G24233,G24234,G24235,G24236,G24237,G24238,G24239,G24240,
       G24241,G24242,G24243,G24244,G24245,G24246,G24247,G24248,G24249,G24250,G24251,G24252,G24253,G24254,G24255,G24256,G24257,G24258,G24259,G24260,
       G24261,G24262,G24263,G24264,G24265,G24266,G24267,G24268,G24269,G24270,G24271,G24272,G24273,G24274,G24275,G24276,G24277,G24278,G24279,G24280,
       G24281,G24282,G24283,G24284,G24285,G24286,G24287,G24288,G24289,G24290,G24291,G24292,G24293,G24294,G24295,G24296,G24297,G24298,G24299,G24300,
       G24301,G24302,G24303,G24304,G24305,G24306,G24307,G24308,G24309,G24310,G24311,G24312,G24313,G24314,G24315,G24316,G24317,G24318,G24319,G24320,
       G24321,G24322,G24323,G24324,G24325,G24326,G24327,G24328,G24329,G24330,G24331,G24332,G24333,G24334,G24335,G24336,G24337,G24338,G24339,G24340,
       G24341,G24342,G24343,G24344,G24345,G24346,G24347,G24348,G24349,G24350,G24351,G24352,G24353,G24354,G24355,G24356,G24357,G24358,G24359,G24360,
       G24361,G24362,G24363,G24364,G24365,G24366,G24367,G24368,G24369,G24370,G24371,G24372,G24373,G24374,G24375,G24376,G24377,G24378,G24379,G24380,
       G24381,G24382,G24383,G24384,G24385,G24386,G24387,G24388,G24389,G24390,G24391,G24392,G24393,G24394,G24395,G24396,G24397,G24398,G24399,G24400,
       G24401,G24402,G24403,G24404,G24405,G24406,G24407,G24408,G24409,G24410,G24411,G24412,G24413,G24414,G24415,G24416,G24417,G24418,G24419,G24420,
       G24421,G24422,G24423,G24424,G24425,G24426,G24427,G24428,G24429,G24430,G24431,G24432,G24433,G24434,G24435,G24436,G24437,G24438,G24439,G24440,
       G24441,G24442,G24443,G24444,G24445,G24446,G24447,G24448,G24449,G24450,G24451,G24452,G24453,G24454,G24455,G24456,G24457,G24458,G24459,G24460,
       G24461,G24462,G24463,G24464,G24465,G24466,G24467,G24468,G24469,G24470,G24471,G24472,G24473,G24474,G24475,G24476,G24477,G24478,G24479,G24480,
       G24481,G24482,G24483,G24484,G24485,G24486,G24487,G24488,G24489,G24490,G24491,G24492,G24493,G24494,G24495,G24496,G24497,G24498,G24499,G24500,
       G24501,G24502,G24503,G24504,G24505,G24506,G24507,G24508,G24509,G24510,G24511,G24512,G24513,G24514,G24515,G24516,G24517,G24518,G24519,G24520,
       G24521,G24522,G24523,G24524,G24525,G24526,G24527,G24528,G24529,G24530,G24531,G24532,G24533,G24534,G24535,G24536,G24537,G24538,G24539,G24540,
       G24541,G24542,G24543,G24544,G24545,G24546,G24547,G24548,G24549,G24550,G24551,G24552,G24553,G24554,G24555,G24556,G24557,G24558,G24559,G24560,
       G24561,G24562,G24563,G24564,G24565,G24566,G24567,G24568,G24569,G24570,G24571,G24572,G24573,G24574,G24575,G24576,G24577,G24578,G24579,G24580,
       G24581,G24582,G24583,G24584,G24585,G24586,G24587,G24588,G24589,G24590,G24591,G24592,G24593,G24594,G24595,G24596,G24597,G24598,G24599,G24600,
       G24601,G24602,G24603,G24604,G24605,G24606,G24607,G24608,G24609,G24610,G24611,G24612,G24613,G24614,G24615,G24616,G24617,G24618,G24619,G24620,
       G24621,G24622,G24623,G24624,G24625,G24626,G24627,G24628,G24629,G24630,G24631,G24632,G24633,G24634,G24635,G24636,G24637,G24638,G24639,G24640,
       G24641,G24642,G24643,G24644,G24645,G24646,G24647,G24648,G24649,G24650,G24651,G24652,G24653,G24654,G24655,G24656,G24657,G24658,G24659,G24660,
       G24661,G24662,G24663,G24664,G24665,G24666,G24667,G24668,G24669,G24670,G24671,G24672,G24673,G24674,G24675,G24676,G24677,G24678,G24679,G24680,
       G24681,G24682,G24683,G24684,G24685,G24686,G24687,G24688,G24689,G24690,G24691,G24692,G24693,G24694,G24695,G24696,G24697,G24698,G24699,G24700,
       G24701,G24702,G24703,G24704,G24705,G24706,G24707,G24708,G24709,G24710,G24711,G24712,G24713,G24714,G24715,G24716,G24717,G24718,G24719,G24720,
       G24721,G24722,G24723,G24724,G24725,G24726,G24727,G24728,G24729,G24730,G24731,G24732,G24733,G24734,G24735,G24736,G24737,G24738,G24739,G24740,
       G24741,G24742,G24743,G24744,G24745,G24746,G24747,G24748,G24749,G24750,G24751,G24752,G24753,G24754,G24755,G24756,G24757,G24758,G24759,G24760,
       G24761,G24762,G24763,G24764,G24765,G24766,G24767,G24768,G24769,G24770,G24771,G24772,G24773,G24774,G24775,G24776,G24777,G24778,G24779,G24780,
       G24781,G24782,G24783,G24784,G24785,G24786,G24787,G24788,G24789,G24790,G24791,G24792,G24793,G24794,G24795,G24796,G24797,G24798,G24799,G24800,
       G24801,G24802,G24803,G24804,G24805,G24806,G24807,G24808,G24809,G24810,G24811,G24812,G24813,G24814,G24815,G24816,G24817,G24818,G24819,G24820,
       G24821,G24822,G24823,G24824,G24825,G24826,G24827,G24828,G24829,G24830,G24831,G24832,G24833,G24834,G24835,G24836,G24837,G24838,G24839,G24840,
       G24841,G24842,G24843,G24844,G24845,G24846,G24847,G24848,G24849,G24850,G24851,G24852,G24853,G24854,G24855,G24856,G24857,G24858,G24859,G24860,
       G24861,G24862,G24863,G24864,G24865,G24866,G24867,G24868,G24869,G24870,G24871,G24872,G24873,G24874,G24875,G24876,G24877,G24878,G24879,G24880,
       G24881,G24882,G24883,G24884,G24885,G24886,G24887,G24888,G24889,G24890,G24891,G24892,G24893,G24894,G24895,G24896,G24897,G24898,G24899,G24900,
       G24901,G24902,G24903,G24904,G24905,G24906,G24907,G24908,G24909,G24910,G24911,G24912,G24913,G24914,G24915,G24916,G24917,G24918,G24919,G24920,
       G24921,G24922,G24923,G24924,G24925,G24926,G24927,G24928,G24929,G24930,G24931,G24932,G24933,G24934,G24935,G24936,G24937,G24938,G24939,G24940,
       G24941,G24942,G24943,G24944,G24945,G24946,G24947,G24948,G24949,G24950,G24951,G24952,G24953,G24954,G24955,G24956,G24957,G24958,G24959,G24960,
       G24961,G24962,G24963,G24964,G24965,G24966,G24967,G24968,G24969,G24970,G24971,G24972,G24973,G24974,G24975,G24976,G24977,G24978,G24979,G24980,
       G24981,G24982,G24983,G24984,G24985,G24986,G24987,G24988,G24989,G24990,G24991,G24992,G24993,G24994,G24995,G24996,G24997,G24998,G24999,G25000,
       G25001,G25002,G25003,G25004,G25005,G25006,G25007,G25008,G25009,G25010,G25011,G25012,G25013,G25014,G25015,G25016,G25017,G25018,G25019,G25020,
       G25021,G25022,G25023,G25024,G25025,G25026,G25027,G25028,G25029,G25030,G25031,G25032,G25033,G25034,G25035,G25036,G25037,G25038,G25039,G25040,
       G25041,G25042,G25043,G25044,G25045,G25046,G25047,G25048,G25049,G25050,G25051,G25052,G25053,G25054,G25055,G25056,G25057,G25058,G25059,G25060,
       G25061,G25062,G25063,G25064,G25065,G25066,G25067,G25068,G25069,G25070,G25071,G25072,G25073,G25074,G25075,G25076,G25077,G25078,G25079,G25080,
       G25081,G25082,G25083,G25084,G25085,G25086,G25087,G25088,G25089,G25090,G25091,G25092,G25093,G25094,G25095,G25096,G25097,G25098,G25099,G25100,
       G25101,G25102,G25103,G25104,G25105,G25106,G25107,G25108,G25109,G25110,G25111,G25112,G25113,G25114,G25115,G25116,G25117,G25118,G25119,G25120,
       G25121,G25122,G25123,G25124,G25125,G25126,G25127,G25128,G25129,G25130,G25131,G25132,G25133,G25134,G25135,G25136,G25137,G25138,G25139,G25140,
       G25141,G25142,G25143,G25144,G25145,G25146,G25147,G25148,G25149,G25150,G25151,G25152,G25153,G25154,G25155,G25156,G25157,G25158,G25159,G25160,
       G25161,G25162,G25163,G25164,G25165,G25166,G25167,G25168,G25169,G25170,G25171,G25172,G25173,G25174,G25175,G25176,G25177,G25178,G25179,G25180,
       G25181,G25182,G25183,G25184,G25185,G25186,G25187,G25188,G25189,G25190,G25191,G25192,G25193,G25194,G25195,G25196,G25197,G25198,G25199,G25200,
       G25201,G25202,G25203,G25204,G25205,G25206,G25207,G25208,G25209,G25210,G25211,G25212,G25213,G25214,G25215,G25216,G25217,G25218,G25219,G25220,
       G25221,G25222,G25223,G25224,G25225,G25226,G25227,G25228,G25229,G25230,G25231,G25232,G25233,G25234,G25235,G25236,G25237,G25238,G25239,G25240,
       G25241,G25242,G25243,G25244,G25245,G25246,G25247,G25248,G25249,G25250,G25251,G25252,G25253,G25254,G25255,G25256,G25257,G25258,G25259,G25260,
       G25261,G25262,G25263,G25264,G25265,G25266,G25267,G25268,G25269,G25270,G25271,G25272,G25273,G25274,G25275,G25276,G25277,G25278,G25279,G25280,
       G25281,G25282,G25283,G25284,G25285,G25286,G25287,G25288,G25289,G25290,G25291,G25292,G25293,G25294,G25295,G25296,G25297,G25298,G25299,G25300,
       G25301,G25302,G25303,G25304,G25305,G25306,G25307,G25308,G25309,G25310,G25311,G25312,G25313,G25314,G25315,G25316,G25317,G25318,G25319,G25320,
       G25321,G25322,G25323,G25324,G25325,G25326,G25327,G25328,G25329,G25330,G25331,G25332,G25333,G25334,G25335,G25336,G25337,G25338,G25339,G25340,
       G25341,G25342,G25343,G25344,G25345,G25346,G25347,G25348,G25349,G25350,G25351,G25352,G25353,G25354,G25355,G25356,G25357,G25358,G25359,G25360,
       G25361,G25362,G25363,G25364,G25365,G25366,G25367,G25368,G25369,G25370,G25371,G25372,G25373,G25374,G25375,G25376,G25377,G25378,G25379,G25380,
       G25381,G25382,G25383,G25384,G25385,G25386,G25387,G25388,G25389,G25390,G25391,G25392,G25393,G25394,G25395,G25396,G25397,G25398,G25399,G25400,
       G25401,G25402,G25403,G25404,G25405,G25406,G25407,G25408,G25409,G25410,G25411,G25412,G25413,G25414,G25415,G25416,G25417,G25418,G25419,G25420,
       G25421,G25422,G25423,G25424,G25425,G25426,G25427,G25428,G25429,G25430,G25431,G25432,G25433,G25434,G25435,G25436,G25437,G25438,G25439,G25440,
       G25441,G25442,G25443,G25444,G25445,G25446,G25447,G25448,G25449,G25450,G25451,G25452,G25453,G25454,G25455,G25456,G25457,G25458,G25459,G25460,
       G25461,G25462,G25463,G25464,G25465,G25466,G25467,G25468,G25469,G25470,G25471,G25472,G25473,G25474,G25475,G25476,G25477,G25478,G25479,G25480,
       G25481,G25482,G25483,G25484,G25485,G25486,G25487,G25488,G25489,G25490,G25491,G25492,G25493,G25494,G25495,G25496,G25497,G25498,G25499,G25500,
       G25501,G25502,G25503,G25504,G25505,G25506,G25507,G25508,G25509,G25510,G25511,G25512,G25513,G25514,G25515,G25516,G25517,G25518,G25519,G25520,
       G25521,G25522,G25523,G25524,G25525,G25526,G25527,G25528,G25529,G25530,G25531,G25532,G25533,G25534,G25535,G25536,G25537,G25538,G25539,G25540,
       G25541,G25542,G25543,G25544,G25545,G25546,G25547,G25548,G25549,G25550,G25551,G25552,G25553,G25554,G25555,G25556,G25557,G25558,G25559,G25560,
       G25561,G25562,G25563,G25564,G25565,G25566,G25567,G25568,G25569,G25570,G25571,G25572,G25573,G25574,G25575,G25576,G25577,G25578,G25579,G25580,
       G25581,G25582,G25583,G25584,G25585,G25586,G25587,G25588,G25589,G25590,G25591,G25592,G25593,G25594,G25595,G25596,G25597,G25598,G25599,G25600,
       G25601,G25602,G25603,G25604,G25605,G25606,G25607,G25608,G25609,G25610,G25611,G25612,G25613,G25614,G25615,G25616,G25617,G25618,G25619,G25620,
       G25621,G25622,G25623,G25624,G25625,G25626,G25627,G25628,G25629,G25630,G25631,G25632,G25633,G25634,G25635,G25636,G25637,G25638,G25639,G25640,
       G25641,G25642,G25643,G25644,G25645,G25646,G25647,G25648,G25649,G25650,G25651,G25652,G25653,G25654,G25655,G25656,G25657,G25658,G25659,G25660,
       G25661,G25662,G25663,G25664,G25665,G25666,G25667,G25668,G25669,G25670,G25671,G25672,G25673,G25674,G25675,G25676,G25677,G25678,G25679,G25680,
       G25681,G25682,G25683,G25684,G25685,G25686,G25687,G25688,G25689,G25690,G25691,G25692,G25693,G25694,G25695,G25696,G25697,G25698,G25699,G25700,
       G25701,G25702,G25703,G25704,G25705,G25706,G25707,G25708,G25709,G25710,G25711,G25712,G25713,G25714,G25715,G25716,G25717,G25718,G25719,G25720,
       G25721,G25722,G25723,G25724,G25725,G25726,G25727,G25728,G25729,G25730,G25731,G25732,G25733,G25734,G25735,G25736,G25737,G25738,G25739,G25740,
       G25741,G25742,G25743,G25744,G25745,G25746,G25747,G25748,G25749,G25750,G25751,G25752,G25753,G25754,G25755,G25756,G25757,G25758,G25759,G25760,
       G25761,G25762,G25763,G25764,G25765,G25766,G25767,G25768,G25769,G25770,G25771,G25772,G25773,G25774,G25775,G25776,G25777,G25778,G25779,G25780,
       G25781,G25782,G25783,G25784,G25785,G25786,G25787,G25788,G25789,G25790,G25791,G25792,G25793,G25794,G25795,G25796,G25797,G25798,G25799,G25800,
       G25801,G25802,G25803,G25804,G25805,G25806,G25807,G25808,G25809,G25810,G25811,G25812,G25813,G25814,G25815,G25816,G25817,G25818,G25819,G25820,
       G25821,G25822,G25823,G25824,G25825,G25826,G25827,G25828,G25829,G25830,G25831,G25832,G25833,G25834,G25835,G25836,G25837,G25838,G25839,G25840,
       G25841,G25842,G25843,G25844,G25845,G25846,G25847,G25848,G25849,G25850,G25851,G25852,G25853,G25854,G25855,G25856,G25857,G25858,G25859,G25860,
       G25861,G25862,G25863,G25864,G25865,G25866,G25867,G25868,G25869,G25870,G25871,G25872,G25873,G25874,G25875,G25876,G25877,G25878,G25879,G25880,
       G25881,G25882,G25883,G25884,G25885,G25886,G25887,G25888,G25889,G25890,G25891,G25892,G25893,G25894,G25895,G25896,G25897,G25898,G25899,G25900,
       G25901,G25902,G25903,G25904,G25905,G25906,G25907,G25908,G25909,G25910,G25911,G25912,G25913,G25914,G25915,G25916,G25917,G25918,G25919,G25920,
       G25921,G25922,G25923,G25924,G25925,G25926,G25927,G25928,G25929,G25930,G25931,G25932,G25933,G25934,G25935,G25936,G25937,G25938,G25939,G25940,
       G25941,G25942,G25943,G25944,G25945,G25946,G25947,G25948,G25949,G25950,G25951,G25952,G25953,G25954,G25955,G25956,G25957,G25958,G25959,G25960,
       G25961,G25962,G25963,G25964,G25965,G25966,G25967,G25968,G25969,G25970,G25971,G25972,G25973,G25974,G25975,G25976,G25977,G25978,G25979,G25980,
       G25981,G25982,G25983,G25984,G25985,G25986,G25987,G25988,G25989,G25990,G25991,G25992,G25993,G25994,G25995,G25996,G25997,G25998,G25999,G26000,
       G26001,G26002,G26003,G26004,G26005,G26006,G26007,G26008,G26009,G26010,G26011,G26012,G26013,G26014,G26015,G26016,G26017,G26018,G26019,G26020,
       G26021,G26022,G26023,G26024,G26025,G26026,G26027,G26028,G26029,G26030,G26031,G26032,G26033,G26034,G26035,G26036,G26037,G26038,G26039,G26040,
       G26041,G26042,G26043,G26044,G26045,G26046,G26047,G26048,G26049,G26050,G26051,G26052,G26053,G26054,G26055,G26056,G26057,G26058,G26059,G26060,
       G26061,G26062,G26063,G26064,G26065,G26066,G26067,G26068,G26069,G26070,G26071,G26072,G26073,G26074,G26075,G26076,G26077,G26078,G26079,G26080,
       G26081,G26082,G26083,G26084,G26085,G26086,G26087,G26088,G26089,G26090,G26091,G26092,G26093,G26094,G26095,G26096,G26097,G26098,G26099,G26100,
       G26101,G26102,G26103,G26104,G26105,G26106,G26107,G26108,G26109,G26110,G26111,G26112,G26113,G26114,G26115,G26116,G26117,G26118,G26119,G26120,
       G26121,G26122,G26123,G26124,G26125,G26126,G26127,G26128,G26129,G26130,G26131,G26132,G26133,G26134,G26135,G26136,G26137,G26138,G26139,G26140,
       G26141,G26142,G26143,G26144,G26145,G26146,G26147,G26148,G26149,G26150,G26151,G26152,G26153,G26154,G26155,G26156,G26157,G26158,G26159,G26160,
       G26161,G26162,G26163,G26164,G26165,G26166,G26167,G26168,G26169,G26170,G26171,G26172,G26173,G26174,G26175,G26176,G26177,G26178,G26179,G26180,
       G26181,G26182,G26183,G26184,G26185,G26186,G26187,G26188,G26189,G26190,G26191,G26192,G26193,G26194,G26195,G26196,G26197,G26198,G26199,G26200,
       G26201,G26202,G26203,G26204,G26205,G26206,G26207,G26208,G26209,G26210,G26211,G26212,G26213,G26214,G26215,G26216,G26217,G26218,G26219,G26220,
       G26221,G26222,G26223,G26224,G26225,G26226,G26227,G26228,G26229,G26230,G26231,G26232,G26233,G26234,G26235,G26236,G26237,G26238,G26239,G26240,
       G26241,G26242,G26243,G26244,G26245,G26246,G26247,G26248,G26249,G26250,G26251,G26252,G26253,G26254,G26255,G26256,G26257,G26258,G26259,G26260,
       G26261,G26262,G26263,G26264,G26265,G26266,G26267,G26268,G26269,G26270,G26271,G26272,G26273,G26274,G26275,G26276,G26277,G26278,G26279,G26280,
       G26281,G26282,G26283,G26284,G26285,G26286,G26287,G26288,G26289,G26290,G26291,G26292,G26293,G26294,G26295,G26296,G26297,G26298,G26299,G26300,
       G26301,G26302,G26303,G26304,G26305,G26306,G26307,G26308,G26309,G26310,G26311,G26312,G26313,G26314,G26315,G26316,G26317,G26318,G26319,G26320,
       G26321,G26322,G26323,G26324,G26325,G26326,G26327,G26328,G26329,G26330,G26331,G26332,G26333,G26334,G26335,G26336,G26337,G26338,G26339,G26340,
       G26341,G26342,G26343,G26344,G26345,G26346,G26347,G26348,G26349,G26350,G26351,G26352,G26353,G26354,G26355,G26356,G26357,G26358,G26359,G26360,
       G26361,G26362,G26363,G26364,G26365,G26366,G26367,G26368,G26369,G26370,G26371,G26372,G26373,G26374,G26375,G26376,G26377,G26378,G26379,G26380,
       G26381,G26382,G26383,G26384,G26385,G26386,G26387,G26388,G26389,G26390,G26391,G26392,G26393,G26394,G26395,G26396,G26397,G26398,G26399,G26400,
       G26401,G26402,G26403,G26404,G26405,G26406,G26407,G26408,G26409,G26410,G26411,G26412,G26413,G26414,G26415,G26416,G26417,G26418,G26419,G26420,
       G26421,G26422,G26423,G26424,G26425,G26426,G26427,G26428,G26429,G26430,G26431,G26432,G26433,G26434,G26435,G26436,G26437,G26438,G26439,G26440,
       G26441,G26442,G26443,G26444,G26445,G26446,G26447,G26448,G26449,G26450,G26451,G26452,G26453,G26454,G26455,G26456,G26457,G26458,G26459,G26460,
       G26461,G26462,G26463,G26464,G26465,G26466,G26467,G26468,G26469,G26470,G26471,G26472,G26473,G26474,G26475,G26476,G26477,G26478,G26479,G26480,
       G26481,G26482,G26483,G26484,G26485,G26486,G26487,G26488,G26489,G26490,G26491,G26492,G26493,G26494,G26495,G26496,G26497,G26498,G26499,G26500,
       G26501,G26502,G26503,G26504,G26505,G26506,G26507,G26508,G26509,G26510,G26511,G26512,G26513,G26514,G26515,G26516,G26517,G26518,G26519,G26520,
       G26521,G26522,G26523,G26524,G26525,G26526,G26527,G26528,G26529,G26530,G26531,G26532,G26533,G26534,G26535,G26536,G26537,G26538,G26539,G26540,
       G26541,G26542,G26543,G26544,G26545,G26546,G26547,G26548,G26549,G26550,G26551,G26552,G26553,G26554,G26555,G26556,G26557,G26558,G26559,G26560,
       G26561,G26562,G26563,G26564,G26565,G26566,G26567,G26568,G26569,G26570,G26571,G26572,G26573,G26574,G26575,G26576,G26577,G26578,G26579,G26580,
       G26581,G26582,G26583,G26584,G26585,G26586,G26587,G26588,G26589,G26590,G26591,G26592,G26593,G26594,G26595,G26596,G26597,G26598,G26599,G26600,
       G26601,G26602,G26603,G26604,G26605,G26606,G26607,G26608,G26609,G26610,G26611,G26612,G26613,G26614,G26615,G26616,G26617,G26618,G26619,G26620,
       G26621,G26622,G26623,G26624,G26625,G26626,G26627,G26628,G26629,G26630,G26631,G26632,G26633,G26634,G26635,G26636,G26637,G26638,G26639,G26640,
       G26641,G26642,G26643,G26644,G26645,G26646,G26647,G26648,G26649,G26650,G26651,G26652,G26653,G26654,G26655,G26656,G26657,G26658,G26659,G26660,
       G26661,G26662,G26663,G26664,G26665,G26666,G26667,G26668,G26669,G26670,G26671,G26672,G26673,G26674,G26675,G26676,G26677,G26678,G26679,G26680,
       G26681,G26682,G26683,G26684,G26685,G26686,G26687,G26688,G26689,G26690,G26691,G26692,G26693,G26694,G26695,G26696,G26697,G26698,G26699,G26700,
       G26701,G26702,G26703,G26704,G26705,G26706,G26707,G26708,G26709,G26710,G26711,G26712,G26713,G26714,G26715,G26716,G26717,G26718,G26719,G26720,
       G26721,G26722,G26723,G26724,G26725,G26726,G26727,G26728,G26729,G26730,G26731,G26732,G26733,G26734,G26735,G26736,G26737,G26738,G26739,G26740,
       G26741,G26742,G26743,G26744,G26745,G26746,G26747,G26748,G26749,G26750,G26751,G26752,G26753,G26754,G26755,G26756,G26757,G26758,G26759,G26760,
       G26761,G26762,G26763,G26764,G26765,G26766,G26767,G26768,G26769,G26770,G26771,G26772,G26773,G26774,G26775,G26776,G26777,G26778,G26779,G26780,
       G26781,G26782,G26783,G26784,G26785,G26786,G26787,G26788,G26789,G26790,G26791,G26792,G26793,G26794,G26795,G26796,G26797,G26798,G26799,G26800,
       G26801,G26802,G26803,G26804,G26805,G26806,G26807,G26808,G26809,G26810,G26811,G26812,G26813,G26814,G26815,G26816,G26817,G26818,G26819,G26820,
       G26821,G26822,G26823,G26824,G26825,G26826,G26827,G26828,G26829,G26830,G26831,G26832,G26833,G26834,G26835,G26836,G26837,G26838,G26839,G26840,
       G26841,G26842,G26843,G26844,G26845,G26846,G26847,G26848,G26849,G26850,G26851,G26852,G26853,G26854,G26855,G26856,G26857,G26858,G26859,G26860,
       G26861,G26862,G26863,G26864,G26865,G26866,G26867,G26868,G26869,G26870,G26871,G26872,G26873,G26874,G26875,G26876,G26877,G26878,G26879,G26880,
       G26881,G26882,G26883,G26884,G26885,G26886,G26887,G26888,G26889,G26890,G26891,G26892,G26893,G26894,G26895,G26896,G26897,G26898,G26899,G26900,
       G26901,G26902,G26903,G26904,G26905,G26906,G26907,G26908,G26909,G26910,G26911,G26912,G26913,G26914,G26915,G26916,G26917,G26918,G26919,G26920,
       G26921,G26922,G26923,G26924,G26925,G26926,G26927,G26928,G26929,G26930,G26931,G26932,G26933,G26934,G26935,G26936,G26937,G26938,G26939,G26940,
       G26941,G26942,G26943,G26944,G26945,G26946,G26947,G26948,G26949,G26950,G26951,G26952,G26953,G26954,G26955,G26956,G26957,G26958,G26959,G26960,
       G26961,G26962,G26963,G26964,G26965,G26966,G26967,G26968,G26969,G26970,G26971,G26972,G26973,G26974,G26975,G26976,G26977,G26978,G26979,G26980,
       G26981,G26982,G26983,G26984,G26985,G26986,G26987,G26988,G26989,G26990,G26991,G26992,G26993,G26994,G26995,G26996,G26997,G26998,G26999,G27000,
       G27001,G27002,G27003,G27004,G27005,G27006,G27007,G27008,G27009,G27010,G27011,G27012,G27013,G27014,G27015,G27016,G27017,G27018,G27019,G27020,
       G27021,G27022,G27023,G27024,G27025,G27026,G27027,G27028,G27029,G27030,G27031,G27032,G27033,G27034,G27035,G27036,G27037,G27038,G27039,G27040,
       G27041,G27042,G27043,G27044,G27045,G27046,G27047,G27048,G27049,G27050,G27051,G27052,G27053,G27054,G27055,G27056,G27057,G27058,G27059,G27060,
       G27061,G27062,G27063,G27064,G27065,G27066,G27067,G27068,G27069,G27070,G27071,G27072,G27073,G27074,G27075,G27076,G27077,G27078,G27079,G27080,
       G27081,G27082,G27083,G27084,G27085,G27086,G27087,G27088,G27089,G27090,G27091,G27092,G27093,G27094,G27095,G27096,G27097,G27098,G27099,G27100,
       G27101,G27102,G27103,G27104,G27105,G27106,G27107,G27108,G27109,G27110,G27111,G27112,G27113,G27114,G27115,G27116,G27117,G27118,G27119,G27120,
       G27121,G27122,G27123,G27124,G27125,G27126,G27127,G27128,G27129,G27130,G27131,G27132,G27133,G27134,G27135,G27136,G27137,G27138,G27139,G27140,
       G27141,G27142,G27143,G27144,G27145,G27146,G27147,G27148,G27149,G27150,G27151,G27152,G27153,G27154,G27155,G27156,G27157,G27158,G27159,G27160,
       G27161,G27162,G27163,G27164,G27165,G27166,G27167,G27168,G27169,G27170,G27171,G27172,G27173,G27174,G27175,G27176,G27177,G27178,G27179,G27180,
       G27181,G27182,G27183,G27184,G27185,G27186,G27187,G27188,G27189,G27190,G27191,G27192,G27193,G27194,G27195,G27196,G27197,G27198,G27199,G27200,
       G27201,G27202,G27203,G27204,G27205,G27206,G27207,G27208,G27209,G27210,G27211,G27212,G27213,G27214,G27215,G27216,G27217,G27218,G27219,G27220,
       G27221,G27222,G27223,G27224,G27225,G27226,G27227,G27228,G27229,G27230,G27231,G27232,G27233,G27234,G27235,G27236,G27237,G27238,G27239,G27240,
       G27241,G27242,G27243,G27244,G27245,G27246,G27247,G27248,G27249,G27250,G27251,G27252,G27253,G27254,G27255,G27256,G27257,G27258,G27259,G27260,
       G27261,G27262,G27263,G27264,G27265,G27266,G27267,G27268,G27269,G27270,G27271,G27272,G27273,G27274,G27275,G27276,G27277,G27278,G27279,G27280,
       G27281,G27282,G27283,G27284,G27285,G27286,G27287,G27288,G27289,G27290,G27291,G27292,G27293,G27294,G27295,G27296,G27297,G27298,G27299,G27300,
       G27301,G27302,G27303,G27304,G27305,G27306,G27307,G27308,G27309,G27310,G27311,G27312,G27313,G27314,G27315,G27316,G27317,G27318,G27319,G27320,
       G27321,G27322,G27323,G27324,G27325,G27326,G27327,G27328,G27329,G27330,G27331,G27332,G27333,G27334,G27335,G27336,G27337,G27338,G27339,G27340,
       G27341,G27342,G27343,G27344,G27345,G27346,G27347,G27348,G27349,G27350,G27351,G27352,G27353,G27354,G27355,G27356,G27357,G27358,G27359,G27360,
       G27361,G27362,G27363,G27364,G27365,G27366,G27367,G27368,G27369,G27370,G27371,G27372,G27373,G27374,G27375,G27376,G27377,G27378,G27379,G27380,
       G27381,G27382,G27383,G27384,G27385,G27386,G27387,G27388,G27389,G27390,G27391,G27392,G27393,G27394,G27395,G27396,G27397,G27398,G27399,G27400,
       G27401,G27402,G27403,G27404,G27405,G27406,G27407,G27408,G27409,G27410,G27411,G27412,G27413,G27414,G27415,G27416,G27417,G27418,G27419,G27420,
       G27421,G27422,G27423,G27424,G27425,G27426,G27427,G27428,G27429,G27430,G27431,G27432,G27433,G27434,G27435,G27436,G27437,G27438,G27439,G27440,
       G27441,G27442,G27443,G27444,G27445,G27446,G27447,G27448,G27449,G27450,G27451,G27452,G27453,G27454,G27455,G27456,G27457,G27458,G27459,G27460,
       G27461,G27462,G27463,G27464,G27465,G27466,G27467,G27468,G27469,G27470,G27471,G27472,G27473,G27474,G27475,G27476,G27477,G27478,G27479,G27480,
       G27481,G27482,G27483,G27484,G27485,G27486,G27487,G27488,G27489,G27490,G27491,G27492,G27493,G27494,G27495,G27496,G27497,G27498,G27499,G27500,
       G27501,G27502,G27503,G27504,G27505,G27506,G27507,G27508,G27509,G27510,G27511,G27512,G27513,G27514,G27515,G27516,G27517,G27518,G27519,G27520,
       G27521,G27522,G27523,G27524,G27525,G27526,G27527,G27528,G27529,G27530,G27531,G27532,G27533,G27534,G27535,G27536,G27537,G27538,G27539,G27540,
       G27541,G27542,G27543,G27544,G27545,G27546,G27547,G27548,G27549,G27550,G27551,G27552,G27553,G27554,G27555,G27556,G27557,G27558,G27559,G27560,
       G27561,G27562,G27563,G27564,G27565,G27566,G27567,G27568,G27569,G27570,G27571,G27572,G27573,G27574,G27575,G27576,G27577,G27578,G27579,G27580,
       G27581,G27582,G27583,G27584,G27585,G27586,G27587,G27588,G27589,G27590,G27591,G27592,G27593,G27594,G27595,G27596,G27597,G27598,G27599,G27600,
       G27601,G27602,G27603,G27604,G27605,G27606,G27607,G27608,G27609,G27610,G27611,G27612,G27613,G27614,G27615,G27616,G27617,G27618,G27619,G27620,
       G27621,G27622,G27623,G27624,G27625,G27626,G27627,G27628,G27629,G27630,G27631,G27632,G27633,G27634,G27635,G27636,G27637,G27638,G27639,G27640,
       G27641,G27642,G27643,G27644,G27645,G27646,G27647,G27648,G27649,G27650,G27651,G27652,G27653,G27654,G27655,G27656,G27657,G27658,G27659,G27660,
       G27661,G27662,G27663,G27664,G27665,G27666,G27667,G27668,G27669,G27670,G27671,G27672,G27673,G27674,G27675,G27676,G27677,G27678,G27679,G27680,
       G27681,G27682,G27683,G27684,G27685,G27686,G27687,G27688,G27689,G27690,G27691,G27692,G27693,G27694,G27695,G27696,G27697,G27698,G27699,G27700,
       G27701,G27702,G27703,G27704,G27705,G27706,G27707,G27708,G27709,G27710,G27711,G27712,G27713,G27714,G27715,G27716,G27717,G27718,G27719,G27720,
       G27721,G27722,G27723,G27724,G27725,G27726,G27727,G27728,G27729,G27730,G27731,G27732,G27733,G27734,G27735,G27736,G27737,G27738,G27739,G27740,
       G27741,G27742,G27743,G27744,G27745,G27746,G27747,G27748,G27749,G27750,G27751,G27752,G27753,G27754,G27755,G27756,G27757,G27758,G27759,G27760,
       G27761,G27762,G27763,G27764,G27765,G27766,G27767,G27768,G27769,G27770,G27771,G27772,G27773,G27774,G27775,G27776,G27777,G27778,G27779,G27780,
       G27781,G27782,G27783,G27784,G27785,G27786,G27787,G27788,G27789,G27790,G27791,G27792,G27793,G27794,G27795,G27796,G27797,G27798,G27799,G27800,
       G27801,G27802,G27803,G27804,G27805,G27806,G27807,G27808,G27809,G27810,G27811,G27812,G27813,G27814,G27815,G27816,G27817,G27818,G27819,G27820,
       G27821,G27822,G27823,G27824,G27825,G27826,G27827,G27828,G27829,G27830,G27831,G27832,G27833,G27834,G27835,G27836,G27837,G27838,G27839,G27840,
       G27841,G27842,G27843,G27844,G27845,G27846,G27847,G27848,G27849,G27850,G27851,G27852,G27853,G27854,G27855,G27856,G27857,G27858,G27859,G27860,
       G27861,G27862,G27863,G27864,G27865,G27866,G27867,G27868,G27869,G27870,G27871,G27872,G27873,G27874,G27875,G27876,G27877,G27878,G27879,G27880,
       G27881,G27882,G27883,G27884,G27885,G27886,G27887,G27888,G27889,G27890,G27891,G27892,G27893,G27894,G27895,G27896,G27897,G27898,G27899,G27900,
       G27901,G27902,G27903,G27904,G27905,G27906,G27907,G27908,G27909,G27910,G27911,G27912,G27913,G27914,G27915,G27916,G27917,G27918,G27919,G27920,
       G27921,G27922,G27923,G27924,G27925,G27926,G27927,G27928,G27929,G27930,G27931,G27932,G27933,G27934,G27935,G27936,G27937,G27938,G27939,G27940,
       G27941,G27942,G27943,G27944,G27945,G27946,G27947,G27948,G27949,G27950,G27951,G27952,G27953,G27954,G27955,G27956,G27957,G27958,G27959,G27960,
       G27961,G27962,G27963,G27964,G27965,G27966,G27967,G27968,G27969,G27970,G27971,G27972,G27973,G27974,G27975,G27976,G27977,G27978,G27979,G27980,
       G27981,G27982,G27983,G27984,G27985,G27986,G27987,G27988,G27989,G27990,G27991,G27992,G27993,G27994,G27995,G27996,G27997,G27998,G27999,G28000,
       G28001,G28002,G28003,G28004,G28005,G28006,G28007,G28008,G28009,G28010,G28011,G28012,G28013,G28014,G28015,G28016,G28017,G28018,G28019,G28020,
       G28021,G28022,G28023,G28024,G28025,G28026,G28027,G28028,G28029,G28030,G28031,G28032,G28033,G28034,G28035,G28036,G28037,G28038,G28039,G28040,
       G28041,G28042,G28043,G28044,G28045,G28046,G28047,G28048,G28049,G28050,G28051,G28052,G28053,G28054,G28055,G28056,G28057,G28058,G28059,G28060,
       G28061,G28062,G28063,G28064,G28065,G28066,G28067,G28068,G28069,G28070,G28071,G28072,G28073,G28074,G28075,G28076,G28077,G28078,G28079,G28080,
       G28081,G28082,G28083,G28084,G28085,G28086,G28087,G28088,G28089,G28090,G28091,G28092,G28093,G28094,G28095,G28096,G28097,G28098,G28099,G28100,
       G28101,G28102,G28103,G28104,G28105,G28106,G28107,G28108,G28109,G28110,G28111,G28112,G28113,G28114,G28115,G28116,G28117,G28118,G28119,G28120,
       G28121,G28122,G28123,G28124,G28125,G28126,G28127,G28128,G28129,G28130,G28131,G28132,G28133,G28134,G28135,G28136,G28137,G28138,G28139,G28140,
       G28141,G28142,G28143,G28144,G28145,G28146,G28147,G28148,G28149,G28150,G28151,G28152,G28153,G28154,G28155,G28156,G28157,G28158,G28159,G28160,
       G28161,G28162,G28163,G28164,G28165,G28166,G28167,G28168,G28169,G28170,G28171,G28172,G28173,G28174,G28175,G28176,G28177,G28178,G28179,G28180,
       G28181,G28182,G28183,G28184,G28185,G28186,G28187,G28188,G28189,G28190,G28191,G28192,G28193,G28194,G28195,G28196,G28197,G28198,G28199,G28200,
       G28201,G28202,G28203,G28204,G28205,G28206,G28207,G28208,G28209,G28210,G28211,G28212,G28213,G28214,G28215,G28216,G28217,G28218,G28219,G28220,
       G28221,G28222,G28223,G28224,G28225,G28226,G28227,G28228,G28229,G28230,G28231,G28232,G28233,G28234,G28235,G28236,G28237,G28238,G28239,G28240,
       G28241,G28242,G28243,G28244,G28245,G28246,G28247,G28248,G28249,G28250,G28251,G28252,G28253,G28254,G28255,G28256,G28257,G28258,G28259,G28260,
       G28261,G28262,G28263,G28264,G28265,G28266,G28267,G28268,G28269,G28270,G28271,G28272,G28273,G28274,G28275,G28276,G28277,G28278,G28279,G28280,
       G28281,G28282,G28283,G28284,G28285,G28286,G28287,G28288,G28289,G28290,G28291,G28292,G28293,G28294,G28295,G28296,G28297,G28298,G28299,G28300,
       G28301,G28302,G28303,G28304,G28305,G28306,G28307,G28308,G28309,G28310,G28311,G28312,G28313,G28314,G28315,G28316,G28317,G28318,G28319,G28320,
       G28321,G28322,G28323,G28324,G28325,G28326,G28327,G28328,G28329,G28330,G28331,G28332,G28333,G28334,G28335,G28336,G28337,G28338,G28339,G28340,
       G28341,G28342,G28343,G28344,G28345,G28346,G28347,G28348,G28349,G28350,G28351,G28352,G28353,G28354,G28355,G28356,G28357,G28358,G28359,G28360,
       G28361,G28362,G28363,G28364,G28365,G28366,G28367,G28368,G28369,G28370,G28371,G28372,G28373,G28374,G28375,G28376,G28377,G28378,G28379,G28380,
       G28381,G28382,G28383,G28384,G28385,G28386,G28387,G28388,G28389,G28390,G28391,G28392,G28393,G28394,G28395,G28396,G28397,G28398,G28399,G28400,
       G28401,G28402,G28403,G28404,G28405,G28406,G28407,G28408,G28409,G28410,G28411,G28412,G28413,G28414,G28415,G28416,G28417,G28418,G28419,G28420,
       G28421,G28422,G28423,G28424,G28425,G28426,G28427,G28428,G28429,G28430,G28431,G28432,G28433,G28434,G28435,G28436,G28437,G28438,G28439,G28440,
       G28441,G28442,G28443,G28444,G28445,G28446,G28447,G28448,G28449,G28450,G28451,G28452,G28453,G28454,G28455,G28456,G28457,G28458,G28459,G28460,
       G28461,G28462,G28463,G28464,G28465,G28466,G28467,G28468,G28469,G28470,G28471,G28472,G28473,G28474,G28475,G28476,G28477,G28478,G28479,G28480,
       G28481,G28482,G28483,G28484,G28485,G28486,G28487,G28488,G28489,G28490,G28491,G28492,G28493,G28494,G28495,G28496,G28497,G28498,G28499,G28500,
       G28501,G28502,G28503,G28504,G28505,G28506,G28507,G28508,G28509,G28510,G28511,G28512,G28513,G28514,G28515,G28516,G28517,G28518,G28519,G28520,
       G28521,G28522,G28523,G28524,G28525,G28526,G28527,G28528,G28529,G28530,G28531,G28532,G28533,G28534,G28535,G28536,G28537,G28538,G28539,G28540,
       G28541,G28542,G28543,G28544,G28545,G28546,G28547,G28548,G28549,G28550,G28551,G28552,G28553,G28554,G28555,G28556,G28557,G28558,G28559,G28560,
       G28561,G28562,G28563,G28564,G28565,G28566,G28567,G28568,G28569,G28570,G28571,G28572,G28573,G28574,G28575,G28576,G28577,G28578,G28579,G28580,
       G28581,G28582,G28583,G28584,G28585,G28586,G28587,G28588,G28589,G28590,G28591,G28592,G28593,G28594,G28595,G28596,G28597,G28598,G28599,G28600,
       G28601,G28602,G28603,G28604,G28605,G28606,G28607,G28608,G28609,G28610,G28611,G28612,G28613,G28614,G28615,G28616,G28617,G28618,G28619,G28620,
       G28621,G28622,G28623,G28624,G28625,G28626,G28627,G28628,G28629,G28630,G28631,G28632,G28633,G28634,G28635,G28636,G28637,G28638,G28639,G28640,
       G28641,G28642,G28643,G28644,G28645,G28646,G28647,G28648,G28649,G28650,G28651,G28652,G28653,G28654,G28655,G28656,G28657,G28658,G28659,G28660,
       G28661,G28662,G28663,G28664,G28665,G28666,G28667,G28668,G28669,G28670,G28671,G28672,G28673,G28674,G28675,G28676,G28677,G28678,G28679,G28680,
       G28681,G28682,G28683,G28684,G28685,G28686,G28687,G28688,G28689,G28690,G28691,G28692,G28693,G28694,G28695,G28696,G28697,G28698,G28699,G28700,
       G28701,G28702,G28703,G28704,G28705,G28706,G28707,G28708,G28709,G28710,G28711,G28712,G28713,G28714,G28715,G28716,G28717,G28718,G28719,G28720,
       G28721,G28722,G28723,G28724,G28725,G28726,G28727,G28728,G28729,G28730,G28731,G28732,G28733,G28734,G28735,G28736,G28737,G28738,G28739,G28740,
       G28741,G28742,G28743,G28744,G28745,G28746,G28747,G28748,G28749,G28750,G28751,G28752,G28753,G28754,G28755,G28756,G28757,G28758,G28759,G28760,
       G28761,G28762,G28763,G28764,G28765,G28766,G28767,G28768,G28769,G28770,G28771,G28772,G28773,G28774,G28775,G28776,G28777,G28778,G28779,G28780,
       G28781,G28782,G28783,G28784,G28785,G28786,G28787,G28788,G28789,G28790,G28791,G28792,G28793,G28794,G28795,G28796,G28797,G28798,G28799,G28800,
       G28801,G28802,G28803,G28804,G28805,G28806,G28807,G28808,G28809,G28810,G28811,G28812,G28813,G28814,G28815,G28816,G28817,G28818,G28819,G28820,
       G28821,G28822,G28823,G28824,G28825,G28826,G28827,G28828,G28829,G28830,G28831,G28832,G28833,G28834,G28835,G28836,G28837,G28838,G28839,G28840,
       G28841,G28842,G28843,G28844,G28845,G28846,G28847,G28848,G28849,G28850,G28851,G28852,G28853,G28854,G28855,G28856,G28857,G28858,G28859,G28860,
       G28861,G28862,G28863,G28864,G28865,G28866,G28867,G28868,G28869,G28870,G28871,G28872,G28873,G28874,G28875,G28876,G28877,G28878,G28879,G28880,
       G28881,G28882,G28883,G28884,G28885,G28886,G28887,G28888,G28889,G28890,G28891,G28892,G28893,G28894,G28895,G28896,G28897,G28898,G28899,G28900,
       G28901,G28902,G28903,G28904,G28905,G28906,G28907,G28908,G28909,G28910,G28911,G28912,G28913,G28914,G28915,G28916,G28917,G28918,G28919,G28920,
       G28921,G28922,G28923,G28924,G28925,G28926,G28927,G28928,G28929,G28930,G28931,G28932,G28933,G28934,G28935,G28936,G28937,G28938,G28939,G28940,
       G28941,G28942,G28943,G28944,G28945,G28946,G28947,G28948,G28949,G28950,G28951,G28952,G28953,G28954,G28955,G28956,G28957,G28958,G28959,G28960,
       G28961,G28962,G28963,G28964,G28965,G28966,G28967,G28968,G28969,G28970,G28971,G28972,G28973,G28974,G28975,G28976,G28977,G28978,G28979,G28980,
       G28981,G28982,G28983,G28984,G28985,G28986,G28987,G28988,G28989,G28990,G28991,G28992,G28993,G28994,G28995,G28996,G28997,G28998,G28999,G29000,
       G29001,G29002,G29003,G29004,G29005,G29006,G29007,G29008,G29009,G29010,G29011,G29012,G29013,G29014,G29015,G29016,G29017,G29018,G29019,G29020,
       G29021,G29022,G29023,G29024,G29025,G29026,G29027,G29028,G29029,G29030,G29031,G29032,G29033,G29034,G29035,G29036,G29037,G29038,G29039,G29040,
       G29041,G29042,G29043,G29044,G29045,G29046,G29047,G29048,G29049,G29050,G29051,G29052,G29053,G29054,G29055,G29056,G29057,G29058,G29059,G29060,
       G29061,G29062,G29063,G29064,G29065,G29066,G29067,G29068,G29069,G29070,G29071,G29072,G29073,G29074,G29075,G29076,G29077,G29078,G29079,G29080,
       G29081,G29082,G29083,G29084,G29085,G29086,G29087,G29088,G29089,G29090,G29091,G29092,G29093,G29094,G29095,G29096,G29097,G29098,G29099,G29100,
       G29101,G29102,G29103,G29104,G29105,G29106,G29107,G29108,G29109,G29110,G29111,G29112,G29113,G29114,G29115,G29116,G29117,G29118,G29119,G29120,
       G29121,G29122,G29123,G29124,G29125,G29126,G29127,G29128,G29129,G29130,G29131,G29132,G29133,G29134,G29135,G29136,G29137,G29138,G29139,G29140,
       G29141,G29142,G29143,G29144,G29145,G29146,G29147,G29148,G29149,G29150,G29151,G29152,G29153,G29154,G29155,G29156,G29157,G29158,G29159,G29160,
       G29161,G29162,G29163,G29164,G29165,G29166,G29167,G29168,G29169,G29170,G29171,G29172,G29173,G29174,G29175,G29176,G29177,G29178,G29179,G29180,
       G29181,G29182,G29183,G29184,G29185,G29186,G29187,G29188,G29189,G29190,G29191,G29192,G29193,G29194,G29195,G29196,G29197,G29198,G29199,G29200,
       G29201,G29202,G29203,G29204,G29205,G29206,G29207,G29208,G29209,G29210,G29211,G29212,G29213,G29214,G29215,G29216,G29217,G29218,G29219,G29220,
       G29221,G29222,G29223,G29224,G29225,G29226,G29227,G29228,G29229,G29230,G29231,G29232,G29233,G29234,G29235,G29236,G29237,G29238,G29239,G29240,
       G29241,G29242,G29243,G29244,G29245,G29246,G29247,G29248,G29249,G29250,G29251,G29252,G29253,G29254,G29255,G29256,G29257,G29258,G29259,G29260,
       G29261,G29262,G29263,G29264,G29265,G29266,G29267,G29268,G29269,G29270,G29271,G29272,G29273,G29274,G29275,G29276,G29277,G29278,G29279,G29280,
       G29281,G29282,G29283,G29284,G29285,G29286,G29287,G29288,G29289,G29290,G29291,G29292,G29293,G29294,G29295,G29296,G29297,G29298,G29299,G29300,
       G29301,G29302,G29303,G29304,G29305,G29306,G29307,G29308,G29309,G29310,G29311,G29312,G29313,G29314,G29315,G29316,G29317,G29318,G29319,G29320,
       G29321,G29322,G29323,G29324,G29325,G29326,G29327,G29328,G29329,G29330,G29331,G29332,G29333,G29334,G29335,G29336,G29337,G29338,G29339,G29340,
       G29341,G29342,G29343,G29344,G29345,G29346,G29347,G29348,G29349,G29350,G29351,G29352,G29353,G29354,G29355,G29356,G29357,G29358,G29359,G29360,
       G29361,G29362,G29363,G29364,G29365,G29366,G29367,G29368,G29369,G29370,G29371,G29372,G29373,G29374,G29375,G29376,G29377,G29378,G29379,G29380,
       G29381,G29382,G29383,G29384,G29385,G29386,G29387,G29388,G29389,G29390,G29391,G29392,G29393,G29394,G29395,G29396,G29397,G29398,G29399,G29400,
       G29401,G29402,G29403,G29404,G29405,G29406,G29407,G29408,G29409,G29410,G29411,G29412,G29413,G29414,G29415,G29416,G29417,G29418,G29419,G29420,
       G29421,G29422,G29423,G29424,G29425,G29426,G29427,G29428,G29429,G29430,G29431,G29432,G29433,G29434,G29435,G29436,G29437,G29438,G29439,G29440,
       G29441,G29442,G29443,G29444,G29445,G29446,G29447,G29448,G29449,G29450,G29451,G29452,G29453,G29454,G29455,G29456,G29457,G29458,G29459,G29460,
       G29461,G29462,G29463,G29464,G29465,G29466,G29467,G29468,G29469,G29470,G29471,G29472,G29473,G29474,G29475,G29476,G29477,G29478,G29479,G29480,
       G29481,G29482,G29483,G29484,G29485,G29486,G29487,G29488,G29489,G29490,G29491,G29492,G29493,G29494,G29495,G29496,G29497,G29498,G29499,G29500,
       G29501,G29502,G29503,G29504,G29505,G29506,G29507,G29508,G29509,G29510,G29511,G29512,G29513,G29514,G29515,G29516,G29517,G29518,G29519,G29520,
       G29521,G29522,G29523,G29524,G29525,G29526,G29527,G29528,G29529,G29530,G29531,G29532,G29533,G29534,G29535,G29536,G29537,G29538,G29539,G29540,
       G29541,G29542,G29543,G29544,G29545,G29546,G29547,G29548,G29549,G29550,G29551,G29552,G29553,G29554,G29555,G29556,G29557,G29558,G29559,G29560,
       G29561,G29562,G29563,G29564,G29565,G29566,G29567,G29568,G29569,G29570,G29571,G29572,G29573,G29574,G29575,G29576,G29577,G29578,G29579,G29580,
       G29581,G29582,G29583,G29584,G29585,G29586,G29587,G29588,G29589,G29590,G29591,G29592,G29593,G29594,G29595,G29596,G29597,G29598,G29599,G29600,
       G29601,G29602,G29603,G29604,G29605,G29606,G29607,G29608,G29609,G29610,G29611,G29612,G29613,G29614,G29615,G29616,G29617,G29618,G29619,G29620,
       G29621,G29622,G29623,G29624,G29625,G29626,G29627,G29628,G29629,G29630,G29631,G29632,G29633,G29634,G29635,G29636,G29637,G29638,G29639,G29640,
       G29641,G29642,G29643,G29644,G29645,G29646,G29647,G29648,G29649,G29650,G29651,G29652,G29653,G29654,G29655,G29656,G29657,G29658,G29659,G29660,
       G29661,G29662,G29663,G29664,G29665,G29666,G29667,G29668,G29669,G29670,G29671,G29672,G29673,G29674,G29675,G29676,G29677,G29678,G29679,G29680,
       G29681,G29682,G29683,G29684,G29685,G29686,G29687,G29688,G29689,G29690,G29691,G29692,G29693,G29694,G29695,G29696,G29697,G29698,G29699,G29700,
       G29701,G29702,G29703,G29704,G29705,G29706,G29707,G29708,G29709,G29710,G29711,G29712,G29713,G29714,G29715,G29716,G29717,G29718,G29719,G29720,
       G29721,G29722,G29723,G29724,G29725,G29726,G29727,G29728,G29729,G29730,G29731,G29732,G29733,G29734,G29735,G29736,G29737,G29738,G29739,G29740,
       G29741,G29742,G29743,G29744,G29745,G29746,G29747,G29748,G29749,G29750,G29751,G29752,G29753,G29754,G29755,G29756,G29757,G29758,G29759,G29760,
       G29761,G29762,G29763,G29764,G29765,G29766,G29767,G29768,G29769,G29770,G29771,G29772,G29773,G29774,G29775,G29776,G29777,G29778,G29779,G29780,
       G29781,G29782,G29783,G29784,G29785,G29786,G29787,G29788,G29789,G29790,G29791,G29792,G29793,G29794,G29795,G29796,G29797,G29798,G29799,G29800,
       G29801,G29802,G29803,G29804,G29805,G29806,G29807,G29808,G29809,G29810,G29811,G29812,G29813,G29814,G29815,G29816,G29817,G29818,G29819,G29820,
       G29821,G29822,G29823,G29824,G29825,G29826,G29827,G29828,G29829,G29830,G29831,G29832,G29833,G29834,G29835,G29836,G29837,G29838,G29839,G29840,
       G29841,G29842,G29843,G29844,G29845,G29846,G29847,G29848,G29849,G29850,G29851,G29852,G29853,G29854,G29855,G29856,G29857,G29858,G29859,G29860,
       G29861,G29862,G29863,G29864,G29865,G29866,G29867,G29868,G29869,G29870,G29871,G29872,G29873,G29874,G29875,G29876,G29877,G29878,G29879,G29880,
       G29881,G29882,G29883,G29884,G29885,G29886,G29887,G29888,G29889,G29890,G29891,G29892,G29893,G29894,G29895,G29896,G29897,G29898,G29899,G29900,
       G29901,G29902,G29903,G29904,G29905,G29906,G29907,G29908,G29909,G29910,G29911,G29912,G29913,G29914,G29915,G29916,G29917,G29918,G29919,G29920,
       G29921,G29922,G29923,G29924,G29925,G29926,G29927,G29928,G29929,G29930,G29931,G29932,G29933,G29934,G29935,G29936,G29937,G29938,G29939,G29940,
       G29941,G29942,G29943,G29944,G29945,G29946,G29947,G29948,G29949,G29950,G29951,G29952,G29953,G29954,G29955,G29956,G29957,G29958,G29959,G29960,
       G29961,G29962,G29963,G29964,G29965,G29966,G29967,G29968,G29969,G29970,G29971,G29972,G29973,G29974,G29975,G29976,G29977,G29978,G29979,G29980,
       G29981,G29982,G29983,G29984,G29985,G29986,G29987,G29988,G29989,G29990,G29991,G29992,G29993,G29994,G29995,G29996,G29997,G29998,G29999,G30000,
       G30001,G30002,G30003,G30004,G30005,G30006,G30007,G30008,G30009,G30010,G30011,G30012,G30013,G30014,G30015,G30016,G30017,G30018,G30019,G30020,
       G30021,G30022,G30023,G30024,G30025,G30026,G30027,G30028,G30029,G30030,G30031,G30032,G30033,G30034,G30035,G30036,G30037,G30038,G30039,G30040,
       G30041,G30042,G30043,G30044,G30045,G30046,G30047,G30048,G30049,G30050,G30051,G30052,G30053,G30054,G30055,G30056,G30057,G30058,G30059,G30060,
       G30061,G30062,G30063,G30064,G30065,G30066,G30067,G30068,G30069,G30070,G30071,G30072,G30073,G30074,G30075,G30076,G30077,G30078,G30079,G30080,
       G30081,G30082,G30083,G30084,G30085,G30086,G30087,G30088,G30089,G30090,G30091,G30092,G30093,G30094,G30095,G30096,G30097,G30098,G30099,G30100,
       G30101,G30102,G30103,G30104,G30105,G30106,G30107,G30108,G30109,G30110,G30111,G30112,G30113,G30114,G30115,G30116,G30117,G30118,G30119,G30120,
       G30121,G30122,G30123,G30124,G30125,G30126,G30127,G30128,G30129,G30130,G30131,G30132,G30133,G30134,G30135,G30136,G30137,G30138,G30139,G30140,
       G30141,G30142,G30143,G30144,G30145,G30146,G30147,G30148,G30149,G30150,G30151,G30152,G30153,G30154,G30155,G30156,G30157,G30158,G30159,G30160,
       G30161,G30162,G30163,G30164,G30165,G30166,G30167,G30168,G30169,G30170,G30171,G30172,G30173,G30174,G30175,G30176,G30177,G30178,G30179,G30180,
       G30181,G30182,G30183,G30184,G30185,G30186,G30187,G30188,G30189,G30190,G30191,G30192,G30193,G30194,G30195,G30196,G30197,G30198,G30199,G30200,
       G30201,G30202,G30203,G30204,G30205,G30206,G30207,G30208,G30209,G30210,G30211,G30212,G30213,G30214,G30215,G30216,G30217,G30218,G30219,G30220,
       G30221,G30222,G30223,G30224,G30225,G30226,G30227,G30228,G30229,G30230,G30231,G30232,G30233,G30234,G30235,G30236,G30237,G30238,G30239,G30240,
       G30241,G30242,G30243,G30244,G30245,G30246,G30247,G30248,G30249,G30250,G30251,G30252,G30253,G30254,G30255,G30256,G30257,G30258,G30259,G30260,
       G30261,G30262,G30263,G30264,G30265,G30266,G30267,G30268,G30269,G30270,G30271,G30272,G30273,G30274,G30275,G30276,G30277,G30278,G30279,G30280,
       G30281,G30282,G30283,G30284,G30285,G30286,G30287,G30288,G30289,G30290,G30291,G30292,G30293,G30294,G30295,G30296,G30297,G30298,G30299,G30300,
       G30301,G30302,G30303,G30304,G30305,G30306,G30307,G30308,G30309,G30310,G30311,G30312,G30313,G30314,G30315,G30316,G30317,G30318,G30319,G30320,
       G30321,G30322,G30323,G30324,G30325,G30326,G30327,G30328,G30329,G30330,G30331,G30332,G30333,G30334,G30335,G30336,G30337,G30338,G30339,G30340,
       G30341,G30342,G30343,G30344,G30345,G30346,G30347,G30348,G30349,G30350,G30351,G30352,G30353,G30354,G30355,G30356,G30357,G30358,G30359,G30360,
       G30361,G30362,G30363,G30364,G30365,G30366,G30367,G30368,G30369,G30370,G30371,G30372,G30373,G30374,G30375,G30376,G30377,G30378,G30379,G30380,
       G30381,G30382,G30383,G30384,G30385,G30386,G30387,G30388,G30389,G30390,G30391,G30392,G30393,G30394,G30395,G30396,G30397,G30398,G30399,G30400,
       G30401,G30402,G30403,G30404,G30405,G30406,G30407,G30408,G30409,G30410,G30411,G30412,G30413,G30414,G30415,G30416,G30417,G30418,G30419,G30420,
       G30421,G30422,G30423,G30424,G30425,G30426,G30427,G30428,G30429,G30430,G30431,G30432,G30433,G30434,G30435,G30436,G30437,G30438,G30439,G30440,
       G30441,G30442,G30443,G30444,G30445,G30446,G30447,G30448,G30449,G30450,G30451,G30452,G30453,G30454,G30455,G30456,G30457,G30458,G30459,G30460,
       G30461,G30462,G30463,G30464,G30465,G30466,G30467,G30468,G30469,G30470,G30471,G30472,G30473,G30474,G30475,G30476,G30477,G30478,G30479,G30480,
       G30481,G30482,G30483,G30484,G30485,G30486,G30487,G30488,G30489,G30490,G30491,G30492,G30493,G30494,G30495,G30496,G30497,G30498,G30499,G30500,
       G30501,G30502,G30503,G30504,G30505,G30506,G30507,G30508,G30509,G30510,G30511,G30512,G30513,G30514,G30515,G30516,G30517,G30518,G30519,G30520,
       G30521,G30522,G30523,G30524,G30525,G30526,G30527,G30528,G30529,G30530,G30531,G30532,G30533,G30534,G30535,G30536,G30537,G30538,G30539,G30540,
       G30541,G30542,G30543,G30544,G30545,G30546,G30547,G30548,G30549,G30550,G30551,G30552,G30553,G30554,G30555,G30556,G30557,G30558,G30559,G30560,
       G30561,G30562,G30563,G30564,G30565,G30566,G30567,G30568,G30569,G30570,G30571,G30572,G30573,G30574,G30575,G30576,G30577,G30578,G30579,G30580,
       G30581,G30582,G30583,G30584,G30585,G30586,G30587,G30588,G30589,G30590,G30591,G30592,G30593,G30594,G30595,G30596,G30597,G30598,G30599,G30600,
       G30601,G30602,G30603,G30604,G30605,G30606,G30607,G30608,G30609,G30610,G30611,G30612,G30613,G30614,G30615,G30616,G30617,G30618,G30619,G30620,
       G30621,G30622,G30623,G30624,G30625,G30626,G30627,G30628,G30629,G30630,G30631,G30632,G30633,G30634,G30635,G30636,G30637,G30638,G30639,G30640,
       G30641,G30642,G30643,G30644,G30645,G30646,G30647,G30648,G30649,G30650,G30651,G30652,G30653,G30654,G30655,G30656,G30657,G30658,G30659,G30660,
       G30661,G30662,G30663,G30664,G30665,G30666,G30667,G30668,G30669,G30670,G30671,G30672,G30673,G30674,G30675,G30676,G30677,G30678,G30679,G30680,
       G30681,G30682,G30683,G30684,G30685,G30686,G30687,G30688,G30689,G30690,G30691,G30692,G30693,G30694,G30695,G30696,G30697,G30698,G30699,G30700,
       G30701,G30702,G30703,G30704,G30705,G30706,G30707,G30708,G30709,G30710,G30711,G30712,G30713,G30714,G30715,G30716,G30717,G30718,G30719,G30720,
       G30721,G30722,G30723,G30724,G30725,G30726,G30727,G30728,G30729,G30730,G30731,G30732,G30733,G30734,G30735,G30736,G30737,G30738,G30739,G30740,
       G30741,G30742,G30743,G30744,G30745,G30746,G30747,G30748,G30749,G30750,G30751,G30752,G30753,G30754,G30755,G30756,G30757,G30758,G30759,G30760,
       G30761,G30762,G30763,G30764,G30765,G30766,G30767,G30768,G30769,G30770,G30771,G30772,G30773,G30774,G30775,G30776,G30777,G30778,G30779,G30780,
       G30781,G30782,G30783,G30784,G30785,G30786,G30787,G30788,G30789,G30790,G30791,G30792,G30793,G30794,G30795,G30796,G30797,G30798,G30799,G30800,
       G30801,G30802,G30803,G30804,G30805,G30806,G30807,G30808,G30809,G30810,G30811,G30812,G30813,G30814,G30815,G30816,G30817,G30818,G30819,G30820,
       G30821,G30822,G30823,G30824,G30825,G30826,G30827,G30828,G30829,G30830,G30831,G30832,G30833,G30834,G30835,G30836,G30837,G30838,G30839,G30840,
       G30841,G30842,G30843,G30844,G30845,G30846,G30847,G30848,G30849,G30850,G30851,G30852,G30853,G30854,G30855,G30856,G30857,G30858,G30859,G30860,
       G30861,G30862,G30863,G30864,G30865,G30866,G30867,G30868,G30869,G30870,G30871,G30872,G30873,G30874,G30875,G30876,G30877,G30878,G30879,G30880,
       G30881,G30882,G30883,G30884,G30885,G30886,G30887,G30888,G30889,G30890,G30891,G30892,G30893,G30894,G30895,G30896,G30897,G30898,G30899,G30900,
       G30901,G30902,G30903,G30904,G30905,G30906,G30907,G30908,G30909,G30910,G30911,G30912,G30913,G30914,G30915,G30916,G30917,G30918,G30919,G30920,
       G30921,G30922,G30923,G30924,G30925,G30926,G30927,G30928,G30929,G30930,G30931,G30932,G30933,G30934,G30935,G30936,G30937,G30938,G30939,G30940,
       G30941,G30942,G30943,G30944,G30945,G30946,G30947,G30948,G30949,G30950,G30951,G30952,G30953,G30954,G30955,G30956,G30957,G30958,G30959,G30960,
       G30961,G30962,G30963,G30964,G30965,G30966,G30967,G30968,G30969,G30970,G30971,G30972,G30973,G30974,G30975,G30976,G30977,G30978,G30979,G30980,
       G30981,G30982,G30983,G30984,G30985,G30986,G30987,G30988,G30989,G30990,G30991,G30992,G30993,G30994,G30995,G30996,G30997,G30998,G30999,G31000,
       G31001,G31002,G31003,G31004,G31005,G31006,G31007,G31008,G31009,G31010,G31011,G31012,G31013,G31014,G31015,G31016,G31017,G31018,G31019,G31020,
       G31021,G31022,G31023,G31024,G31025,G31026,G31027,G31028,G31029,G31030,G31031,G31032,G31033,G31034,G31035,G31036,G31037,G31038,G31039,G31040,
       G31041,G31042,G31043,G31044,G31045,G31046,G31047,G31048,G31049,G31050,G31051,G31052,G31053,G31054,G31055,G31056,G31057,G31058,G31059,G31060,
       G31061,G31062,G31063,G31064,G31065,G31066,G31067,G31068,G31069,G31070,G31071,G31072,G31073,G31074,G31075,G31076,G31077,G31078,G31079,G31080,
       G31081,G31082,G31083,G31084,G31085,G31086,G31087,G31088,G31089,G31090,G31091,G31092,G31093,G31094,G31095,G31096,G31097,G31098,G31099,G31100,
       G31101,G31102,G31103,G31104,G31105,G31106,G31107,G31108,G31109,G31110,G31111,G31112,G31113,G31114,G31115,G31116,G31117,G31118,G31119,G31120,
       G31121,G31122,G31123,G31124,G31125,G31126,G31127,G31128,G31129,G31130,G31131,G31132,G31133,G31134,G31135,G31136,G31137,G31138,G31139,G31140,
       G31141,G31142,G31143,G31144,G31145,G31146,G31147,G31148,G31149,G31150,G31151,G31152,G31153,G31154,G31155,G31156,G31157,G31158,G31159,G31160,
       G31161,G31162,G31163,G31164,G31165,G31166,G31167,G31168,G31169,G31170,G31171,G31172,G31173,G31174,G31175,G31176,G31177,G31178,G31179,G31180,
       G31181,G31182,G31183,G31184,G31185,G31186,G31187,G31188,G31189,G31190,G31191,G31192,G31193,G31194,G31195,G31196,G31197,G31198,G31199,G31200,
       G31201,G31202,G31203,G31204,G31205,G31206,G31207,G31208,G31209,G31210,G31211,G31212,G31213,G31214,G31215,G31216,G31217,G31218,G31219,G31220,
       G31221,G31222,G31223,G31224,G31225,G31226,G31227,G31228,G31229,G31230,G31231,G31232,G31233,G31234,G31235,G31236,G31237,G31238,G31239,G31240,
       G31241,G31242,G31243,G31244,G31245,G31246,G31247,G31248,G31249,G31250,G31251,G31252,G31253,G31254,G31255,G31256,G31257,G31258,G31259,G31260,
       G31261,G31262,G31263,G31264,G31265,G31266,G31267,G31268,G31269,G31270,G31271,G31272,G31273,G31274,G31275,G31276,G31277,G31278,G31279,G31280,
       G31281,G31282,G31283,G31284,G31285,G31286,G31287,G31288,G31289,G31290,G31291,G31292,G31293,G31294,G31295,G31296,G31297,G31298,G31299,G31300,
       G31301,G31302,G31303,G31304,G31305,G31306,G31307,G31308,G31309,G31310,G31311,G31312,G31313,G31314,G31315,G31316,G31317,G31318,G31319,G31320,
       G31321,G31322,G31323,G31324,G31325,G31326,G31327,G31328,G31329,G31330,G31331,G31332,G31333,G31334,G31335,G31336,G31337,G31338,G31339,G31340,
       G31341,G31342,G31343,G31344,G31345,G31346,G31347,G31348,G31349,G31350,G31351,G31352,G31353,G31354,G31355,G31356,G31357,G31358,G31359,G31360,
       G31361,G31362,G31363,G31364,G31365,G31366,G31367,G31368,G31369,G31370,G31371,G31372,G31373,G31374,G31375,G31376,G31377,G31378,G31379,G31380,
       G31381,G31382,G31383,G31384,G31385,G31386,G31387,G31388,G31389,G31390,G31391,G31392,G31393,G31394,G31395,G31396,G31397,G31398,G31399,G31400,
       G31401,G31402,G31403,G31404,G31405,G31406,G31407,G31408,G31409,G31410,G31411,G31412,G31413,G31414,G31415,G31416,G31417,G31418,G31419,G31420,
       G31421,G31422,G31423,G31424,G31425,G31426,G31427,G31428,G31429,G31430,G31431,G31432,G31433,G31434,G31435,G31436,G31437,G31438,G31439,G31440,
       G31441,G31442,G31443,G31444,G31445,G31446,G31447,G31448,G31449,G31450,G31451,G31452,G31453,G31454,G31455,G31456,G31457,G31458,G31459,G31460,
       G31461,G31462,G31463,G31464,G31465,G31466,G31467,G31468,G31469,G31470,G31471,G31472,G31473,G31474,G31475,G31476,G31477,G31478,G31479,G31480,
       G31481,G31482,G31483,G31484,G31485,G31486,G31487,G31488,G31489,G31490,G31491,G31492,G31493,G31494,G31495,G31496,G31497,G31498,G31499,G31500,
       G31501,G31502,G31503,G31504,G31505,G31506,G31507,G31508,G31509,G31510,G31511,G31512,G31513,G31514,G31515,G31516,G31517,G31518,G31519,G31520,
       G31521,G31522,G31523,G31524,G31525,G31526,G31527,G31528,G31529,G31530,G31531,G31532,G31533,G31534,G31535,G31536,G31537,G31538,G31539,G31540,
       G31541,G31542,G31543,G31544,G31545,G31546,G31547,G31548,G31549,G31550,G31551,G31552,G31553,G31554,G31555,G31556,G31557,G31558,G31559,G31560,
       G31561,G31562,G31563,G31564,G31565,G31566,G31567,G31568,G31569,G31570,G31571,G31572,G31573,G31574,G31575,G31576,G31577,G31578,G31579,G31580,
       G31581,G31582,G31583,G31584,G31585,G31586,G31587,G31588,G31589,G31590,G31591,G31592,G31593,G31594,G31595,G31596,G31597,G31598,G31599,G31600,
       G31601,G31602,G31603,G31604,G31605,G31606,G31607,G31608,G31609,G31610,G31611,G31612,G31613,G31614,G31615,G31616,G31617,G31618,G31619,G31620,
       G31621,G31622,G31623,G31624,G31625,G31626,G31627,G31628,G31629,G31630,G31631,G31632,G31633,G31634,G31635,G31636,G31637,G31638,G31639,G31640,
       G31641,G31642,G31643,G31644,G31645,G31646,G31647,G31648,G31649,G31650,G31651,G31652,G31653,G31654,G31655,G31656,G31657,G31658,G31659,G31660,
       G31661,G31662,G31663,G31664,G31665,G31666,G31667,G31668,G31669,G31670,G31671,G31672,G31673,G31674,G31675,G31676,G31677,G31678,G31679,G31680,
       G31681,G31682,G31683,G31684,G31685,G31686,G31687,G31688,G31689,G31690,G31691,G31692,G31693,G31694,G31695,G31696,G31697,G31698,G31699,G31700,
       G31701,G31702,G31703,G31704,G31705,G31706,G31707,G31708,G31709,G31710,G31711,G31712,G31713,G31714,G31715,G31716,G31717,G31718,G31719,G31720,
       G31721,G31722,G31723,G31724,G31725,G31726,G31727,G31728,G31729,G31730,G31731,G31732,G31733,G31734,G31735,G31736,G31737,G31738,G31739,G31740,
       G31741,G31742,G31743,G31744,G31745,G31746,G31747,G31748,G31749,G31750,G31751,G31752,G31753,G31754,G31755,G31756,G31757,G31758,G31759,G31760,
       G31761,G31762,G31763,G31764,G31765,G31766,G31767,G31768,G31769,G31770,G31771,G31772,G31773,G31774,G31775,G31776,G31777,G31778,G31779,G31780,
       G31781,G31782,G31783,G31784,G31785,G31786,G31787,G31788,G31789,G31790,G31791,G31792,G31793,G31794,G31795,G31796,G31797,G31798,G31799,G31800,
       G31801,G31802,G31803,G31804,G31805,G31806,G31807,G31808,G31809,G31810,G31811,G31812,G31813,G31814,G31815,G31816,G31817,G31818,G31819,G31820,
       G31821,G31822,G31823,G31824,G31825,G31826,G31827,G31828,G31829,G31830,G31831,G31832,G31833,G31834,G31835,G31836,G31837,G31838,G31839,G31840,
       G31841,G31842,G31843,G31844,G31845,G31846,G31847,G31848,G31849,G31850,G31851,G31852,G31853,G31854,G31855,G31856,G31857,G31858,G31859,G31860,
       G31861,G31862,G31863,G31864,G31865,G31866,G31867,G31868,G31869,G31870,G31871,G31872,G31873,G31874,G31875,G31876,G31877,G31878,G31879,G31880,
       G31881,G31882,G31883,G31884,G31885,G31886,G31887,G31888,G31889,G31890,G31891,G31892,G31893,G31894,G31895,G31896,G31897,G31898,G31899,G31900,
       G31901,G31902,G31903,G31904,G31905,G31906,G31907,G31908,G31909,G31910,G31911,G31912,G31913,G31914,G31915,G31916,G31917,G31918,G31919,G31920,
       G31921,G31922,G31923,G31924,G31925,G31926,G31927,G31928,G31929,G31930,G31931,G31932,G31933,G31934,G31935,G31936,G31937,G31938,G31939,G31940,
       G31941,G31942,G31943,G31944,G31945,G31946,G31947,G31948,G31949,G31950,G31951,G31952,G31953,G31954,G31955,G31956,G31957,G31958,G31959,G31960,
       G31961,G31962,G31963,G31964,G31965,G31966,G31967,G31968,G31969,G31970,G31971,G31972,G31973,G31974,G31975,G31976,G31977,G31978,G31979,G31980,
       G31981,G31982,G31983,G31984,G31985,G31986,G31987,G31988,G31989,G31990,G31991,G31992,G31993,G31994,G31995,G31996,G31997,G31998,G31999,G32000,
       G32001,G32002,G32003,G32004,G32005,G32006,G32007,G32008,G32009,G32010,G32011,G32012,G32013,G32014,G32015,G32016,G32017,G32018,G32019,G32020,
       G32021,G32022,G32023,G32024,G32025,G32026,G32027,G32028,G32029,G32030,G32031,G32032,G32033,G32034,G32035,G32036,G32037,G32038,G32039,G32040,
       G32041,G32042,G32043,G32044,G32045,G32046,G32047,G32048,G32049,G32050,G32051,G32052,G32053,G32054,G32055,G32056,G32057,G32058,G32059,G32060,
       G32061,G32062,G32063,G32064,G32065,G32066,G32067,G32068,G32069,G32070,G32071,G32072,G32073,G32074,G32075,G32076,G32077,G32078,G32079,G32080,
       G32081,G32082,G32083,G32084,G32085,G32086,G32087,G32088,G32089,G32090,G32091,G32092,G32093,G32094,G32095,G32096,G32097,G32098,G32099,G32100,
       G32101,G32102,G32103,G32104,G32105,G32106,G32107,G32108,G32109,G32110,G32111,G32112,G32113,G32114,G32115,G32116,G32117,G32118,G32119,G32120,
       G32121,G32122,G32123,G32124,G32125,G32126,G32127,G32128,G32129,G32130,G32131,G32132,G32133,G32134,G32135,G32136,G32137,G32138,G32139,G32140,
       G32141,G32142,G32143,G32144,G32145,G32146,G32147,G32148,G32149,G32150,G32151,G32152,G32153,G32154,G32155,G32156,G32157,G32158,G32159,G32160,
       G32161,G32162,G32163,G32164,G32165,G32166,G32167,G32168,G32169,G32170,G32171,G32172,G32173,G32174,G32175,G32176,G32177,G32178,G32179,G32180,
       G32181,G32182,G32183,G32184,G32185,G32186,G32187,G32188,G32189,G32190,G32191,G32192,G32193,G32194,G32195,G32196,G32197,G32198,G32199,G32200,
       G32201,G32202,G32203,G32204,G32205,G32206,G32207,G32208,G32209,G32210,G32211,G32212,G32213,G32214,G32215,G32216,G32217,G32218,G32219,G32220,
       G32221,G32222,G32223,G32224,G32225,G32226,G32227,G32228,G32229,G32230,G32231,G32232,G32233,G32234,G32235,G32236,G32237,G32238,G32239,G32240,
       G32241,G32242,G32243,G32244,G32245,G32246,G32247,G32248,G32249,G32250,G32251,G32252,G32253,G32254,G32255,G32256,G32257,G32258,G32259,G32260,
       G32261,G32262,G32263,G32264,G32265,G32266,G32267,G32268,G32269,G32270,G32271,G32272,G32273,G32274,G32275,G32276,G32277,G32278,G32279,G32280,
       G32281,G32282,G32283,G32284,G32285,G32286,G32287,G32288,G32289,G32290,G32291,G32292,G32293,G32294,G32295,G32296,G32297,G32298,G32299,G32300,
       G32301,G32302,G32303,G32304,G32305,G32306,G32307,G32308,G32309,G32310,G32311,G32312,G32313,G32314,G32315,G32316,G32317,G32318,G32319,G32320,
       G32321,G32322,G32323,G32324,G32325,G32326,G32327,G32328,G32329,G32330,G32331,G32332,G32333,G32334,G32335,G32336,G32337,G32338,G32339,G32340,
       G32341,G32342,G32343,G32344,G32345,G32346,G32347,G32348,G32349,G32350,G32351,G32352,G32353,G32354,G32355,G32356,G32357,G32358,G32359,G32360,
       G32361,G32362,G32363,G32364,G32365,G32366,G32367,G32368,G32369,G32370,G32371,G32372,G32373,G32374,G32375,G32376,G32377,G32378,G32379,G32380,
       G32381,G32382,G32383,G32384,G32385,G32386,G32387,G32388,G32389,G32390,G32391,G32392,G32393,G32394,G32395,G32396,G32397,G32398,G32399,G32400,
       G32401,G32402,G32403,G32404,G32405,G32406,G32407,G32408,G32409,G32410,G32411,G32412,G32413,G32414,G32415,G32416,G32417,G32418,G32419,G32420,
       G32421,G32422,G32423,G32424,G32425,G32426,G32427,G32428,G32429,G32430,G32431,G32432,G32433,G32434,G32435,G32436,G32437,G32438,G32439,G32440,
       G32441,G32442,G32443,G32444,G32445,G32446,G32447,G32448,G32449,G32450,G32451,G32452,G32453,G32454,G32455,G32456,G32457,G32458,G32459,G32460,
       G32461,G32462,G32463,G32464,G32465,G32466,G32467,G32468,G32469,G32470,G32471,G32472,G32473,G32474,G32475,G32476,G32477,G32478,G32479,G32480,
       G32481,G32482,G32483,G32484,G32485,G32486,G32487,G32488,G32489,G32490,G32491,G32492,G32493,G32494,G32495,G32496,G32497,G32498,G32499,G32500,
       G32501,G32502,G32503,G32504,G32505,G32506,G32507,G32508,G32509,G32510,G32511,G32512,G32513,G32514,G32515,G32516,G32517,G32518,G32519,G32520,
       G32521,G32522,G32523,G32524,G32525,G32526,G32527,G32528,G32529,G32530,G32531,G32532,G32533,G32534,G32535,G32536,G32537,G32538,G32539,G32540,
       G32541,G32542,G32543,G32544,G32545,G32546,G32547,G32548,G32549,G32550,G32551,G32552,G32553,G32554,G32555,G32556,G32557,G32558,G32559,G32560,
       G32561,G32562,G32563,G32564,G32565,G32566,G32567,G32568,G32569,G32570,G32571,G32572,G32573,G32574,G32575,G32576,G32577,G32578,G32579,G32580,
       G32581,G32582,G32583,G32584,G32585,G32586,G32587,G32588,G32589,G32590,G32591,G32592,G32593,G32594,G32595,G32596,G32597,G32598,G32599,G32600,
       G32601,G32602,G32603,G32604,G32605,G32606,G32607,G32608,G32609,G32610,G32611,G32612,G32613,G32614,G32615,G32616,G32617,G32618,G32619,G32620,
       G32621,G32622,G32623,G32624,G32625,G32626,G32627,G32628,G32629,G32630,G32631,G32632,G32633,G32634,G32635,G32636,G32637,G32638,G32639,G32640,
       G32641,G32642,G32643,G32644,G32645,G32646,G32647,G32648,G32649,G32650,G32651,G32652,G32653,G32654,G32655,G32656,G32657,G32658,G32659,G32660,
       G32661,G32662,G32663,G32664,G32665,G32666,G32667,G32668,G32669,G32670,G32671,G32672,G32673,G32674,G32675,G32676,G32677,G32678,G32679,G32680,
       G32681,G32682,G32683,G32684,G32685,G32686,G32687,G32688,G32689,G32690,G32691,G32692,G32693,G32694,G32695,G32696,G32697,G32698,G32699,G32700,
       G32701,G32702,G32703,G32704,G32705,G32706,G32707,G32708,G32709,G32710,G32711,G32712,G32713,G32714,G32715,G32716,G32717,G32718,G32719,G32720,
       G32721,G32722,G32723,G32724,G32725,G32726,G32727,G32728,G32729,G32730,G32731,G32732,G32733,G32734,G32735,G32736,G32737,G32738,G32739,G32740,
       G32741,G32742,G32743,G32744,G32745,G32746,G32747,G32748,G32749,G32750,G32751,G32752,G32753,G32754,G32755,G32756,G32757,G32758,G32759,G32760,
       G32761,G32762,G32763,G32764,G32765,G32766,G32767,G32768,G32769,G32770,G32771,G32772,G32773,G32774,G32775,G32776,G32777,G32778,G32779,G32780,
       G32781,G32782,G32783,G32784,G32785,G32786,G32787,G32788,G32789,G32790,G32791,G32792,G32793,G32794,G32795,G32796,G32797,G32798,G32799,G32800,
       G32801,G32802,G32803,G32804,G32805,G32806,G32807,G32808,G32809,G32810,G32811,G32812,G32813,G32814,G32815,G32816,G32817,G32818,G32819,G32820,
       G32821,G32822,G32823,G32824,G32825,G32826,G32827,G32828,G32829,G32830,G32831,G32832,G32833,G32834,G32835,G32836,G32837,G32838,G32839,G32840,
       G32841,G32842,G32843,G32844,G32845,G32846,G32847,G32848,G32849,G32850,G32851,G32852,G32853,G32854,G32855,G32856,G32857,G32858,G32859,G32860,
       G32861,G32862,G32863,G32864,G32865,G32866,G32867,G32868,G32869,G32870,G32871,G32872,G32873,G32874,G32875,G32876,G32877,G32878,G32879,G32880,
       G32881,G32882,G32883,G32884,G32885,G32886,G32887,G32888,G32889,G32890,G32891,G32892,G32893,G32894,G32895,G32896,G32897,G32898,G32899,G32900,
       G32901,G32902,G32903,G32904,G32905,G32906,G32907,G32908,G32909,G32910,G32911,G32912,G32913,G32914,G32915,G32916,G32917,G32918,G32919,G32920,
       G32921,G32922,G32923,G32924,G32925,G32926,G32927,G32928,G32929,G32930,G32931,G32932,G32933,G32934,G32935,G32936,G32937,G32938,G32939,G32940,
       G32941,G32942,G32943,G32944,G32945,G32946,G32947,G32948,G32949,G32950,G32951,G32952,G32953,G32954,G32955,G32956,G32957,G32958,G32959,G32960,
       G32961,G32962,G32963,G32964,G32965,G32966,G32967,G32968,G32969,G32970,G32971,G32972,G32973,G32974,G32975,G32976,G32977,G32978,G32979,G32980,
       G32981,G32982,G32983,G32984,G32985,G32986,G32987,G32988,G32989,G32990,G32991,G32992,G32993,G32994,G32995,G32996,G32997,G32998,G32999,G33000,
       G33001,G33002,G33003,G33004,G33005,G33006,G33007,G33008,G33009,G33010,G33011,G33012,G33013,G33014,G33015,G33016,G33017,G33018,G33019,G33020,
       G33021,G33022,G33023,G33024,G33025,G33026,G33027,G33028,G33029,G33030,G33031,G33032,G33033,G33034,G33035,G33036,G33037,G33038,G33039,G33040,
       G33041,G33042,G33043,G33044,G33045,G33046,G33047,G33048,G33049,G33050,G33051,G33052,G33053,G33054,G33055,G33056,G33057,G33058,G33059,G33060,
       G33061,G33062,G33063,G33064,G33065,G33066,G33067,G33068,G33069,G33070,G33071,G33072,G33073,G33074,G33075,G33076,G33077,G33078,G33079,G33080,
       G33081,G33082,G33083,G33084,G33085,G33086,G33087,G33088,G33089,G33090,G33091,G33092,G33093,G33094,G33095,G33096,G33097,G33098,G33099,G33100,
       G33101,G33102,G33103,G33104,G33105,G33106,G33107,G33108,G33109,G33110,G33111,G33112,G33113,G33114,G33115,G33116,G33117,G33118,G33119,G33120,
       G33121,G33122,G33123,G33124,G33125,G33126,G33127,G33128,G33129,G33130,G33131,G33132,G33133,G33134,G33135,G33136,G33137,G33138,G33139,G33140,
       G33141,G33142,G33143,G33144,G33145,G33146,G33147,G33148,G33149,G33150,G33151,G33152,G33153,G33154,G33155,G33156,G33157,G33158,G33159,G33160,
       G33161,G33162,G33163,G33164,G33165,G33166,G33167,G33168,G33169,G33170,G33171,G33172,G33173,G33174,G33175,G33176,G33177,G33178,G33179,G33180,
       G33181,G33182,G33183,G33184,G33185,G33186,G33187,G33188,G33189,G33190,G33191,G33192,G33193,G33194,G33195,G33196,G33197,G33198,G33199,G33200,
       G33201,G33202,G33203,G33204,G33205,G33206,G33207,G33208,G33209,G33210,G33211,G33212,G33213,G33214,G33215,G33216,G33217,G33218,G33219,G33220,
       G33221,G33222,G33223,G33224,G33225,G33226,G33227,G33228,G33229,G33230,G33231,G33232,G33233,G33234,G33235,G33236,G33237,G33238,G33239,G33240,
       G33241,G33242,G33243,G33244,G33245,G33246,G33247,G33248,G33249,G33250,G33251,G33252,G33253,G33254,G33255,G33256,G33257,G33258,G33259,G33260,
       G33261,G33262,G33263,G33264,G33265,G33266,G33267,G33268,G33269,G33270,G33271,G33272,G33273,G33274,G33275,G33276,G33277,G33278,G33279,G33280,
       G33281,G33282,G33283,G33284,G33285,G33286,G33287,G33288,G33289,G33290,G33291,G33292,G33293,G33294,G33295,G33296,G33297,G33298,G33299,G33300,
       G33301,G33302,G33303,G33304,G33305,G33306,G33307,G33308,G33309,G33310,G33311,G33312,G33313,G33314,G33315,G33316,G33317,G33318,G33319,G33320,
       G33321,G33322,G33323,G33324,G33325,G33326,G33327,G33328,G33329,G33330,G33331,G33332,G33333,G33334,G33335,G33336,G33337,G33338,G33339,G33340,
       G33341,G33342,G33343,G33344,G33345,G33346,G33347,G33348,G33349,G33350,G33351,G33352,G33353,G33354,G33355,G33356,G33357,G33358,G33359,G33360,
       G33361,G33362,G33363,G33364,G33365,G33366,G33367,G33368,G33369,G33370,G33371,G33372,G33373,G33374,G33375,G33376,G33377,G33378,G33379,G33380,
       G33381,G33382,G33383,G33384,G33385,G33386,G33387,G33388,G33389,G33390,G33391,G33392,G33393,G33394,G33395,G33396,G33397,G33398,G33399,G33400,
       G33401,G33402,G33403,G33404,G33405,G33406,G33407,G33408,G33409,G33410,G33411,G33412,G33413,G33414,G33415,G33416,G33417,G33418,G33419,G33420,
       G33421,G33422,G33423,G33424,G33425,G33426,G33427,G33428,G33429,G33430,G33431,G33432,G33433,G33434,G33435,G33436,G33437,G33438,G33439,G33440,
       G33441,G33442,G33443,G33444,G33445,G33446,G33447,G33448,G33449,G33450,G33451,G33452,G33453,G33454,G33455,G33456,G33457,G33458,G33459,G33460,
       G33461,G33462,G33463,G33464,G33465,G33466,G33467,G33468,G33469,G33470,G33471,G33472,G33473,G33474,G33475,G33476,G33477,G33478,G33479,G33480,
       G33481,G33482,G33483,G33484,G33485,G33486,G33487,G33488,G33489,G33490,G33491,G33492,G33493,G33494,G33495,G33496,G33497,G33498,G33499,G33500,
       G33501,G33502,G33503,G33504,G33505,G33506,G33507,G33508,G33509,G33510,G33511,G33512,G33513,G33514,G33515,G33516,G33517,G33518,G33519,G33520,
       G33521,G33522,G33523,G33524,G33525,G33526,G33527,G33528,G33529,G33530,G33531,G33532,G33533,G33534,G33535,G33536,G33537,G33538,G33539,G33540,
       G33541,G33542,G33543,G33544,G33545,G33546,G33547,G33548,G33549,G33550,G33551,G33552,G33553,G33554,G33555,G33556,G33557,G33558,G33559,G33560,
       G33561,G33562,G33563,G33564,G33565,G33566,G33567,G33568,G33569,G33570,G33571,G33572,G33573,G33574,G33575,G33576,G33577,G33578,G33579,G33580,
       G33581,G33582,G33583,G33584,G33585,G33586,G33587,G33588,G33589,G33590,G33591,G33592,G33593,G33594,G33595,G33596,G33597,G33598,G33599,G33600,
       G33601,G33602,G33603,G33604,G33605,G33606,G33607,G33608,G33609,G33610,G33611,G33612,G33613,G33614,G33615,G33616,G33617,G33618,G33619,G33620,
       G33621,G33622,G33623,G33624,G33625,G33626,G33627,G33628,G33629,G33630,G33631,G33632,G33633,G33634,G33635,G33636,G33637,G33638,G33639,G33640,
       G33641,G33642,G33643,G33644,G33645,G33646,G33647,G33648,G33649,G33650,G33651,G33652,G33653,G33654,G33655,G33656,G33657,G33658,G33659,G33660,
       G33661,G33662,G33663,G33664,G33665,G33666,G33667,G33668,G33669,G33670,G33671,G33672,G33673,G33674,G33675,G33676,G33677,G33678,G33679,G33680,
       G33681,G33682,G33683,G33684,G33685,G33686,G33687,G33688,G33689,G33690,G33691,G33692,G33693,G33694,G33695,G33696,G33697,G33698,G33699,G33700,
       G33701,G33702,G33703,G33704,G33705,G33706,G33707,G33708,G33709,G33710,G33711,G33712,G33713,G33714,G33715,G33716,G33717,G33718,G33719,G33720,
       G33721,G33722,G33723,G33724,G33725,G33726,G33727,G33728,G33729,G33730,G33731,G33732,G33733,G33734,G33735,G33736,G33737,G33738,G33739,G33740,
       G33741,G33742,G33743,G33744,G33745,G33746,G33747,G33748,G33749,G33750,G33751,G33752,G33753,G33754,G33755,G33756,G33757,G33758,G33759,G33760,
       G33761,G33762,G33763,G33764,G33765,G33766,G33767,G33768,G33769,G33770,G33771,G33772,G33773,G33774,G33775,G33776,G33777,G33778,G33779,G33780,
       G33781,G33782,G33783,G33784,G33785,G33786,G33787,G33788,G33789,G33790,G33791,G33792,G33793,G33794,G33795,G33796,G33797,G33798,G33799,G33800,
       G33801,G33802,G33803,G33804,G33805,G33806,G33807,G33808,G33809,G33810,G33811,G33812,G33813,G33814,G33815,G33816,G33817,G33818,G33819,G33820,
       G33821,G33822,G33823,G33824,G33825,G33826,G33827,G33828,G33829,G33830,G33831,G33832,G33833,G33834,G33835,G33836,G33837,G33838,G33839,G33840,
       G33841,G33842,G33843,G33844,G33845,G33846,G33847,G33848,G33849,G33850,G33851,G33852,G33853,G33854,G33855,G33856,G33857,G33858,G33859,G33860,
       G33861,G33862,G33863,G33864,G33865,G33866,G33867,G33868,G33869,G33870,G33871,G33872,G33873,G33874,G33875,G33876,G33877,G33878,G33879,G33880,
       G33881,G33882,G33883,G33884,G33885,G33886,G33887,G33888,G33889,G33890,G33891,G33892,G33893,G33894,G33895,G33896,G33897,G33898,G33899,G33900,
       G33901,G33902,G33903,G33904,G33905,G33906,G33907,G33908,G33909,G33910,G33911,G33912,G33913,G33914,G33915,G33916,G33917,G33918,G33919,G33920,
       G33921,G33922,G33923,G33924,G33925,G33926,G33927,G33928,G33929,G33930,G33931,G33932,G33933,G33934,G33935,G33936,G33937,G33938,G33939,G33940,
       G33941,G33942,G33943,G33944,G33945,G33946,G33947,G33948,G33949,G33950,G33951,G33952,G33953,G33954,G33955,G33956,G33957,G33958,G33959,G33960,
       G33961,G33962,G33963,G33964,G33965,G33966,G33967,G33968,G33969,G33970,G33971,G33972,G33973,G33974,G33975,G33976,G33977,G33978,G33979,G33980,
       G33981,G33982,G33983,G33984,G33985,G33986,G33987,G33988,G33989,G33990,G33991,G33992,G33993,G33994,G33995,G33996,G33997,G33998,G33999,G34000,
       G34001,G34002,G34003,G34004,G34005,G34006,G34007,G34008,G34009,G34010,G34011,G34012,G34013,G34014,G34015,G34016,G34017,G34018,G34019,G34020,
       G34021,G34022,G34023,G34024,G34025,G34026,G34027,G34028,G34029,G34030,G34031,G34032,G34033,G34034,G34035,G34036,G34037,G34038,G34039,G34040,
       G34041,G34042,G34043,G34044,G34045,G34046,G34047,G34048,G34049,G34050,G34051,G34052,G34053,G34054,G34055,G34056,G34057,G34058,G34059,G34060,
       G34061,G34062,G34063,G34064,G34065,G34066,G34067,G34068,G34069,G34070,G34071,G34072,G34073,G34074,G34075,G34076,G34077,G34078,G34079,G34080,
       G34081,G34082,G34083,G34084,G34085,G34086,G34087,G34088,G34089,G34090,G34091,G34092,G34093,G34094,G34095,G34096,G34097,G34098,G34099,G34100,
       G34101,G34102,G34103,G34104,G34105,G34106,G34107,G34108,G34109,G34110,G34111,G34112,G34113,G34114,G34115,G34116,G34117,G34118,G34119,G34120,
       G34121,G34122,G34123,G34124,G34125,G34126,G34127,G34128,G34129,G34130,G34131,G34132,G34133,G34134,G34135,G34136,G34137,G34138,G34139,G34140,
       G34141,G34142,G34143,G34144,G34145,G34146,G34147,G34148,G34149,G34150,G34151,G34152,G34153,G34154,G34155,G34156,G34157,G34158,G34159,G34160,
       G34161,G34162,G34163,G34164,G34165,G34166,G34167,G34168,G34169,G34170,G34171,G34172,G34173,G34174,G34175,G34176,G34177,G34178,G34179,G34180,
       G34181,G34182,G34183,G34184,G34185,G34186,G34187,G34188,G34189,G34190,G34191,G34192,G34193,G34194,G34195,G34196,G34197,G34198,G34199,G34200,
       G34201,G34202,G34203,G34204,G34205,G34206,G34207,G34208,G34209,G34210,G34211,G34212,G34213,G34214,G34215,G34216,G34217,G34218,G34219,G34220,
       G34221,G34222,G34223,G34224,G34225,G34226,G34227,G34228,G34229,G34230,G34231,G34232,G34233,G34234,G34235,G34236,G34237,G34238,G34239,G34240,
       G34241,G34242,G34243,G34244,G34245,G34246,G34247,G34248,G34249,G34250,G34251,G34252,G34253,G34254,G34255,G34256,G34257,G34258,G34259,G34260,
       G34261,G34262,G34263,G34264,G34265,G34266,G34267,G34268,G34269,G34270,G34271,G34272,G34273,G34274,G34275,G34276,G34277,G34278,G34279,G34280,
       G34281,G34282,G34283,G34284,G34285,G34286,G34287,G34288,G34289,G34290,G34291,G34292,G34293,G34294,G34295,G34296,G34297,G34298,G34299,G34300,
       G34301,G34302,G34303,G34304,G34305,G34306,G34307,G34308,G34309,G34310,G34311,G34312,G34313,G34314,G34315,G34316,G34317,G34318,G34319,G34320,
       G34321,G34322,G34323,G34324,G34325,G34326,G34327,G34328,G34329,G34330,G34331,G34332,G34333,G34334,G34335,G34336,G34337,G34338,G34339,G34340,
       G34341,G34342,G34343,G34344,G34345,G34346,G34347,G34348,G34349,G34350,G34351,G34352,G34353,G34354,G34355,G34356,G34357,G34358,G34359,G34360,
       G34361,G34362,G34363,G34364,G34365,G34366,G34367,G34368,G34369,G34370,G34371,G34372,G34373,G34374,G34375,G34376,G34377,G34378,G34379,G34380,
       G34381,G34382,G34383,G34384,G34385,G34386,G34387,G34388,G34389,G34390,G34391,G34392,G34393,G34394,G34395,G34396,G34397,G34398,G34399,G34400,
       G34401,G34402,G34403,G34404,G34405,G34406,G34407,G34408,G34409,G34410,G34411,G34412,G34413,G34414,G34415,G34416,G34417,G34418,G34419,G34420,
       G34421,G34422,G34423,G34424,G34425,G34426,G34427,G34428,G34429,G34430,G34431,G34432,G34433,G34434,G34435,G34436,G34437,G34438,G34439,G34440,
       G34441,G34442,G34443,G34444,G34445,G34446,G34447,G34448,G34449,G34450,G34451,G34452,G34453,G34454,G34455,G34456,G34457,G34458,G34459,G34460,
       G34461,G34462,G34463,G34464,G34465,G34466,G34467,G34468,G34469,G34470,G34471,G34472,G34473,G34474,G34475,G34476,G34477,G34478,G34479,G34480,
       G34481,G34482,G34483,G34484,G34485,G34486,G34487,G34488,G34489,G34490,G34491,G34492,G34493,G34494,G34495,G34496,G34497,G34498,G34499,G34500,
       G34501,G34502,G34503,G34504,G34505,G34506,G34507,G34508,G34509,G34510,G34511,G34512,G34513,G34514,G34515,G34516,G34517,G34518,G34519,G34520,
       G34521,G34522,G34523,G34524,G34525,G34526,G34527,G34528,G34529,G34530,G34531,G34532,G34533,G34534,G34535,G34536,G34537,G34538,G34539,G34540,
       G34541,G34542,G34543,G34544,G34545,G34546,G34547,G34548,G34549,G34550,G34551,G34552,G34553,G34554,G34555,G34556,G34557,G34558,G34559,G34560,
       G34561,G34562,G34563,G34564,G34565,G34566,G34567,G34568,G34569,G34570,G34571,G34572,G34573,G34574,G34575,G34576,G34577,G34578,G34579,G34580,
       G34581,G34582,G34583,G34584,G34585,G34586,G34587,G34588,G34589,G34590,G34591,G34592,G34593,G34594,G34595,G34596,G34597,G34598,G34599,G34600,
       G34601,G34602,G34603,G34604,G34605,G34606,G34607,G34608,G34609,G34610,G34611,G34612,G34613,G34614,G34615,G34616,G34617,G34618,G34619,G34620,
       G34621,G34622,G34623,G34624,G34625,G34626,G34627,G34628,G34629,G34630,G34631,G34632,G34633,G34634,G34635,G34636,G34637,G34638,G34639,G34640,
       G34641,G34642,G34643,G34644,G34645,G34646,G34647,G34648,G34649,G34650,G34651,G34652,G34653,G34654,G34655,G34656,G34657,G34658,G34659,G34660,
       G34661,G34662,G34663,G34664,G34665,G34666,G34667,G34668,G34669,G34670,G34671,G34672,G34673,G34674,G34675,G34676,G34677,G34678,G34679,G34680,
       G34681,G34682,G34683,G34684,G34685,G34686,G34687,G34688,G34689,G34690,G34691,G34692,G34693,G34694,G34695,G34696,G34697,G34698,G34699,G34700,
       G34701,G34702,G34703,G34704,G34705,G34706,G34707,G34708,G34709,G34710,G34711,G34712,G34713,G34714,G34715,G34716,G34717,G34718,G34719,G34720,
       G34721,G34722,G34723,G34724,G34725,G34726,G34727,G34728,G34729,G34730,G34731,G34732,G34733,G34734,G34735,G34736,G34737,G34738,G34739,G34740,
       G34741,G34742,G34743,G34744,G34745,G34746,G34747,G34748,G34749,G34750,G34751,G34752,G34753,G34754,G34755,G34756,G34757,G34758,G34759,G34760,
       G34761,G34762,G34763,G34764,G34765,G34766,G34767,G34768,G34769,G34770,G34771,G34772,G34773,G34774,G34775,G34776,G34777,G34778,G34779,G34780,
       G34781,G34782,G34783,G34784,G34785,G34786,G34787,G34788,G34789,G34790,G34791,G34792,G34793,G34794,G34795,G34796,G34797,G34798,G34799,G34800,
       G34801,G34802,G34803,G34804,G34805,G34806,G34807,G34808,G34809,G34810,G34811,G34812,G34813,G34814,G34815,G34816,G34817,G34818,G34819,G34820,
       G34821,G34822,G34823,G34824,G34825,G34826,G34827,G34828,G34829,G34830,G34831,G34832,G34833,G34834,G34835,G34836,G34837,G34838,G34839,G34840,
       G34841,G34842,G34843,G34844,G34845,G34846,G34847,G34848,G34849,G34850,G34851,G34852,G34853,G34854,G34855,G34856,G34857,G34858,G34859,G34860,
       G34861,G34862,G34863,G34864,G34865,G34866,G34867,G34868,G34869,G34870,G34871,G34872,G34873,G34874,G34875,G34876,G34877,G34878,G34879,G34880,
       G34881,G34882,G34883,G34884,G34885,G34886,G34887,G34888,G34889,G34890,G34891,G34892,G34893,G34894,G34895,G34896,G34897,G34898,G34899,G34900,
       G34901,G34902,G34903,G34904,G34905,G34906,G34907,G34908,G34909,G34910,G34911,G34912,G34913,G34914,G34915,G34916,G34917,G34918,G34919,G34920,
       G34921,G34922,G34923,G34924,G34925,G34926,G34927,G34928,G34929,G34930,G34931,G34932,G34933,G34934,G34935,G34936,G34937,G34938,G34939,G34940,
       G34941,G34942,G34943,G34944,G34945,G34946,G34947,G34948,G34949,G34950,G34951,G34952,G34953,G34954,G34955,G34956,G34957,G34958,G34959,G34960,
       G34961,G34962,G34963,G34964,G34965,G34966,G34967,G34968,G34969,G34970,G34971,G34972,G34973,G34974,G34975,G34976,G34977,G34978,G34979,G34980,
       G34981,G34982,G34983,G34984,G34985,G34986,G34987,G34988,G34989,G34990,G34991,G34992,G34993,G34994,G34995,G34996,G34997,G34998,G34999,G35000,
       G35001,G35002,G35003,G35004,G35005,G35006,G35007,G35008,G35009,G35010,G35011,G35012,G35013,G35014,G35015,G35016,G35017,G35018,G35019,G35020,
       G35021,G35022,G35023,G35024,G35025,G35026,G35027,G35028,G35029,G35030,G35031,G35032,G35033,G35034,G35035,G35036,G35037,G35038,G35039,G35040,
       G35041,G35042,G35043,G35044,G35045,G35046,G35047,G35048,G35049,G35050,G35051,G35052,G35053,G35054,G35055,G35056,G35057,G35058,G35059,G35060,
       G35061,G35062,G35063,G35064,G35065,G35066,G35067,G35068,G35069,G35070,G35071,G35072,G35073,G35074,G35075,G35076,G35077,G35078,G35079,G35080,
       G35081,G35082,G35083,G35084,G35085,G35086,G35087,G35088,G35089,G35090,G35091,G35092,G35093,G35094,G35095,G35096,G35097,G35098,G35099,G35100,
       G35101,G35102,G35103,G35104,G35105,G35106,G35107,G35108,G35109,G35110,G35111,G35112,G35113,G35114,G35115,G35116,G35117,G35118,G35119,G35120,
       G35121,G35122,G35123,G35124,G35125,G35126,G35127,G35128,G35129,G35130,G35131,G35132,G35133,G35134,G35135,G35136,G35137,G35138,G35139,G35140,
       G35141,G35142,G35143,G35144,G35145,G35146,G35147,G35148,G35149,G35150,G35151,G35152,G35153,G35154,G35155,G35156,G35157,G35158,G35159,G35160,
       G35161,G35162,G35163,G35164,G35165,G35166,G35167,G35168,G35169,G35170,G35171,G35172,G35173,G35174,G35175,G35176,G35177,G35178,G35179,G35180,
       G35181,G35182,G35183,G35184,G35185,G35186,G35187,G35188,G35189,G35190,G35191,G35192,G35193,G35194,G35195,G35196,G35197,G35198,G35199,G35200,
       G35201,G35202,G35203,G35204,G35205,G35206,G35207,G35208,G35209,G35210,G35211,G35212,G35213,G35214,G35215,G35216,G35217,G35218,G35219,G35220,
       G35221,G35222,G35223,G35224,G35225,G35226,G35227,G35228,G35229,G35230,G35231,G35232,G35233,G35234,G35235,G35236,G35237,G35238,G35239,G35240,
       G35241,G35242,G35243,G35244,G35245,G35246,G35247,G35248,G35249,G35250,G35251,G35252,G35253,G35254,G35255,G35256,G35257,G35258,G35259,G35260,
       G35261,G35262,G35263,G35264,G35265,G35266,G35267,G35268,G35269,G35270,G35271,G35272,G35273,G35274,G35275,G35276,G35277,G35278,G35279,G35280,
       G35281,G35282,G35283,G35284,G35285,G35286,G35287,G35288,G35289,G35290,G35291,G35292,G35293,G35294,G35295,G35296,G35297,G35298,G35299,G35300,
       G35301,G35302,G35303,G35304,G35305,G35306,G35307,G35308,G35309,G35310,G35311,G35312,G35313,G35314,G35315,G35316,G35317,G35318,G35319,G35320,
       G35321,G35322,G35323,G35324,G35325,G35326,G35327,G35328,G35329,G35330,G35331,G35332,G35333,G35334,G35335,G35336,G35337,G35338,G35339,G35340,
       G35341,G35342,G35343,G35344,G35345,G35346,G35347,G35348,G35349,G35350,G35351,G35352,G35353,G35354,G35355,G35356,G35357,G35358,G35359,G35360,
       G35361,G35362,G35363,G35364,G35365,G35366,G35367,G35368,G35369,G35370,G35371,G35372,G35373,G35374,G35375,G35376,G35377,G35378,G35379,G35380,
       G35381,G35382,G35383,G35384,G35385,G35386,G35387,G35388,G35389,G35390,G35391,G35392,G35393,G35394,G35395,G35396,G35397,G35398,G35399,G35400,
       G35401,G35402,G35403,G35404,G35405,G35406,G35407,G35408,G35409,G35410,G35411,G35412,G35413,G35414,G35415,G35416,G35417,G35418,G35419,G35420,
       G35421,G35422,G35423,G35424,G35425,G35426,G35427,G35428,G35429,G35430,G35431,G35432,G35433,G35434,G35435,G35436,G35437,G35438,G35439,G35440,
       G35441,G35442,G35443,G35444,G35445,G35446,G35447,G35448,G35449,G35450,G35451,G35452,G35453,G35454,G35455,G35456,G35457,G35458,G35459,G35460,
       G35461,G35462,G35463,G35464,G35465,G35466,G35467,G35468,G35469,G35470,G35471,G35472,G35473,G35474,G35475,G35476,G35477,G35478,G35479,G35480,
       G35481,G35482,G35483,G35484,G35485,G35486,G35487,G35488,G35489,G35490,G35491,G35492,G35493,G35494,G35495,G35496,G35497,G35498,G35499,G35500,
       G35501,G35502,G35503,G35504,G35505,G35506,G35507,G35508,G35509,G35510,G35511,G35512,G35513,G35514,G35515,G35516,G35517,G35518,G35519,G35520,
       G35521,G35522,G35523,G35524,G35525,G35526,G35527,G35528,G35529,G35530,G35531,G35532,G35533,G35534,G35535,G35536,G35537,G35538,G35539,G35540,
       G35541,G35542,G35543,G35544,G35545,G35546,G35547,G35548,G35549,G35550,G35551,G35552,G35553,G35554,G35555,G35556,G35557,G35558,G35559,G35560,
       G35561,G35562,G35563,G35564,G35565,G35566,G35567,G35568,G35569,G35570,G35571,G35572,G35573,G35574,G35575,G35576,G35577,G35578,G35579,G35580,
       G35581,G35582,G35583,G35584,G35585,G35586,G35587,G35588,G35589,G35590,G35591,G35592,G35593,G35594,G35595,G35596,G35597,G35598,G35599,G35600,
       G35601,G35602,G35603,G35604,G35605,G35606,G35607,G35608,G35609,G35610,G35611,G35612,G35613,G35614,G35615,G35616,G35617,G35618,G35619,G35620,
       G35621,G35622,G35623,G35624,G35625,G35626,G35627,G35628,G35629,G35630,G35631,G35632,G35633,G35634,G35635,G35636,G35637,G35638,G35639,G35640,
       G35641,G35642,G35643,G35644,G35645,G35646,G35647,G35648,G35649,G35650,G35651,G35652,G35653,G35654,G35655,G35656,G35657,G35658,G35659,G35660,
       G35661,G35662,G35663,G35664,G35665,G35666,G35667,G35668,G35669,G35670,G35671,G35672,G35673,G35674,G35675,G35676,G35677,G35678,G35679,G35680,
       G35681,G35682,G35683,G35684,G35685,G35686,G35687,G35688,G35689,G35690,G35691,G35692,G35693,G35694,G35695,G35696,G35697,G35698,G35699,G35700,
       G35701,G35702,G35703,G35704,G35705,G35706,G35707,G35708,G35709,G35710,G35711,G35712,G35713,G35714,G35715,G35716,G35717,G35718,G35719,G35720,
       G35721,G35722,G35723,G35724,G35725,G35726,G35727,G35728,G35729,G35730,G35731,G35732,G35733,G35734,G35735,G35736,G35737,G35738,G35739,G35740,
       G35741,G35742,G35743,G35744,G35745,G35746,G35747,G35748,G35749,G35750,G35751,G35752,G35753,G35754,G35755,G35756,G35757,G35758,G35759,G35760,
       G35761,G35762,G35763,G35764,G35765,G35766,G35767,G35768,G35769,G35770,G35771,G35772,G35773,G35774,G35775,G35776,G35777,G35778,G35779,G35780,
       G35781,G35782,G35783,G35784,G35785,G35786,G35787,G35788,G35789,G35790,G35791,G35792,G35793,G35794,G35795,G35796,G35797,G35798,G35799,G35800,
       G35801,G35802,G35803,G35804,G35805,G35806,G35807,G35808,G35809,G35810,G35811,G35812,G35813,G35814,G35815,G35816,G35817,G35818,G35819,G35820,
       G35821,G35822,G35823,G35824,G35825,G35826,G35827,G35828,G35829,G35830,G35831,G35832,G35833,G35834,G35835,G35836,G35837,G35838,G35839,G35840,
       G35841,G35842,G35843,G35844,G35845,G35846,G35847,G35848,G35849,G35850,G35851,G35852,G35853,G35854,G35855,G35856,G35857,G35858,G35859,G35860,
       G35861,G35862,G35863,G35864,G35865,G35866,G35867,G35868,G35869,G35870,G35871,G35872,G35873,G35874,G35875,G35876,G35877,G35878,G35879,G35880,
       G35881,G35882,G35883,G35884,G35885,G35886,G35887,G35888,G35889,G35890,G35891,G35892,G35893,G35894,G35895,G35896,G35897,G35898,G35899,G35900,
       G35901,G35902,G35903,G35904,G35905,G35906,G35907,G35908,G35909,G35910,G35911,G35912,G35913,G35914,G35915,G35916,G35917,G35918,G35919,G35920,
       G35921,G35922,G35923,G35924,G35925,G35926,G35927,G35928,G35929,G35930,G35931,G35932,G35933,G35934,G35935,G35936,G35937,G35938,G35939,G35940,
       G35941,G35942,G35943,G35944,G35945,G35946,G35947,G35948,G35949,G35950,G35951,G35952,G35953,G35954,G35955,G35956,G35957,G35958,G35959,G35960,
       G35961,G35962,G35963,G35964,G35965,G35966,G35967,G35968,G35969,G35970,G35971,G35972,G35973,G35974,G35975,G35976,G35977,G35978,G35979,G35980,
       G35981,G35982,G35983,G35984,G35985,G35986,G35987,G35988,G35989,G35990,G35991,G35992,G35993,G35994,G35995,G35996,G35997,G35998,G35999,G36000,
       G36001,G36002,G36003,G36004,G36005,G36006,G36007,G36008,G36009,G36010,G36011,G36012,G36013,G36014,G36015,G36016,G36017,G36018,G36019,G36020,
       G36021,G36022,G36023,G36024,G36025,G36026,G36027,G36028,G36029,G36030,G36031,G36032,G36033,G36034,G36035,G36036,G36037,G36038,G36039,G36040,
       G36041,G36042,G36043,G36044,G36045,G36046,G36047,G36048,G36049,G36050,G36051,G36052,G36053,G36054,G36055,G36056,G36057,G36058,G36059,G36060,
       G36061,G36062,G36063,G36064,G36065,G36066,G36067,G36068,G36069,G36070,G36071,G36072,G36073,G36074,G36075,G36076,G36077,G36078,G36079,G36080,
       G36081,G36082,G36083,G36084,G36085,G36086,G36087,G36088,G36089,G36090,G36091,G36092,G36093,G36094,G36095,G36096,G36097,G36098,G36099,G36100,
       G36101,G36102,G36103,G36104,G36105,G36106,G36107,G36108,G36109,G36110,G36111,G36112,G36113,G36114,G36115,G36116,G36117,G36118,G36119,G36120,
       G36121,G36122,G36123,G36124,G36125,G36126,G36127,G36128,G36129,G36130,G36131,G36132,G36133,G36134,G36135,G36136,G36137,G36138,G36139,G36140,
       G36141,G36142,G36143,G36144,G36145,G36146,G36147,G36148,G36149,G36150,G36151,G36152,G36153,G36154,G36155,G36156,G36157,G36158,G36159,G36160,
       G36161,G36162,G36163,G36164,G36165,G36166,G36167,G36168,G36169,G36170,G36171,G36172,G36173,G36174,G36175,G36176,G36177,G36178,G36179,G36180,
       G36181,G36182,G36183,G36184,G36185,G36186,G36187,G36188,G36189,G36190,G36191,G36192,G36193,G36194,G36195,G36196,G36197,G36198,G36199,G36200,
       G36201,G36202,G36203,G36204,G36205,G36206,G36207,G36208,G36209,G36210,G36211,G36212,G36213,G36214,G36215,G36216,G36217,G36218,G36219,G36220,
       G36221,G36222,G36223,G36224,G36225,G36226,G36227,G36228,G36229,G36230,G36231,G36232,G36233,G36234,G36235,G36236,G36237,G36238,G36239,G36240,
       G36241,G36242,G36243,G36244,G36245,G36246,G36247,G36248,G36249,G36250,G36251,G36252,G36253,G36254,G36255,G36256,G36257,G36258,G36259,G36260,
       G36261,G36262,G36263,G36264,G36265,G36266,G36267,G36268,G36269,G36270,G36271,G36272,G36273,G36274,G36275,G36276,G36277,G36278,G36279,G36280,
       G36281,G36282,G36283,G36284,G36285,G36286,G36287,G36288,G36289,G36290,G36291,G36292,G36293,G36294,G36295,G36296,G36297,G36298,G36299,G36300,
       G36301,G36302,G36303,G36304,G36305,G36306,G36307,G36308,G36309,G36310,G36311,G36312,G36313,G36314,G36315,G36316,G36317,G36318,G36319,G36320,
       G36321,G36322,G36323,G36324,G36325,G36326,G36327,G36328,G36329,G36330,G36331,G36332,G36333,G36334,G36335,G36336,G36337,G36338,G36339,G36340,
       G36341,G36342,G36343,G36344,G36345,G36346,G36347,G36348,G36349,G36350,G36351,G36352,G36353,G36354,G36355,G36356,G36357,G36358,G36359,G36360,
       G36361,G36362,G36363,G36364,G36365,G36366,G36367,G36368,G36369,G36370,G36371,G36372,G36373,G36374,G36375,G36376,G36377,G36378,G36379,G36380,
       G36381,G36382,G36383,G36384,G36385,G36386,G36387,G36388,G36389,G36390,G36391,G36392,G36393,G36394,G36395,G36396,G36397,G36398,G36399,G36400,
       G36401,G36402,G36403,G36404,G36405,G36406,G36407,G36408,G36409,G36410,G36411,G36412,G36413,G36414,G36415,G36416,G36417,G36418,G36419,G36420,
       G36421,G36422,G36423,G36424,G36425,G36426,G36427,G36428,G36429,G36430,G36431,G36432,G36433,G36434,G36435,G36436,G36437,G36438,G36439,G36440,
       G36441,G36442,G36443,G36444,G36445,G36446,G36447,G36448,G36449,G36450,G36451,G36452,G36453,G36454,G36455,G36456,G36457,G36458,G36459,G36460,
       G36461,G36462,G36463,G36464,G36465,G36466,G36467,G36468,G36469,G36470,G36471,G36472,G36473,G36474,G36475,G36476,G36477,G36478,G36479,G36480,
       G36481,G36482,G36483,G36484,G36485,G36486,G36487,G36488,G36489,G36490,G36491,G36492,G36493,G36494,G36495,G36496,G36497,G36498,G36499,G36500,
       G36501,G36502,G36503,G36504,G36505,G36506,G36507,G36508,G36509,G36510,G36511,G36512,G36513,G36514,G36515,G36516,G36517,G36518,G36519,G36520,
       G36521,G36522,G36523,G36524,G36525,G36526,G36527,G36528,G36529,G36530,G36531,G36532,G36533,G36534,G36535,G36536,G36537,G36538,G36539,G36540,
       G36541,G36542,G36543,G36544,G36545,G36546,G36547,G36548,G36549,G36550,G36551,G36552,G36553,G36554,G36555,G36556,G36557,G36558,G36559,G36560,
       G36561,G36562,G36563,G36564,G36565,G36566,G36567,G36568,G36569,G36570,G36571,G36572,G36573,G36574,G36575,G36576,G36577,G36578,G36579,G36580,
       G36581,G36582,G36583,G36584,G36585,G36586,G36587,G36588,G36589,G36590,G36591,G36592,G36593,G36594,G36595,G36596,G36597,G36598,G36599,G36600,
       G36601,G36602,G36603,G36604,G36605,G36606,G36607,G36608,G36609,G36610,G36611,G36612,G36613,G36614,G36615,G36616,G36617,G36618,G36619,G36620,
       G36621,G36622,G36623,G36624,G36625,G36626,G36627,G36628,G36629,G36630,G36631,G36632,G36633,G36634,G36635,G36636,G36637,G36638,G36639,G36640,
       G36641,G36642,G36643,G36644,G36645,G36646,G36647,G36648,G36649,G36650,G36651,G36652,G36653,G36654,G36655,G36656,G36657,G36658,G36659,G36660,
       G36661,G36662,G36663,G36664,G36665,G36666,G36667,G36668,G36669,G36670,G36671,G36672,G36673,G36674,G36675,G36676,G36677,G36678,G36679,G36680,
       G36681,G36682,G36683,G36684,G36685,G36686,G36687,G36688,G36689,G36690,G36691,G36692,G36693,G36694,G36695,G36696,G36697,G36698,G36699,G36700,
       G36701,G36702,G36703,G36704,G36705,G36706,G36707;

  dff DFF_55(CK,G35973,G1407);
  dff DFF_56(CK,G35974,G1408);
  dff DFF_57(CK,G35975,G1409);
  dff DFF_58(CK,G35976,G1410);
  dff DFF_59(CK,G35977,G1411);
  dff DFF_60(CK,G35978,G1412);
  dff DFF_61(CK,G35979,G1413);
  dff DFF_62(CK,G35980,G1414);
  dff DFF_63(CK,G35981,G1415);
  dff DFF_64(CK,G35982,G1416);
  dff DFF_65(CK,G35983,G1417);
  dff DFF_66(CK,G35984,G1418);
  dff DFF_67(CK,G35985,G1419);
  dff DFF_68(CK,G35986,G1420);
  dff DFF_69(CK,G35987,G1421);
  dff DFF_70(CK,G35988,G1422);
  dff DFF_71(CK,G35989,G1423);
  dff DFF_72(CK,G35990,G1424);
  dff DFF_73(CK,G35991,G1425);
  dff DFF_74(CK,G35992,G1426);
  dff DFF_75(CK,G35993,G1427);
  dff DFF_76(CK,G35994,G1428);
  dff DFF_77(CK,G35995,G1429);
  dff DFF_78(CK,G35996,G1430);
  dff DFF_79(CK,G35997,G1431);
  dff DFF_80(CK,G35998,G1432);
  dff DFF_81(CK,G35999,G1433);
  dff DFF_82(CK,G36000,G1434);
  dff DFF_83(CK,G36001,G1435);
  dff DFF_84(CK,G36002,G1436);
  dff DFF_85(CK,G36003,G1437);
  dff DFF_86(CK,G36004,G1438);
  dff DFF_87(CK,G36005,G1715);
  dff DFF_88(CK,G36006,G1716);
  dff DFF_89(CK,G36007,G1439);
  dff DFF_90(CK,G36008,G1440);
  dff DFF_91(CK,G36009,G1441);
  dff DFF_92(CK,G36010,G1442);
  dff DFF_93(CK,G36011,G1443);
  dff DFF_94(CK,G36012,G1444);
  dff DFF_95(CK,G36013,G1445);
  dff DFF_96(CK,G36014,G1446);
  dff DFF_97(CK,G36015,G1447);
  dff DFF_98(CK,G36016,G1448);
  dff DFF_99(CK,G36017,G1449);
  dff DFF_100(CK,G36018,G1450);
  dff DFF_101(CK,G36019,G1451);
  dff DFF_102(CK,G36020,G1452);
  dff DFF_103(CK,G36021,G1453);
  dff DFF_104(CK,G36022,G1454);
  dff DFF_105(CK,G36023,G1455);
  dff DFF_106(CK,G36024,G1456);
  dff DFF_107(CK,G36025,G1457);
  dff DFF_108(CK,G36026,G1458);
  dff DFF_109(CK,G36027,G1459);
  dff DFF_110(CK,G36028,G1460);
  dff DFF_111(CK,G36029,G1461);
  dff DFF_112(CK,G36030,G1462);
  dff DFF_113(CK,G36031,G1463);
  dff DFF_114(CK,G36032,G1464);
  dff DFF_115(CK,G36033,G1465);
  dff DFF_116(CK,G36034,G1466);
  dff DFF_117(CK,G36035,G1467);
  dff DFF_118(CK,G36036,G1468);
  dff DFF_119(CK,G36037,G1727);
  dff DFF_120(CK,G36038,G1730);
  dff DFF_121(CK,G36039,G1733);
  dff DFF_122(CK,G36040,G1736);
  dff DFF_123(CK,G36041,G1739);
  dff DFF_124(CK,G36042,G1742);
  dff DFF_125(CK,G36043,G1745);
  dff DFF_126(CK,G36044,G1748);
  dff DFF_127(CK,G36045,G1751);
  dff DFF_128(CK,G36046,G1754);
  dff DFF_129(CK,G36047,G1757);
  dff DFF_130(CK,G36048,G1760);
  dff DFF_131(CK,G36049,G1763);
  dff DFF_132(CK,G36050,G1766);
  dff DFF_133(CK,G36051,G1769);
  dff DFF_134(CK,G36052,G1772);
  dff DFF_135(CK,G36053,G1775);
  dff DFF_136(CK,G36054,G1778);
  dff DFF_137(CK,G36055,G1781);
  dff DFF_138(CK,G36056,G1783);
  dff DFF_139(CK,G36057,G1784);
  dff DFF_140(CK,G36058,G1785);
  dff DFF_141(CK,G36059,G1786);
  dff DFF_142(CK,G36060,G1787);
  dff DFF_143(CK,G36061,G1788);
  dff DFF_144(CK,G36062,G1789);
  dff DFF_145(CK,G36063,G1790);
  dff DFF_146(CK,G36064,G1791);
  dff DFF_147(CK,G36065,G1792);
  dff DFF_148(CK,G36066,G1793);
  dff DFF_149(CK,G36067,G1794);
  dff DFF_150(CK,G36068,G1795);
  dff DFF_151(CK,G36069,G1796);
  dff DFF_152(CK,G36070,G1797);
  dff DFF_153(CK,G36071,G1798);
  dff DFF_154(CK,G36072,G1799);
  dff DFF_155(CK,G36073,G1800);
  dff DFF_156(CK,G36074,G1801);
  dff DFF_157(CK,G36075,G1802);
  dff DFF_158(CK,G36076,G1803);
  dff DFF_159(CK,G36077,G1804);
  dff DFF_160(CK,G36078,G1805);
  dff DFF_161(CK,G36079,G1806);
  dff DFF_162(CK,G36080,G1807);
  dff DFF_163(CK,G36081,G1808);
  dff DFF_164(CK,G36082,G1809);
  dff DFF_165(CK,G36083,G1810);
  dff DFF_166(CK,G36084,G1811);
  dff DFF_167(CK,G36085,G1812);
  dff DFF_168(CK,G36086,G1813);
  dff DFF_169(CK,G36087,G1814);
  dff DFF_170(CK,G36088,G1815);
  dff DFF_171(CK,G36089,G1816);
  dff DFF_172(CK,G36090,G1817);
  dff DFF_173(CK,G36091,G1818);
  dff DFF_174(CK,G36092,G1819);
  dff DFF_175(CK,G36093,G1820);
  dff DFF_176(CK,G36094,G1821);
  dff DFF_177(CK,G36095,G1822);
  dff DFF_178(CK,G36096,G1823);
  dff DFF_179(CK,G36097,G1824);
  dff DFF_180(CK,G36098,G1825);
  dff DFF_181(CK,G36099,G1826);
  dff DFF_182(CK,G36100,G1827);
  dff DFF_183(CK,G36101,G1469);
  dff DFF_184(CK,G36102,G1828);
  dff DFF_185(CK,G36103,G1470);
  dff DFF_186(CK,G36104,G1471);
  dff DFF_187(CK,G36105,G1472);
  dff DFF_188(CK,G36106,G1473);
  dff DFF_189(CK,G36107,G1474);
  dff DFF_190(CK,G36108,G1475);
  dff DFF_191(CK,G36109,G1476);
  dff DFF_192(CK,G36110,G1477);
  dff DFF_193(CK,G36111,G1478);
  dff DFF_194(CK,G36112,G1479);
  dff DFF_195(CK,G36113,G1480);
  dff DFF_196(CK,G36114,G1481);
  dff DFF_197(CK,G36115,G1482);
  dff DFF_198(CK,G36116,G1483);
  dff DFF_199(CK,G36117,G1484);
  dff DFF_200(CK,G36118,G1485);
  dff DFF_201(CK,G36119,G1486);
  dff DFF_202(CK,G36120,G1487);
  dff DFF_203(CK,G36121,G1488);
  dff DFF_204(CK,G36122,G1489);
  dff DFF_205(CK,G36123,G1490);
  dff DFF_206(CK,G36124,G1491);
  dff DFF_207(CK,G36125,G1492);
  dff DFF_208(CK,G36126,G1493);
  dff DFF_209(CK,G36127,G1494);
  dff DFF_210(CK,G36128,G1495);
  dff DFF_211(CK,G36129,G1496);
  dff DFF_212(CK,G36130,G1497);
  dff DFF_213(CK,G36131,G1498);
  dff DFF_214(CK,G36132,G1499);
  dff DFF_215(CK,G36133,G1500);
  dff DFF_216(CK,G36134,G1501);
  dff DFF_217(CK,G36135,G1502);
  dff DFF_218(CK,G36136,G1503);
  dff DFF_219(CK,G36137,G1504);
  dff DFF_220(CK,G36138,G1505);
  dff DFF_221(CK,G36139,G1506);
  dff DFF_222(CK,G36140,G1507);
  dff DFF_223(CK,G36141,G1508);
  dff DFF_224(CK,G36142,G1509);
  dff DFF_225(CK,G36143,G1510);
  dff DFF_226(CK,G36144,G1511);
  dff DFF_227(CK,G36145,G1512);
  dff DFF_228(CK,G36146,G1513);
  dff DFF_229(CK,G36147,G1514);
  dff DFF_230(CK,G36148,G1515);
  dff DFF_231(CK,G36149,G1516);
  dff DFF_232(CK,G36150,G1517);
  dff DFF_233(CK,G36151,G1518);
  dff DFF_234(CK,G36152,G1519);
  dff DFF_235(CK,G36153,G1829);
  dff DFF_236(CK,G36154,G1830);
  dff DFF_237(CK,G36155,G1831);
  dff DFF_238(CK,G36156,G1832);
  dff DFF_239(CK,G36157,G1833);
  dff DFF_240(CK,G36158,G1834);
  dff DFF_241(CK,G36159,G1835);
  dff DFF_242(CK,G36160,G1836);
  dff DFF_243(CK,G36161,G1837);
  dff DFF_244(CK,G36162,G1838);
  dff DFF_245(CK,G36163,G1839);
  dff DFF_246(CK,G36164,G1840);
  dff DFF_247(CK,G36165,G1841);
  dff DFF_248(CK,G36166,G1842);
  dff DFF_249(CK,G36167,G1843);
  dff DFF_250(CK,G36168,G1844);
  dff DFF_251(CK,G36169,G1845);
  dff DFF_252(CK,G36170,G1846);
  dff DFF_253(CK,G36171,G1847);
  dff DFF_254(CK,G36172,G1848);
  dff DFF_255(CK,G36173,G1849);
  dff DFF_256(CK,G36174,G1850);
  dff DFF_257(CK,G36175,G1851);
  dff DFF_258(CK,G36176,G1852);
  dff DFF_259(CK,G36177,G1853);
  dff DFF_260(CK,G36178,G1854);
  dff DFF_261(CK,G36179,G1855);
  dff DFF_262(CK,G36180,G1856);
  dff DFF_263(CK,G36181,G1857);
  dff DFF_264(CK,G36182,G1858);
  dff DFF_265(CK,G36183,G1859);
  dff DFF_266(CK,G36184,G1860);
  dff DFF_267(CK,G36185,G1520);
  dff DFF_268(CK,G36186,G1521);
  dff DFF_269(CK,G36187,G1522);
  dff DFF_270(CK,G36188,G1523);
  dff DFF_271(CK,G36189,G1524);
  dff DFF_272(CK,G36190,G1525);
  dff DFF_273(CK,G36191,G1526);
  dff DFF_274(CK,G36192,G1527);
  dff DFF_275(CK,G36193,G1528);
  dff DFF_276(CK,G36194,G1529);
  dff DFF_277(CK,G36195,G1530);
  dff DFF_278(CK,G36196,G1531);
  dff DFF_279(CK,G36197,G1532);
  dff DFF_280(CK,G36198,G1533);
  dff DFF_281(CK,G36199,G1534);
  dff DFF_282(CK,G36200,G1535);
  dff DFF_283(CK,G36201,G1536);
  dff DFF_284(CK,G36202,G1537);
  dff DFF_285(CK,G36203,G1538);
  dff DFF_286(CK,G36204,G1539);
  dff DFF_287(CK,G36205,G1540);
  dff DFF_288(CK,G36206,G1541);
  dff DFF_289(CK,G36207,G1542);
  dff DFF_290(CK,G36208,G1543);
  dff DFF_291(CK,G36209,G1544);
  dff DFF_292(CK,G36210,G1545);
  dff DFF_293(CK,G36211,G1546);
  dff DFF_294(CK,G36212,G1547);
  dff DFF_295(CK,G36213,G1548);
  dff DFF_296(CK,G36214,G1549);
  dff DFF_297(CK,G36215,G1406);
  dff DFF_298(CK,G36216,G1341);
  dff DFF_299(CK,G36217,G1625);
  dff DFF_300(CK,G36218,G4390);
  dff DFF_301(CK,G36219,G4391);
  dff DFF_302(CK,G36220,G4392);
  dff DFF_303(CK,G36221,G4393);
  dff DFF_304(CK,G36222,G4394);
  dff DFF_305(CK,G36223,G4395);
  dff DFF_306(CK,G36224,G4396);
  dff DFF_307(CK,G36225,G4397);
  dff DFF_308(CK,G36226,G4398);
  dff DFF_309(CK,G36227,G4399);
  dff DFF_310(CK,G36228,G4400);
  dff DFF_311(CK,G36229,G4401);
  dff DFF_312(CK,G36230,G4402);
  dff DFF_313(CK,G36231,G4403);
  dff DFF_314(CK,G36232,G4404);
  dff DFF_315(CK,G36233,G4405);
  dff DFF_316(CK,G36234,G4406);
  dff DFF_317(CK,G36235,G4407);
  dff DFF_318(CK,G36236,G4408);
  dff DFF_319(CK,G36237,G4409);
  dff DFF_320(CK,G36238,G4410);
  dff DFF_321(CK,G36239,G4411);
  dff DFF_322(CK,G36240,G4412);
  dff DFF_323(CK,G36241,G4413);
  dff DFF_324(CK,G36242,G4414);
  dff DFF_325(CK,G36243,G4415);
  dff DFF_326(CK,G36244,G4416);
  dff DFF_327(CK,G36245,G4417);
  dff DFF_328(CK,G36246,G4418);
  dff DFF_329(CK,G36247,G4419);
  dff DFF_330(CK,G36248,G4420);
  dff DFF_331(CK,G36249,G4421);
  dff DFF_332(CK,G36250,G4692);
  dff DFF_333(CK,G36251,G4693);
  dff DFF_334(CK,G36252,G4422);
  dff DFF_335(CK,G36253,G4423);
  dff DFF_336(CK,G36254,G4424);
  dff DFF_337(CK,G36255,G4425);
  dff DFF_338(CK,G36256,G4426);
  dff DFF_339(CK,G36257,G4427);
  dff DFF_340(CK,G36258,G4428);
  dff DFF_341(CK,G36259,G4429);
  dff DFF_342(CK,G36260,G4430);
  dff DFF_343(CK,G36261,G4431);
  dff DFF_344(CK,G36262,G4432);
  dff DFF_345(CK,G36263,G4433);
  dff DFF_346(CK,G36264,G4434);
  dff DFF_347(CK,G36265,G4435);
  dff DFF_348(CK,G36266,G4436);
  dff DFF_349(CK,G36267,G4437);
  dff DFF_350(CK,G36268,G4438);
  dff DFF_351(CK,G36269,G4439);
  dff DFF_352(CK,G36270,G4440);
  dff DFF_353(CK,G36271,G4441);
  dff DFF_354(CK,G36272,G4442);
  dff DFF_355(CK,G36273,G4443);
  dff DFF_356(CK,G36274,G4444);
  dff DFF_357(CK,G36275,G4445);
  dff DFF_358(CK,G36276,G4446);
  dff DFF_359(CK,G36277,G4447);
  dff DFF_360(CK,G36278,G4448);
  dff DFF_361(CK,G36279,G4449);
  dff DFF_362(CK,G36280,G4450);
  dff DFF_363(CK,G36281,G4451);
  dff DFF_364(CK,G36282,G4704);
  dff DFF_365(CK,G36283,G4707);
  dff DFF_366(CK,G36284,G4710);
  dff DFF_367(CK,G36285,G4713);
  dff DFF_368(CK,G36286,G4716);
  dff DFF_369(CK,G36287,G4719);
  dff DFF_370(CK,G36288,G4722);
  dff DFF_371(CK,G36289,G4725);
  dff DFF_372(CK,G36290,G4728);
  dff DFF_373(CK,G36291,G4731);
  dff DFF_374(CK,G36292,G4734);
  dff DFF_375(CK,G36293,G4737);
  dff DFF_376(CK,G36294,G4740);
  dff DFF_377(CK,G36295,G4743);
  dff DFF_378(CK,G36296,G4746);
  dff DFF_379(CK,G36297,G4749);
  dff DFF_380(CK,G36298,G4752);
  dff DFF_381(CK,G36299,G4755);
  dff DFF_382(CK,G36300,G4758);
  dff DFF_383(CK,G36301,G4760);
  dff DFF_384(CK,G36302,G4761);
  dff DFF_385(CK,G36303,G4762);
  dff DFF_386(CK,G36304,G4763);
  dff DFF_387(CK,G36305,G4764);
  dff DFF_388(CK,G36306,G4765);
  dff DFF_389(CK,G36307,G4766);
  dff DFF_390(CK,G36308,G4767);
  dff DFF_391(CK,G36309,G4768);
  dff DFF_392(CK,G36310,G4769);
  dff DFF_393(CK,G36311,G4770);
  dff DFF_394(CK,G36312,G4771);
  dff DFF_395(CK,G36313,G4772);
  dff DFF_396(CK,G36314,G4773);
  dff DFF_397(CK,G36315,G4774);
  dff DFF_398(CK,G36316,G4775);
  dff DFF_399(CK,G36317,G4776);
  dff DFF_400(CK,G36318,G4777);
  dff DFF_401(CK,G36319,G4778);
  dff DFF_402(CK,G36320,G4779);
  dff DFF_403(CK,G36321,G4780);
  dff DFF_404(CK,G36322,G4781);
  dff DFF_405(CK,G36323,G4782);
  dff DFF_406(CK,G36324,G4783);
  dff DFF_407(CK,G36325,G4784);
  dff DFF_408(CK,G36326,G4785);
  dff DFF_409(CK,G36327,G4786);
  dff DFF_410(CK,G36328,G4787);
  dff DFF_411(CK,G36329,G4788);
  dff DFF_412(CK,G36330,G4789);
  dff DFF_413(CK,G36331,G4790);
  dff DFF_414(CK,G36332,G4791);
  dff DFF_415(CK,G36333,G4792);
  dff DFF_416(CK,G36334,G4793);
  dff DFF_417(CK,G36335,G4794);
  dff DFF_418(CK,G36336,G4795);
  dff DFF_419(CK,G36337,G4796);
  dff DFF_420(CK,G36338,G4797);
  dff DFF_421(CK,G36339,G4798);
  dff DFF_422(CK,G36340,G4799);
  dff DFF_423(CK,G36341,G4800);
  dff DFF_424(CK,G36342,G4801);
  dff DFF_425(CK,G36343,G4802);
  dff DFF_426(CK,G36344,G4803);
  dff DFF_427(CK,G36345,G4804);
  dff DFF_428(CK,G36346,G4452);
  dff DFF_429(CK,G36347,G4453);
  dff DFF_430(CK,G36348,G4454);
  dff DFF_431(CK,G36349,G4455);
  dff DFF_432(CK,G36350,G4456);
  dff DFF_433(CK,G36351,G4457);
  dff DFF_434(CK,G36352,G4458);
  dff DFF_435(CK,G36353,G4459);
  dff DFF_436(CK,G36354,G4460);
  dff DFF_437(CK,G36355,G4461);
  dff DFF_438(CK,G36356,G4462);
  dff DFF_439(CK,G36357,G4463);
  dff DFF_440(CK,G36358,G4464);
  dff DFF_441(CK,G36359,G4465);
  dff DFF_442(CK,G36360,G4466);
  dff DFF_443(CK,G36361,G4467);
  dff DFF_444(CK,G36362,G4468);
  dff DFF_445(CK,G36363,G4469);
  dff DFF_446(CK,G36364,G4470);
  dff DFF_447(CK,G36365,G4471);
  dff DFF_448(CK,G36366,G4472);
  dff DFF_449(CK,G36367,G4473);
  dff DFF_450(CK,G36368,G4474);
  dff DFF_451(CK,G36369,G4475);
  dff DFF_452(CK,G36370,G4476);
  dff DFF_453(CK,G36371,G4477);
  dff DFF_454(CK,G36372,G4478);
  dff DFF_455(CK,G36373,G4479);
  dff DFF_456(CK,G36374,G4480);
  dff DFF_457(CK,G36375,G4481);
  dff DFF_458(CK,G36376,G4482);
  dff DFF_459(CK,G36377,G4483);
  dff DFF_460(CK,G36378,G4484);
  dff DFF_461(CK,G36379,G4485);
  dff DFF_462(CK,G36380,G4486);
  dff DFF_463(CK,G36381,G4487);
  dff DFF_464(CK,G36382,G4488);
  dff DFF_465(CK,G36383,G4489);
  dff DFF_466(CK,G36384,G4490);
  dff DFF_467(CK,G36385,G4491);
  dff DFF_468(CK,G36386,G4492);
  dff DFF_469(CK,G36387,G4493);
  dff DFF_470(CK,G36388,G4494);
  dff DFF_471(CK,G36389,G4495);
  dff DFF_472(CK,G36390,G4496);
  dff DFF_473(CK,G36391,G4497);
  dff DFF_474(CK,G36392,G4498);
  dff DFF_475(CK,G36393,G4499);
  dff DFF_476(CK,G36394,G4500);
  dff DFF_477(CK,G36395,G4501);
  dff DFF_478(CK,G36396,G4502);
  dff DFF_479(CK,G36397,G4503);
  dff DFF_480(CK,G36398,G4805);
  dff DFF_481(CK,G36399,G4806);
  dff DFF_482(CK,G36400,G4807);
  dff DFF_483(CK,G36401,G4808);
  dff DFF_484(CK,G36402,G4809);
  dff DFF_485(CK,G36403,G4810);
  dff DFF_486(CK,G36404,G4811);
  dff DFF_487(CK,G36405,G4812);
  dff DFF_488(CK,G36406,G4813);
  dff DFF_489(CK,G36407,G4814);
  dff DFF_490(CK,G36408,G4815);
  dff DFF_491(CK,G36409,G4816);
  dff DFF_492(CK,G36410,G4817);
  dff DFF_493(CK,G36411,G4818);
  dff DFF_494(CK,G36412,G4819);
  dff DFF_495(CK,G36413,G4820);
  dff DFF_496(CK,G36414,G4821);
  dff DFF_497(CK,G36415,G4822);
  dff DFF_498(CK,G36416,G4823);
  dff DFF_499(CK,G36417,G4824);
  dff DFF_500(CK,G36418,G4825);
  dff DFF_501(CK,G36419,G4826);
  dff DFF_502(CK,G36420,G4827);
  dff DFF_503(CK,G36421,G4828);
  dff DFF_504(CK,G36422,G4829);
  dff DFF_505(CK,G36423,G4830);
  dff DFF_506(CK,G36424,G4831);
  dff DFF_507(CK,G36425,G4832);
  dff DFF_508(CK,G36426,G4833);
  dff DFF_509(CK,G36427,G4834);
  dff DFF_510(CK,G36428,G4835);
  dff DFF_511(CK,G36429,G4836);
  dff DFF_512(CK,G36430,G4504);
  dff DFF_513(CK,G36431,G4505);
  dff DFF_514(CK,G36432,G4506);
  dff DFF_515(CK,G36433,G4507);
  dff DFF_516(CK,G36434,G4508);
  dff DFF_517(CK,G36435,G4509);
  dff DFF_518(CK,G36436,G4510);
  dff DFF_519(CK,G36437,G4511);
  dff DFF_520(CK,G36438,G4512);
  dff DFF_521(CK,G36439,G4513);
  dff DFF_522(CK,G36440,G4514);
  dff DFF_523(CK,G36441,G4515);
  dff DFF_524(CK,G36442,G4516);
  dff DFF_525(CK,G36443,G4517);
  dff DFF_526(CK,G36444,G4518);
  dff DFF_527(CK,G36445,G4519);
  dff DFF_528(CK,G36446,G4520);
  dff DFF_529(CK,G36447,G4521);
  dff DFF_530(CK,G36448,G4522);
  dff DFF_531(CK,G36449,G4523);
  dff DFF_532(CK,G36450,G4524);
  dff DFF_533(CK,G36451,G4525);
  dff DFF_534(CK,G36452,G4526);
  dff DFF_535(CK,G36453,G4527);
  dff DFF_536(CK,G36454,G4528);
  dff DFF_537(CK,G36455,G4529);
  dff DFF_538(CK,G36456,G4530);
  dff DFF_539(CK,G36457,G4531);
  dff DFF_540(CK,G36458,G4532);
  dff DFF_541(CK,G36459,G4533);
  dff DFF_542(CK,G36460,G4389);
  dff DFF_543(CK,G36461,G4388);
  dff DFF_544(CK,G36462,G4591);
  dff DFF_545(CK,G36463,G7318);
  dff DFF_546(CK,G36464,G7319);
  dff DFF_547(CK,G36465,G7320);
  dff DFF_548(CK,G36466,G7321);
  dff DFF_549(CK,G36467,G7322);
  dff DFF_550(CK,G36468,G7323);
  dff DFF_551(CK,G36469,G7324);
  dff DFF_552(CK,G36470,G7325);
  dff DFF_553(CK,G36471,G7326);
  dff DFF_554(CK,G36472,G7327);
  dff DFF_555(CK,G36473,G7328);
  dff DFF_556(CK,G36474,G7329);
  dff DFF_557(CK,G36475,G7330);
  dff DFF_558(CK,G36476,G7331);
  dff DFF_559(CK,G36477,G7332);
  dff DFF_560(CK,G36478,G7333);
  dff DFF_561(CK,G36479,G7334);
  dff DFF_562(CK,G36480,G7335);
  dff DFF_563(CK,G36481,G7336);
  dff DFF_564(CK,G36482,G7337);
  dff DFF_565(CK,G36483,G7338);
  dff DFF_566(CK,G36484,G7339);
  dff DFF_567(CK,G36485,G7340);
  dff DFF_568(CK,G36486,G7341);
  dff DFF_569(CK,G36487,G7342);
  dff DFF_570(CK,G36488,G7343);
  dff DFF_571(CK,G36489,G7344);
  dff DFF_572(CK,G36490,G7345);
  dff DFF_573(CK,G36491,G7346);
  dff DFF_574(CK,G36492,G7347);
  dff DFF_575(CK,G36493,G7348);
  dff DFF_576(CK,G36494,G7349);
  dff DFF_577(CK,G36495,G7660);
  dff DFF_578(CK,G36496,G7661);
  dff DFF_579(CK,G36497,G7350);
  dff DFF_580(CK,G36498,G7351);
  dff DFF_581(CK,G36499,G7352);
  dff DFF_582(CK,G36500,G7353);
  dff DFF_583(CK,G36501,G7354);
  dff DFF_584(CK,G36502,G7355);
  dff DFF_585(CK,G36503,G7356);
  dff DFF_586(CK,G36504,G7357);
  dff DFF_587(CK,G36505,G7358);
  dff DFF_588(CK,G36506,G7359);
  dff DFF_589(CK,G36507,G7360);
  dff DFF_590(CK,G36508,G7361);
  dff DFF_591(CK,G36509,G7362);
  dff DFF_592(CK,G36510,G7363);
  dff DFF_593(CK,G36511,G7364);
  dff DFF_594(CK,G36512,G7365);
  dff DFF_595(CK,G36513,G7366);
  dff DFF_596(CK,G36514,G7367);
  dff DFF_597(CK,G36515,G7368);
  dff DFF_598(CK,G36516,G7369);
  dff DFF_599(CK,G36517,G7370);
  dff DFF_600(CK,G36518,G7371);
  dff DFF_601(CK,G36519,G7372);
  dff DFF_602(CK,G36520,G7373);
  dff DFF_603(CK,G36521,G7374);
  dff DFF_604(CK,G36522,G7375);
  dff DFF_605(CK,G36523,G7376);
  dff DFF_606(CK,G36524,G7377);
  dff DFF_607(CK,G36525,G7378);
  dff DFF_608(CK,G36526,G7379);
  dff DFF_609(CK,G36527,G7380);
  dff DFF_610(CK,G36528,G7381);
  dff DFF_611(CK,G36529,G7382);
  dff DFF_612(CK,G36530,G7383);
  dff DFF_613(CK,G36531,G7384);
  dff DFF_614(CK,G36532,G7385);
  dff DFF_615(CK,G36533,G7386);
  dff DFF_616(CK,G36534,G7387);
  dff DFF_617(CK,G36535,G7388);
  dff DFF_618(CK,G36536,G7389);
  dff DFF_619(CK,G36537,G7390);
  dff DFF_620(CK,G36538,G7391);
  dff DFF_621(CK,G36539,G7392);
  dff DFF_622(CK,G36540,G7393);
  dff DFF_623(CK,G36541,G7394);
  dff DFF_624(CK,G36542,G7395);
  dff DFF_625(CK,G36543,G7396);
  dff DFF_626(CK,G36544,G7397);
  dff DFF_627(CK,G36545,G7398);
  dff DFF_628(CK,G36546,G7399);
  dff DFF_629(CK,G36547,G7400);
  dff DFF_630(CK,G36548,G7401);
  dff DFF_631(CK,G36549,G7402);
  dff DFF_632(CK,G36550,G7403);
  dff DFF_633(CK,G36551,G7404);
  dff DFF_634(CK,G36552,G7405);
  dff DFF_635(CK,G36553,G7406);
  dff DFF_636(CK,G36554,G7407);
  dff DFF_637(CK,G36555,G7408);
  dff DFF_638(CK,G36556,G7409);
  dff DFF_639(CK,G36557,G7410);
  dff DFF_640(CK,G36558,G7411);
  dff DFF_641(CK,G36559,G7412);
  dff DFF_642(CK,G36560,G7413);
  dff DFF_643(CK,G36561,G7414);
  dff DFF_644(CK,G36562,G7415);
  dff DFF_645(CK,G36563,G7416);
  dff DFF_646(CK,G36564,G7417);
  dff DFF_647(CK,G36565,G7418);
  dff DFF_648(CK,G36566,G7419);
  dff DFF_649(CK,G36567,G7420);
  dff DFF_650(CK,G36568,G7421);
  dff DFF_651(CK,G36569,G7422);
  dff DFF_652(CK,G36570,G7423);
  dff DFF_653(CK,G36571,G7424);
  dff DFF_654(CK,G36572,G7425);
  dff DFF_655(CK,G36573,G7426);
  dff DFF_656(CK,G36574,G7427);
  dff DFF_657(CK,G36575,G7428);
  dff DFF_658(CK,G36576,G7429);
  dff DFF_659(CK,G36577,G7430);
  dff DFF_660(CK,G36578,G7431);
  dff DFF_661(CK,G36579,G7432);
  dff DFF_662(CK,G36580,G7433);
  dff DFF_663(CK,G36581,G7434);
  dff DFF_664(CK,G36582,G7435);
  dff DFF_665(CK,G36583,G7436);
  dff DFF_666(CK,G36584,G7437);
  dff DFF_667(CK,G36585,G7438);
  dff DFF_668(CK,G36586,G7439);
  dff DFF_669(CK,G36587,G7440);
  dff DFF_670(CK,G36588,G7441);
  dff DFF_671(CK,G36589,G7442);
  dff DFF_672(CK,G36590,G7443);
  dff DFF_673(CK,G36591,G7444);
  dff DFF_674(CK,G36592,G7445);
  dff DFF_675(CK,G36593,G7446);
  dff DFF_676(CK,G36594,G7447);
  dff DFF_677(CK,G36595,G7448);
  dff DFF_678(CK,G36596,G7449);
  dff DFF_679(CK,G36597,G7450);
  dff DFF_680(CK,G36598,G7451);
  dff DFF_681(CK,G36599,G7452);
  dff DFF_682(CK,G36600,G7453);
  dff DFF_683(CK,G36601,G7454);
  dff DFF_684(CK,G36602,G7455);
  dff DFF_685(CK,G36603,G7456);
  dff DFF_686(CK,G36604,G7457);
  dff DFF_687(CK,G36605,G7458);
  dff DFF_688(CK,G36606,G7459);
  dff DFF_689(CK,G36607,G7460);
  dff DFF_690(CK,G36608,G7461);
  dff DFF_691(CK,G36609,G7462);
  dff DFF_692(CK,G36610,G7463);
  dff DFF_693(CK,G36611,G7464);
  dff DFF_694(CK,G36612,G7465);
  dff DFF_695(CK,G36613,G7466);
  dff DFF_696(CK,G36614,G7467);
  dff DFF_697(CK,G36615,G7468);
  dff DFF_698(CK,G36616,G7469);
  dff DFF_699(CK,G36617,G7470);
  dff DFF_700(CK,G36618,G7471);
  dff DFF_701(CK,G36619,G7472);
  dff DFF_702(CK,G36620,G7473);
  dff DFF_703(CK,G36621,G7474);
  dff DFF_704(CK,G36622,G7475);
  dff DFF_705(CK,G36623,G7476);
  dff DFF_706(CK,G36624,G7477);
  dff DFF_707(CK,G36625,G7478);
  dff DFF_708(CK,G36626,G7479);
  dff DFF_709(CK,G36627,G7480);
  dff DFF_710(CK,G36628,G7481);
  dff DFF_711(CK,G36629,G7482);
  dff DFF_712(CK,G36630,G7483);
  dff DFF_713(CK,G36631,G7484);
  dff DFF_714(CK,G36632,G7485);
  dff DFF_715(CK,G36633,G7486);
  dff DFF_716(CK,G36634,G7487);
  dff DFF_717(CK,G36635,G7488);
  dff DFF_718(CK,G36636,G7489);
  dff DFF_719(CK,G36637,G7490);
  dff DFF_720(CK,G36638,G7491);
  dff DFF_721(CK,G36639,G7492);
  dff DFF_722(CK,G36640,G7493);
  dff DFF_723(CK,G36641,G7494);
  dff DFF_724(CK,G36642,G7495);
  dff DFF_725(CK,G36643,G7689);
  dff DFF_726(CK,G36644,G7690);
  dff DFF_727(CK,G36645,G7691);
  dff DFF_728(CK,G36646,G7692);
  dff DFF_729(CK,G36647,G7693);
  dff DFF_730(CK,G36648,G7694);
  dff DFF_731(CK,G36649,G7695);
  dff DFF_732(CK,G36650,G7696);
  dff DFF_733(CK,G36651,G7697);
  dff DFF_734(CK,G36652,G7698);
  dff DFF_735(CK,G36653,G7699);
  dff DFF_736(CK,G36654,G7700);
  dff DFF_737(CK,G36655,G7701);
  dff DFF_738(CK,G36656,G7702);
  dff DFF_739(CK,G36657,G7703);
  dff DFF_740(CK,G36658,G7704);
  dff DFF_741(CK,G36659,G7705);
  dff DFF_742(CK,G36660,G7706);
  dff DFF_743(CK,G36661,G7707);
  dff DFF_744(CK,G36662,G7708);
  dff DFF_745(CK,G36663,G7709);
  dff DFF_746(CK,G36664,G7710);
  dff DFF_747(CK,G36665,G7711);
  dff DFF_748(CK,G36666,G7712);
  dff DFF_749(CK,G36667,G7713);
  dff DFF_750(CK,G36668,G7714);
  dff DFF_751(CK,G36669,G7715);
  dff DFF_752(CK,G36670,G7716);
  dff DFF_753(CK,G36671,G7717);
  dff DFF_754(CK,G36672,G7718);
  dff DFF_755(CK,G36673,G7719);
  dff DFF_756(CK,G36674,G7720);
  dff DFF_757(CK,G36675,G7496);
  dff DFF_758(CK,G36676,G7497);
  dff DFF_759(CK,G36677,G7498);
  dff DFF_760(CK,G36678,G7499);
  dff DFF_761(CK,G36679,G7500);
  dff DFF_762(CK,G36680,G7501);
  dff DFF_763(CK,G36681,G7502);
  dff DFF_764(CK,G36682,G7503);
  dff DFF_765(CK,G36683,G7504);
  dff DFF_766(CK,G36684,G7505);
  dff DFF_767(CK,G36685,G7506);
  dff DFF_768(CK,G36686,G7507);
  dff DFF_769(CK,G36687,G7508);
  dff DFF_770(CK,G36688,G7509);
  dff DFF_771(CK,G36689,G7510);
  dff DFF_772(CK,G36690,G7511);
  dff DFF_773(CK,G36691,G7512);
  dff DFF_774(CK,G36692,G7513);
  dff DFF_775(CK,G36693,G7514);
  dff DFF_776(CK,G36694,G7515);
  dff DFF_777(CK,G36695,G7516);
  dff DFF_778(CK,G36696,G7517);
  dff DFF_779(CK,G36697,G7518);
  dff DFF_780(CK,G36698,G7519);
  dff DFF_781(CK,G36699,G7520);
  dff DFF_782(CK,G36700,G7521);
  dff DFF_783(CK,G36701,G7522);
  dff DFF_784(CK,G36702,G7523);
  dff DFF_785(CK,G36703,G7524);
  dff DFF_786(CK,G36704,G7525);
  dff DFF_787(CK,G36705,G7317);
  dff DFF_788(CK,G36706,G7316);
  dff DFF_789(CK,G36707,G7605);
  not GNAME790(G790,G7157);
  and GNAME791(G791,G790,G7159);
  or GNAME792(G792,G926,G36706);
  or GNAME793(G793,G923,G36707);
  nand GNAME794(G794,G935,G936);
  nand GNAME795(G795,G937,G938);
  nand GNAME796(G796,G939,G940);
  nand GNAME797(G797,G941,G942);
  nand GNAME798(G798,G943,G944);
  nand GNAME799(G799,G945,G946);
  nand GNAME800(G800,G947,G948);
  nand GNAME801(G801,G949,G950);
  nand GNAME802(G802,G951,G952);
  nand GNAME803(G803,G953,G954);
  nand GNAME804(G804,G955,G956);
  nand GNAME805(G805,G957,G958);
  nand GNAME806(G806,G959,G960);
  nand GNAME807(G807,G961,G962);
  nand GNAME808(G808,G963,G964);
  nand GNAME809(G809,G965,G966);
  nand GNAME810(G810,G967,G968);
  nand GNAME811(G811,G969,G970);
  nand GNAME812(G812,G971,G972);
  nand GNAME813(G813,G973,G974);
  nand GNAME814(G814,G975,G976);
  nand GNAME815(G815,G977,G978);
  nand GNAME816(G816,G979,G980);
  nand GNAME817(G817,G981,G982);
  nand GNAME818(G818,G983,G984);
  nand GNAME819(G819,G985,G986);
  nand GNAME820(G820,G987,G988);
  nand GNAME821(G821,G989,G990);
  nand GNAME822(G822,G991,G992);
  nand GNAME823(G823,G993,G994);
  nand GNAME824(G824,G995,G996);
  nand GNAME825(G825,G997,G998);
  nand GNAME826(G826,G999,G1000);
  nand GNAME827(G827,G1001,G1002);
  nand GNAME828(G828,G1003,G1004);
  nand GNAME829(G829,G1005,G1006);
  nand GNAME830(G830,G1007,G1008);
  nand GNAME831(G831,G1009,G1010);
  nand GNAME832(G832,G1011,G1012);
  nand GNAME833(G833,G1013,G1014);
  nand GNAME834(G834,G1015,G1016);
  nand GNAME835(G835,G1017,G1018);
  nand GNAME836(G836,G1019,G1020);
  nand GNAME837(G837,G1021,G1022);
  nand GNAME838(G838,G1023,G1024);
  nand GNAME839(G839,G1025,G1026);
  nand GNAME840(G840,G1027,G1028);
  nand GNAME841(G841,G1029,G1030);
  nand GNAME842(G842,G1031,G1032);
  nand GNAME843(G843,G1033,G1034);
  nand GNAME844(G844,G1035,G1036);
  nand GNAME845(G845,G1037,G1038);
  nand GNAME846(G846,G1039,G1040);
  nand GNAME847(G847,G1041,G1042);
  nand GNAME848(G848,G1043,G1044);
  nand GNAME849(G849,G1045,G1046);
  nand GNAME850(G850,G1047,G1048);
  nand GNAME851(G851,G1049,G1050);
  nand GNAME852(G852,G1051,G1052);
  nand GNAME853(G853,G1053,G1054);
  nand GNAME854(G854,G1055,G1056);
  nand GNAME855(G855,G1057,G1058);
  nand GNAME856(G856,G1059,G1060);
  nand GNAME857(G857,G1061,G1062);
  nand GNAME858(G858,G1063,G1064);
  nand GNAME859(G859,G1065,G1066);
  nand GNAME860(G860,G1067,G1068);
  nand GNAME861(G861,G1069,G1070);
  nand GNAME862(G862,G1071,G1072);
  nand GNAME863(G863,G1073,G1074);
  nand GNAME864(G864,G1075,G1076);
  nand GNAME865(G865,G1077,G1078);
  nand GNAME866(G866,G1079,G1080);
  nand GNAME867(G867,G1081,G1082);
  nand GNAME868(G868,G1083,G1084);
  nand GNAME869(G869,G1085,G1086);
  nand GNAME870(G870,G1087,G1088);
  nand GNAME871(G871,G1089,G1090);
  nand GNAME872(G872,G1091,G1092);
  nand GNAME873(G873,G1093,G1094);
  nand GNAME874(G874,G1095,G1096);
  nand GNAME875(G875,G1097,G1098);
  nand GNAME876(G876,G1099,G1100);
  nand GNAME877(G877,G1101,G1102);
  nand GNAME878(G878,G1103,G1104);
  nand GNAME879(G879,G1105,G1106);
  nand GNAME880(G880,G1107,G1108);
  nand GNAME881(G881,G1109,G1110);
  nand GNAME882(G882,G1111,G1112);
  nand GNAME883(G883,G1113,G1114);
  nand GNAME884(G884,G1115,G1116);
  nand GNAME885(G885,G1117,G1118);
  nand GNAME886(G886,G1119,G1120);
  nand GNAME887(G887,G1121,G1122);
  nand GNAME888(G888,G1123,G1124);
  nand GNAME889(G889,G1125,G1126);
  nand GNAME890(G890,G1127,G1128);
  nand GNAME891(G891,G1129,G1130);
  nand GNAME892(G892,G1131,G1132);
  nand GNAME893(G893,G1133,G1134);
  nand GNAME894(G894,G1135,G1136);
  nand GNAME895(G895,G1137,G1138);
  nand GNAME896(G896,G1139,G1140);
  nand GNAME897(G897,G1141,G1142);
  nand GNAME898(G898,G1143,G1144);
  nand GNAME899(G899,G1145,G1146);
  nand GNAME900(G900,G1147,G1148);
  nand GNAME901(G901,G1149,G1150);
  nand GNAME902(G902,G1151,G1152);
  nand GNAME903(G903,G1153,G1154);
  nand GNAME904(G904,G1155,G1156);
  nand GNAME905(G905,G1157,G1158);
  nand GNAME906(G906,G1159,G1160);
  nand GNAME907(G907,G1161,G1162);
  nand GNAME908(G908,G1163,G1164);
  nand GNAME909(G909,G1165,G1166);
  nand GNAME910(G910,G1167,G1168);
  nand GNAME911(G911,G1169,G1170);
  nand GNAME912(G912,G1171,G1172);
  nand GNAME913(G913,G1173,G1174);
  nand GNAME914(G914,G1175,G1176);
  nand GNAME915(G915,G1177,G1178);
  nand GNAME916(G916,G1179,G1180);
  nand GNAME917(G917,G1181,G1182);
  nand GNAME918(G918,G1183,G1184);
  nand GNAME919(G919,G1185,G1186);
  nand GNAME920(G920,G1187,G1188);
  nand GNAME921(G921,G1189,G1190);
  not GNAME922(G922,G36462);
  and GNAME923(G923,G931,G932);
  not GNAME924(G924,G36216);
  not GNAME925(G925,G36461);
  and GNAME926(G926,G933,G934);
  and GNAME927(G927,G928,G929);
  nand GNAME928(G928,G924,G36623,G10360,G9932);
  nand GNAME929(G929,G925,G9933,G36378,G36133);
  not GNAME930(G930,G927);
  nand GNAME931(G931,G922,G36217);
  or GNAME932(G932,G36217,G922);
  or GNAME933(G933,G36461,G924);
  or GNAME934(G934,G36216,G925);
  nand GNAME935(G935,G930,G10815);
  nand GNAME936(G936,G927,G23);
  nand GNAME937(G937,G930,G10817);
  nand GNAME938(G938,G927,G24);
  nand GNAME939(G939,G930,G10819);
  nand GNAME940(G940,G927,G25);
  nand GNAME941(G941,G930,G10821);
  nand GNAME942(G942,G927,G26);
  nand GNAME943(G943,G930,G10823);
  nand GNAME944(G944,G927,G27);
  nand GNAME945(G945,G930,G10825);
  nand GNAME946(G946,G927,G28);
  nand GNAME947(G947,G930,G10827);
  nand GNAME948(G948,G927,G29);
  nand GNAME949(G949,G930,G10719);
  nand GNAME950(G950,G927,G1);
  nand GNAME951(G951,G930,G10830);
  nand GNAME952(G952,G927,G2);
  nand GNAME953(G953,G930,G10832);
  nand GNAME954(G954,G927,G30);
  nand GNAME955(G955,G930,G10834);
  nand GNAME956(G956,G927,G3);
  nand GNAME957(G957,G930,G10836);
  nand GNAME958(G958,G927,G4);
  nand GNAME959(G959,G930,G10838);
  nand GNAME960(G960,G927,G5);
  nand GNAME961(G961,G930,G10840);
  nand GNAME962(G962,G927,G6);
  nand GNAME963(G963,G930,G10842);
  nand GNAME964(G964,G927,G7);
  nand GNAME965(G965,G930,G10844);
  nand GNAME966(G966,G927,G8);
  nand GNAME967(G967,G930,G10846);
  nand GNAME968(G968,G927,G9);
  nand GNAME969(G969,G930,G10848);
  nand GNAME970(G970,G927,G10);
  nand GNAME971(G971,G930,G10850);
  nand GNAME972(G972,G927,G11);
  nand GNAME973(G973,G930,G10852);
  nand GNAME974(G974,G927,G12);
  nand GNAME975(G975,G930,G10783);
  nand GNAME976(G976,G927,G31);
  nand GNAME977(G977,G930,G10855);
  nand GNAME978(G978,G927,G13);
  nand GNAME979(G979,G930,G10857);
  nand GNAME980(G980,G927,G14);
  nand GNAME981(G981,G930,G10859);
  nand GNAME982(G982,G927,G15);
  nand GNAME983(G983,G930,G10861);
  nand GNAME984(G984,G927,G16);
  nand GNAME985(G985,G930,G10863);
  nand GNAME986(G986,G927,G17);
  nand GNAME987(G987,G930,G10865);
  nand GNAME988(G988,G927,G18);
  nand GNAME989(G989,G930,G10867);
  nand GNAME990(G990,G927,G19);
  nand GNAME991(G991,G930,G10869);
  nand GNAME992(G992,G927,G20);
  nand GNAME993(G993,G930,G10871);
  nand GNAME994(G994,G927,G21);
  nand GNAME995(G995,G930,G10873);
  nand GNAME996(G996,G927,G22);
  nand GNAME997(G997,G930,G10720);
  nand GNAME998(G998,G927,G32);
  nand GNAME999(G999,G930,G36162);
  nand GNAME1000(G1000,G927,G10426);
  nand GNAME1001(G1001,G930,G36161);
  nand GNAME1002(G1002,G927,G10427);
  nand GNAME1003(G1003,G930,G36160);
  nand GNAME1004(G1004,G927,G10428);
  nand GNAME1005(G1005,G930,G36159);
  nand GNAME1006(G1006,G927,G10429);
  nand GNAME1007(G1007,G930,G36158);
  nand GNAME1008(G1008,G927,G10430);
  nand GNAME1009(G1009,G930,G36157);
  nand GNAME1010(G1010,G927,G10431);
  nand GNAME1011(G1011,G930,G36156);
  nand GNAME1012(G1012,G927,G10432);
  nand GNAME1013(G1013,G930,G36184);
  nand GNAME1014(G1014,G927,G10366);
  nand GNAME1015(G1015,G930,G36183);
  nand GNAME1016(G1016,G927,G10433);
  nand GNAME1017(G1017,G930,G36155);
  nand GNAME1018(G1018,G927,G10434);
  nand GNAME1019(G1019,G930,G36182);
  nand GNAME1020(G1020,G927,G10435);
  nand GNAME1021(G1021,G930,G36181);
  nand GNAME1022(G1022,G927,G10436);
  nand GNAME1023(G1023,G930,G36180);
  nand GNAME1024(G1024,G927,G10365);
  nand GNAME1025(G1025,G930,G36179);
  nand GNAME1026(G1026,G927,G10437);
  nand GNAME1027(G1027,G930,G36178);
  nand GNAME1028(G1028,G927,G10438);
  nand GNAME1029(G1029,G930,G36177);
  nand GNAME1030(G1030,G927,G10439);
  nand GNAME1031(G1031,G930,G36176);
  nand GNAME1032(G1032,G927,G10440);
  nand GNAME1033(G1033,G930,G36175);
  nand GNAME1034(G1034,G927,G10441);
  nand GNAME1035(G1035,G930,G36174);
  nand GNAME1036(G1036,G927,G10442);
  nand GNAME1037(G1037,G930,G36173);
  nand GNAME1038(G1038,G927,G10443);
  nand GNAME1039(G1039,G930,G36154);
  nand GNAME1040(G1040,G927,G10367);
  nand GNAME1041(G1041,G930,G36172);
  nand GNAME1042(G1042,G927,G10444);
  nand GNAME1043(G1043,G930,G36171);
  nand GNAME1044(G1044,G927,G10445);
  nand GNAME1045(G1045,G930,G36170);
  nand GNAME1046(G1046,G927,G10446);
  nand GNAME1047(G1047,G930,G36169);
  nand GNAME1048(G1048,G927,G10447);
  nand GNAME1049(G1049,G930,G36168);
  nand GNAME1050(G1050,G927,G10364);
  nand GNAME1051(G1051,G930,G36167);
  nand GNAME1052(G1052,G927,G10363);
  nand GNAME1053(G1053,G930,G36166);
  nand GNAME1054(G1054,G927,G10448);
  nand GNAME1055(G1055,G930,G36165);
  nand GNAME1056(G1056,G927,G10449);
  nand GNAME1057(G1057,G930,G36164);
  nand GNAME1058(G1058,G927,G10362);
  nand GNAME1059(G1059,G930,G36163);
  nand GNAME1060(G1060,G927,G10361);
  nand GNAME1061(G1061,G930,G36153);
  nand GNAME1062(G1062,G927,G10425);
  nand GNAME1063(G1063,G930,G10426);
  nand GNAME1064(G1064,G927,G36407);
  nand GNAME1065(G1065,G930,G10427);
  nand GNAME1066(G1066,G927,G36406);
  nand GNAME1067(G1067,G930,G10428);
  nand GNAME1068(G1068,G927,G36405);
  nand GNAME1069(G1069,G930,G10429);
  nand GNAME1070(G1070,G927,G36404);
  nand GNAME1071(G1071,G930,G10430);
  nand GNAME1072(G1072,G927,G36403);
  nand GNAME1073(G1073,G930,G10431);
  nand GNAME1074(G1074,G927,G36402);
  nand GNAME1075(G1075,G930,G10432);
  nand GNAME1076(G1076,G927,G36401);
  nand GNAME1077(G1077,G930,G10366);
  nand GNAME1078(G1078,G927,G36429);
  nand GNAME1079(G1079,G930,G10433);
  nand GNAME1080(G1080,G927,G36428);
  nand GNAME1081(G1081,G930,G10434);
  nand GNAME1082(G1082,G927,G36400);
  nand GNAME1083(G1083,G930,G10435);
  nand GNAME1084(G1084,G927,G36427);
  nand GNAME1085(G1085,G930,G10436);
  nand GNAME1086(G1086,G927,G36426);
  nand GNAME1087(G1087,G930,G10365);
  nand GNAME1088(G1088,G927,G36425);
  nand GNAME1089(G1089,G930,G10437);
  nand GNAME1090(G1090,G927,G36424);
  nand GNAME1091(G1091,G930,G10438);
  nand GNAME1092(G1092,G927,G36423);
  nand GNAME1093(G1093,G930,G10439);
  nand GNAME1094(G1094,G927,G36422);
  nand GNAME1095(G1095,G930,G10440);
  nand GNAME1096(G1096,G927,G36421);
  nand GNAME1097(G1097,G930,G10441);
  nand GNAME1098(G1098,G927,G36420);
  nand GNAME1099(G1099,G930,G10442);
  nand GNAME1100(G1100,G927,G36419);
  nand GNAME1101(G1101,G930,G10443);
  nand GNAME1102(G1102,G927,G36418);
  nand GNAME1103(G1103,G930,G10367);
  nand GNAME1104(G1104,G927,G36399);
  nand GNAME1105(G1105,G930,G10444);
  nand GNAME1106(G1106,G927,G36417);
  nand GNAME1107(G1107,G930,G10445);
  nand GNAME1108(G1108,G927,G36416);
  nand GNAME1109(G1109,G930,G10446);
  nand GNAME1110(G1110,G927,G36415);
  nand GNAME1111(G1111,G930,G10447);
  nand GNAME1112(G1112,G927,G36414);
  nand GNAME1113(G1113,G930,G10364);
  nand GNAME1114(G1114,G927,G36413);
  nand GNAME1115(G1115,G930,G10363);
  nand GNAME1116(G1116,G927,G36412);
  nand GNAME1117(G1117,G930,G10448);
  nand GNAME1118(G1118,G927,G36411);
  nand GNAME1119(G1119,G930,G10449);
  nand GNAME1120(G1120,G927,G36410);
  nand GNAME1121(G1121,G930,G10362);
  nand GNAME1122(G1122,G927,G36409);
  nand GNAME1123(G1123,G930,G10361);
  nand GNAME1124(G1124,G927,G36408);
  nand GNAME1125(G1125,G930,G10425);
  nand GNAME1126(G1126,G927,G36398);
  nand GNAME1127(G1127,G930,G36407);
  nand GNAME1128(G1128,G927,G36162);
  nand GNAME1129(G1129,G930,G36406);
  nand GNAME1130(G1130,G927,G36161);
  nand GNAME1131(G1131,G930,G36405);
  nand GNAME1132(G1132,G927,G36160);
  nand GNAME1133(G1133,G930,G36404);
  nand GNAME1134(G1134,G927,G36159);
  nand GNAME1135(G1135,G930,G36403);
  nand GNAME1136(G1136,G927,G36158);
  nand GNAME1137(G1137,G930,G36402);
  nand GNAME1138(G1138,G927,G36157);
  nand GNAME1139(G1139,G930,G36429);
  nand GNAME1140(G1140,G927,G36184);
  nand GNAME1141(G1141,G930,G36428);
  nand GNAME1142(G1142,G927,G36183);
  nand GNAME1143(G1143,G930,G36401);
  nand GNAME1144(G1144,G927,G36156);
  nand GNAME1145(G1145,G930,G36427);
  nand GNAME1146(G1146,G927,G36182);
  nand GNAME1147(G1147,G930,G36426);
  nand GNAME1148(G1148,G927,G36181);
  nand GNAME1149(G1149,G930,G36425);
  nand GNAME1150(G1150,G927,G36180);
  nand GNAME1151(G1151,G930,G36424);
  nand GNAME1152(G1152,G927,G36179);
  nand GNAME1153(G1153,G930,G36423);
  nand GNAME1154(G1154,G927,G36178);
  nand GNAME1155(G1155,G930,G36422);
  nand GNAME1156(G1156,G927,G36177);
  nand GNAME1157(G1157,G930,G36421);
  nand GNAME1158(G1158,G927,G36176);
  nand GNAME1159(G1159,G930,G36420);
  nand GNAME1160(G1160,G927,G36175);
  nand GNAME1161(G1161,G930,G36419);
  nand GNAME1162(G1162,G927,G36174);
  nand GNAME1163(G1163,G930,G36418);
  nand GNAME1164(G1164,G927,G36173);
  nand GNAME1165(G1165,G930,G36400);
  nand GNAME1166(G1166,G927,G36155);
  nand GNAME1167(G1167,G930,G36417);
  nand GNAME1168(G1168,G927,G36172);
  nand GNAME1169(G1169,G930,G36416);
  nand GNAME1170(G1170,G927,G36171);
  nand GNAME1171(G1171,G930,G36415);
  nand GNAME1172(G1172,G927,G36170);
  nand GNAME1173(G1173,G930,G36414);
  nand GNAME1174(G1174,G927,G36169);
  nand GNAME1175(G1175,G930,G36413);
  nand GNAME1176(G1176,G927,G36168);
  nand GNAME1177(G1177,G930,G36412);
  nand GNAME1178(G1178,G927,G36167);
  nand GNAME1179(G1179,G930,G36411);
  nand GNAME1180(G1180,G927,G36166);
  nand GNAME1181(G1181,G930,G36410);
  nand GNAME1182(G1182,G927,G36165);
  nand GNAME1183(G1183,G930,G36409);
  nand GNAME1184(G1184,G927,G36164);
  nand GNAME1185(G1185,G930,G36408);
  nand GNAME1186(G1186,G927,G36163);
  nand GNAME1187(G1187,G930,G36399);
  nand GNAME1188(G1188,G927,G36154);
  nand GNAME1189(G1189,G930,G36398);
  nand GNAME1190(G1190,G927,G36153);
  nand GNAME1191(G1191,G15024,G7747);
  nand GNAME1192(G1192,G1193,G1195,G1194);
  or GNAME1193(G1193,G7747,G15024);
  or GNAME1194(G1194,G7578,G15023);
  nand GNAME1195(G1195,G1196,G1198,G1197);
  nand GNAME1196(G1196,G15023,G7578);
  or GNAME1197(G1197,G7750,G15022);
  nand GNAME1198(G1198,G1199,G1201,G1200);
  nand GNAME1199(G1199,G15022,G7750);
  or GNAME1200(G1200,G7574,G15021);
  nand GNAME1201(G1201,G1202,G1204,G1203);
  nand GNAME1202(G1202,G15021,G7574);
  or GNAME1203(G1203,G7752,G15020);
  nand GNAME1204(G1204,G1205,G1207,G1206);
  nand GNAME1205(G1205,G15020,G7752);
  or GNAME1206(G1206,G7572,G15019);
  nand GNAME1207(G1207,G1208,G4164,G4163);
  nand GNAME1208(G1208,G15019,G7572);
  or GNAME1209(G1209,G1680,G1714);
  or GNAME1210(G1210,G1211,G1714);
  nand GNAME1211(G1211,G3191,G3192,G3190,G2032,G3189);
  nand GNAME1212(G1212,G3197,G2032,G3196);
  nand GNAME1213(G1213,G3199,G2032,G3198);
  nand GNAME1214(G1214,G3201,G2032,G3200);
  nand GNAME1215(G1215,G3203,G2032,G3202);
  nand GNAME1216(G1216,G3205,G2032,G3204);
  nand GNAME1217(G1217,G3207,G2032,G3206);
  nand GNAME1218(G1218,G3209,G2032,G3208);
  nand GNAME1219(G1219,G3211,G2032,G3210);
  nand GNAME1220(G1220,G3213,G2032,G3212);
  nand GNAME1221(G1221,G3218,G2032,G3217);
  nand GNAME1222(G1222,G3221,G3219,G3220);
  nand GNAME1223(G1223,G3224,G3222,G3223);
  nand GNAME1224(G1224,G3227,G3225,G3226);
  nand GNAME1225(G1225,G3230,G3228,G3229);
  nand GNAME1226(G1226,G3233,G3231,G3232);
  nand GNAME1227(G1227,G3236,G3234,G3235);
  nand GNAME1228(G1228,G3239,G3237,G3238);
  nand GNAME1229(G1229,G3242,G3240,G3241);
  nand GNAME1230(G1230,G3245,G3243,G3244);
  nand GNAME1231(G1231,G3171,G3169,G3170);
  nand GNAME1232(G1232,G3174,G3172,G3173);
  nand GNAME1233(G1233,G3177,G3175,G3176);
  nand GNAME1234(G1234,G3180,G3178,G3179);
  nand GNAME1235(G1235,G3183,G3181,G3182);
  nand GNAME1236(G1236,G3186,G3184,G3185);
  nand GNAME1237(G1237,G3195,G3193,G3194);
  nand GNAME1238(G1238,G3216,G3214,G3215);
  nand GNAME1239(G1239,G3248,G3246,G3247);
  nand GNAME1240(G1240,G3249,G3250,G3251,G3252);
  nand GNAME1241(G1241,G3530,G1711);
  nand GNAME1242(G1242,G2458,G2456,G2457);
  nand GNAME1243(G1243,G3531,G1711);
  nand GNAME1244(G1244,G2445,G2443,G2444);
  nand GNAME1245(G1245,G3536,G1711);
  nand GNAME1246(G1246,G1710,G3537,G3538);
  nand GNAME1247(G1247,G1710,G3539,G3540);
  nand GNAME1248(G1248,G1710,G3541,G3542);
  nand GNAME1249(G1249,G1710,G3543,G3544);
  nand GNAME1250(G1250,G1710,G3545,G3546);
  nand GNAME1251(G1251,G1710,G3547,G3548);
  nand GNAME1252(G1252,G1710,G3549,G3550);
  nand GNAME1253(G1253,G1710,G3551,G3552);
  nand GNAME1254(G1254,G1710,G3553,G3554);
  nand GNAME1255(G1255,G1710,G3559,G3560);
  nand GNAME1256(G1256,G3561,G3562,G3563,G3564);
  nand GNAME1257(G1257,G3565,G3566,G3567,G3568);
  nand GNAME1258(G1258,G3569,G3570,G3571,G3572);
  nand GNAME1259(G1259,G3573,G3574,G3575,G3576);
  nand GNAME1260(G1260,G3577,G3578,G3579,G3580);
  nand GNAME1261(G1261,G3581,G3582,G3583,G3584);
  nand GNAME1262(G1262,G3585,G3586,G3587,G3588);
  nand GNAME1263(G1263,G3589,G3590,G3591,G3592);
  nand GNAME1264(G1264,G3593,G3594,G3595,G3596);
  nand GNAME1265(G1265,G3500,G3501,G3502,G3503);
  nand GNAME1266(G1266,G3504,G3505,G3506,G3507);
  nand GNAME1267(G1267,G3508,G3509,G3510,G3511);
  nand GNAME1268(G1268,G3512,G3513,G3514,G3515);
  nand GNAME1269(G1269,G3516,G3517,G3518,G3519);
  nand GNAME1270(G1270,G3520,G3521,G3522,G3523);
  nand GNAME1271(G1271,G3532,G3533,G3534,G3535);
  nand GNAME1272(G1272,G3555,G3556,G3557,G3558);
  nand GNAME1273(G1273,G3597,G3598,G3599,G3600);
  nand GNAME1274(G1274,G3604,G3605,G3603,G3601,G3602);
  nand GNAME1275(G1275,G3624,G1626);
  nand GNAME1276(G1276,G1693,G2033,G1714,G4117,G4118);
  nand GNAME1277(G1277,G3407,G3405,G3406);
  nand GNAME1278(G1278,G3410,G3408,G3409);
  nand GNAME1279(G1279,G3414,G3415,G3416,G1696);
  nand GNAME1280(G1280,G3417,G3418,G3419,G1696);
  nand GNAME1281(G1281,G3420,G3421,G3422,G1696);
  nand GNAME1282(G1282,G3423,G3424,G3425,G1696);
  nand GNAME1283(G1283,G3426,G3427,G3428,G1696);
  nand GNAME1284(G1284,G3429,G3430,G3431,G1696);
  nand GNAME1285(G1285,G3432,G3433,G3434,G1696);
  nand GNAME1286(G1286,G3435,G3436,G3437,G1696);
  nand GNAME1287(G1287,G3438,G3439,G3440,G1696);
  nand GNAME1288(G1288,G3441,G3442,G3443,G1696);
  nand GNAME1289(G1289,G3447,G3448,G3449,G1696);
  nand GNAME1290(G1290,G3450,G3451,G3452,G1696);
  nand GNAME1291(G1291,G3453,G3454,G3455,G1696);
  nand GNAME1292(G1292,G3456,G3457,G3458,G1696);
  nand GNAME1293(G1293,G3459,G3460,G3461,G1696);
  nand GNAME1294(G1294,G3462,G3463,G3464,G1696);
  nand GNAME1295(G1295,G3465,G3466,G3467,G1696);
  nand GNAME1296(G1296,G3468,G3469,G3470,G1696);
  nand GNAME1297(G1297,G3471,G3472,G3473,G1696);
  nand GNAME1298(G1298,G3474,G3475,G3476,G1696);
  nand GNAME1299(G1299,G3387,G3388,G3389,G1696);
  nand GNAME1300(G1300,G3390,G3391,G3392,G1696);
  nand GNAME1301(G1301,G3393,G3394,G3395,G1696);
  nand GNAME1302(G1302,G3396,G3397,G3398,G1696);
  nand GNAME1303(G1303,G3399,G3400,G3401,G1696);
  nand GNAME1304(G1304,G3402,G3403,G3404,G1696);
  nand GNAME1305(G1305,G3411,G3412,G3413,G1696);
  nand GNAME1306(G1306,G3444,G3445,G3446,G1696);
  nand GNAME1307(G1307,G3477,G3478,G3479,G1696);
  nand GNAME1308(G1308,G3480,G3481,G3482,G1696);
  nand GNAME1309(G1309,G3285,G3283,G3284);
  nand GNAME1310(G1310,G3288,G3286,G3287);
  nand GNAME1311(G1311,G3293,G3294,G3295,G3296);
  nand GNAME1312(G1312,G3297,G3298,G3299,G3300);
  nand GNAME1313(G1313,G3301,G3302,G3303,G3304);
  nand GNAME1314(G1314,G3305,G3306,G3307,G3308);
  nand GNAME1315(G1315,G3309,G3310,G3311,G3312);
  nand GNAME1316(G1316,G3313,G3314,G3315,G3316);
  nand GNAME1317(G1317,G3317,G3318,G3319,G3320);
  nand GNAME1318(G1318,G3321,G3322,G3323,G3324);
  nand GNAME1319(G1319,G3325,G3326,G3327,G3328);
  nand GNAME1320(G1320,G3329,G3330,G3331,G3332);
  nand GNAME1321(G1321,G3337,G3338,G3339,G3340);
  nand GNAME1322(G1322,G3341,G3342,G3343,G3344);
  nand GNAME1323(G1323,G3345,G3346,G3347,G3348);
  nand GNAME1324(G1324,G3349,G3350,G3351,G3352);
  nand GNAME1325(G1325,G3353,G3354,G3355,G3356);
  nand GNAME1326(G1326,G3357,G3358,G3359,G3360);
  nand GNAME1327(G1327,G3361,G3362,G3363,G3364);
  nand GNAME1328(G1328,G3365,G3366,G3367,G3368);
  nand GNAME1329(G1329,G3369,G3370,G3371,G3372);
  nand GNAME1330(G1330,G3373,G3374,G3375,G3376);
  nand GNAME1331(G1331,G3259,G3260,G3261,G3262);
  nand GNAME1332(G1332,G3263,G3264,G3265,G3266);
  nand GNAME1333(G1333,G3267,G3268,G3269,G3270);
  nand GNAME1334(G1334,G3271,G3272,G3273,G3274);
  nand GNAME1335(G1335,G3275,G3276,G3277,G3278);
  nand GNAME1336(G1336,G3279,G3280,G3281,G3282);
  nand GNAME1337(G1337,G3289,G3290,G3291,G3292);
  nand GNAME1338(G1338,G3333,G3334,G3335,G3336);
  nand GNAME1339(G1339,G3377,G3378,G3379,G3380);
  nand GNAME1340(G1340,G3383,G3381,G3382);
  nand GNAME1341(G1341,G36215,G2693);
  nand GNAME1342(G1342,G3494,G1705);
  nand GNAME1343(G1343,G1705,G3495,G3646);
  nand GNAME1344(G1344,G3496,G1705);
  and GNAME1345(G1345,G3497,G1587);
  and GNAME1346(G1346,G3497,G1586);
  and GNAME1347(G1347,G3497,G1585);
  and GNAME1348(G1348,G3497,G1584);
  and GNAME1349(G1349,G3497,G1583);
  and GNAME1350(G1350,G3497,G1582);
  and GNAME1351(G1351,G3497,G1581);
  and GNAME1352(G1352,G3497,G1580);
  and GNAME1353(G1353,G3497,G1579);
  and GNAME1354(G1354,G3490,G1782);
  and GNAME1355(G1355,G3490,G1780);
  and GNAME1356(G1356,G3490,G1777);
  and GNAME1357(G1357,G3490,G1774);
  and GNAME1358(G1358,G3490,G1771);
  and GNAME1359(G1359,G3490,G1768);
  and GNAME1360(G1360,G3490,G1765);
  and GNAME1361(G1361,G3490,G1762);
  and GNAME1362(G1362,G3490,G1759);
  and GNAME1363(G1363,G3490,G1756);
  and GNAME1364(G1364,G3490,G1753);
  and GNAME1365(G1365,G3490,G1750);
  and GNAME1366(G1366,G3490,G1747);
  and GNAME1367(G1367,G3490,G1744);
  and GNAME1368(G1368,G3490,G1741);
  and GNAME1369(G1369,G3490,G1738);
  and GNAME1370(G1370,G3490,G1735);
  and GNAME1371(G1371,G3490,G1732);
  and GNAME1372(G1372,G3490,G1729);
  and GNAME1373(G1373,G3490,G1724);
  nand GNAME1374(G1374,G3487,G1702);
  nand GNAME1375(G1375,G3488,G1702);
  nand GNAME1376(G1376,G3489,G1702);
  and GNAME1377(G1377,G1647,G3484);
  and GNAME1378(G1378,G1646,G3484);
  and GNAME1379(G1379,G1649,G3484);
  and GNAME1380(G1380,G1642,G3484);
  and GNAME1381(G1381,G1639,G3484);
  and GNAME1382(G1382,G1643,G3484);
  and GNAME1383(G1383,G1645,G3484);
  and GNAME1384(G1384,G1640,G3484);
  and GNAME1385(G1385,G1644,G3484);
  and GNAME1386(G1386,G1656,G3484);
  and GNAME1387(G1387,G1657,G3484);
  and GNAME1388(G1388,G1655,G3484);
  and GNAME1389(G1389,G1653,G3484);
  and GNAME1390(G1390,G1648,G3484);
  and GNAME1391(G1391,G1651,G3484);
  and GNAME1392(G1392,G1652,G3484);
  and GNAME1393(G1393,G1654,G3484);
  and GNAME1394(G1394,G1650,G3484);
  and GNAME1395(G1395,G1637,G3484);
  and GNAME1396(G1396,G1638,G3484);
  and GNAME1397(G1397,G1630,G3484);
  and GNAME1398(G1398,G1635,G3484);
  and GNAME1399(G1399,G1634,G3484);
  and GNAME1400(G1400,G1636,G3484);
  and GNAME1401(G1401,G1632,G3484);
  and GNAME1402(G1402,G1629,G3484);
  and GNAME1403(G1403,G1633,G3484);
  and GNAME1404(G1404,G1631,G3484);
  and GNAME1405(G1405,G1658,G3484);
  not GNAME1406(G1406,G36215);
  nand GNAME1407(G1407,G2042,G2040,G2041);
  nand GNAME1408(G1408,G2045,G2043,G2044);
  nand GNAME1409(G1409,G2048,G2046,G2047);
  nand GNAME1410(G1410,G2051,G2049,G2050);
  nand GNAME1411(G1411,G2054,G2052,G2053);
  nand GNAME1412(G1412,G2057,G2055,G2056);
  nand GNAME1413(G1413,G2060,G2058,G2059);
  nand GNAME1414(G1414,G2063,G2061,G2062);
  nand GNAME1415(G1415,G2066,G2064,G2065);
  nand GNAME1416(G1416,G2069,G2067,G2068);
  nand GNAME1417(G1417,G2072,G2070,G2071);
  nand GNAME1418(G1418,G2075,G2073,G2074);
  nand GNAME1419(G1419,G2078,G2076,G2077);
  nand GNAME1420(G1420,G2081,G2079,G2080);
  nand GNAME1421(G1421,G2084,G2082,G2083);
  nand GNAME1422(G1422,G2087,G2085,G2086);
  nand GNAME1423(G1423,G2090,G2088,G2089);
  nand GNAME1424(G1424,G2093,G2091,G2092);
  nand GNAME1425(G1425,G2096,G2094,G2095);
  nand GNAME1426(G1426,G2099,G2097,G2098);
  nand GNAME1427(G1427,G2102,G2100,G2101);
  nand GNAME1428(G1428,G2105,G2103,G2104);
  nand GNAME1429(G1429,G2108,G2106,G2107);
  nand GNAME1430(G1430,G2111,G2109,G2110);
  nand GNAME1431(G1431,G2114,G2112,G2113);
  nand GNAME1432(G1432,G2117,G2115,G2116);
  nand GNAME1433(G1433,G2120,G2118,G2119);
  nand GNAME1434(G1434,G2123,G2121,G2122);
  nand GNAME1435(G1435,G2126,G2124,G2125);
  nand GNAME1436(G1436,G2129,G2127,G2128);
  nand GNAME1437(G1437,G2132,G2130,G2131);
  nand GNAME1438(G1438,G2135,G2133,G2134);
  and GNAME1439(G1439,G1989,G36007);
  and GNAME1440(G1440,G1989,G36008);
  and GNAME1441(G1441,G1989,G36009);
  and GNAME1442(G1442,G1989,G36010);
  and GNAME1443(G1443,G1989,G36011);
  and GNAME1444(G1444,G1989,G36012);
  and GNAME1445(G1445,G1989,G36013);
  and GNAME1446(G1446,G1989,G36014);
  and GNAME1447(G1447,G1989,G36015);
  and GNAME1448(G1448,G1989,G36016);
  and GNAME1449(G1449,G1989,G36017);
  and GNAME1450(G1450,G1989,G36018);
  and GNAME1451(G1451,G1989,G36019);
  and GNAME1452(G1452,G1989,G36020);
  and GNAME1453(G1453,G1989,G36021);
  and GNAME1454(G1454,G1989,G36022);
  and GNAME1455(G1455,G1989,G36023);
  and GNAME1456(G1456,G1989,G36024);
  and GNAME1457(G1457,G1989,G36025);
  and GNAME1458(G1458,G1989,G36026);
  and GNAME1459(G1459,G1989,G36027);
  and GNAME1460(G1460,G1989,G36028);
  and GNAME1461(G1461,G1989,G36029);
  and GNAME1462(G1462,G1989,G36030);
  and GNAME1463(G1463,G1989,G36031);
  and GNAME1464(G1464,G1989,G36032);
  and GNAME1465(G1465,G1989,G36033);
  and GNAME1466(G1466,G1989,G36034);
  and GNAME1467(G1467,G1989,G36035);
  and GNAME1468(G1468,G1989,G36036);
  nand GNAME1469(G1469,G1922,G2479,G2477,G2478);
  nand GNAME1470(G1470,G1923,G2492,G2490,G2491);
  nand GNAME1471(G1471,G1924,G2499,G2497,G2498);
  nand GNAME1472(G1472,G1925,G2503,G2504,G2505);
  nand GNAME1473(G1473,G1926,G2510,G2511,G2512);
  nand GNAME1474(G1474,G1927,G2517,G2518,G2519);
  nand GNAME1475(G1475,G1928,G2524,G2525,G2526);
  nand GNAME1476(G1476,G1929,G2531,G2532,G2533);
  nand GNAME1477(G1477,G1930,G2538,G2539,G2540);
  nand GNAME1478(G1478,G1931,G2545,G2546,G2547);
  nand GNAME1479(G1479,G1932,G2552,G2553,G2554);
  nand GNAME1480(G1480,G1933,G2559,G2560,G2561);
  nand GNAME1481(G1481,G1934,G2566,G2567,G2568);
  nand GNAME1482(G1482,G1935,G2573,G2574,G2575);
  nand GNAME1483(G1483,G1936,G2580,G2581,G2582);
  nand GNAME1484(G1484,G1937,G2587,G2588,G2589);
  nand GNAME1485(G1485,G1938,G2594,G2595,G2596);
  nand GNAME1486(G1486,G1939,G2601,G2602,G2603);
  nand GNAME1487(G1487,G1940,G2608,G2609,G2610);
  nand GNAME1488(G1488,G1941,G2615,G2616,G2617);
  nand GNAME1489(G1489,G1942,G2622,G2623,G2624);
  nand GNAME1490(G1490,G1943,G2629,G2630,G2631);
  nand GNAME1491(G1491,G1944,G2636,G2637,G2638);
  nand GNAME1492(G1492,G1945,G2643,G2644,G2645);
  nand GNAME1493(G1493,G1946,G2650,G2651,G2652);
  nand GNAME1494(G1494,G1947,G2657,G2658,G2659);
  nand GNAME1495(G1495,G1948,G2664,G2665,G2666);
  nand GNAME1496(G1496,G1949,G2671,G2672,G2673);
  nand GNAME1497(G1497,G2678,G1993,G2677,G2675,G2676);
  nand GNAME1498(G1498,G2681,G3878,G3879);
  nand GNAME1499(G1499,G2684,G3880,G3881);
  nand GNAME1500(G1500,G2699,G2700,G3106,G2697,G2698);
  nand GNAME1501(G1501,G2707,G2708,G2706,G2705,G2917);
  nand GNAME1502(G1502,G2715,G2716,G2714,G2713,G3016);
  nand GNAME1503(G1503,G2723,G2724,G2722,G2721,G3036);
  nand GNAME1504(G1504,G2731,G2732,G2730,G2729,G2885);
  nand GNAME1505(G1505,G2739,G2740,G2738,G2737,G3146);
  nand GNAME1506(G1506,G2747,G2748,G2746,G2745,G2957);
  nand GNAME1507(G1507,G2755,G2756,G2754,G2753,G3056);
  nand GNAME1508(G1508,G2763,G2764,G2762,G2761,G2937);
  nand GNAME1509(G1509,G2771,G2772,G2770,G2769,G3126);
  nand GNAME1510(G1510,G2779,G2780,G2778,G2777,G2986);
  nand GNAME1511(G1511,G2787,G2788,G2786,G2785,G3086);
  nand GNAME1512(G1512,G2795,G2796,G2794,G2793,G3166);
  nand GNAME1513(G1513,G2803,G2804,G2802,G2801,G2907);
  nand GNAME1514(G1514,G2811,G2812,G2810,G2809,G3026);
  nand GNAME1515(G1515,G1950,G2817,G2818,G2819);
  nand GNAME1516(G1516,G2827,G2828,G2826,G2825,G3116);
  nand GNAME1517(G1517,G1951,G2833,G2834,G2835);
  nand GNAME1518(G1518,G2843,G2844,G2842,G2841,G3076);
  nand GNAME1519(G1519,G2851,G2852,G2850,G2849,G2976);
  nand GNAME1520(G1520,G2868,G2866,G2867);
  nand GNAME1521(G1521,G1959,G2882,G2880,G2883);
  nand GNAME1522(G1522,G1960,G2894,G2895,G2896);
  nand GNAME1523(G1523,G1961,G2904,G2905,G2903);
  nand GNAME1524(G1524,G1962,G2914,G2912,G2915);
  nand GNAME1525(G1525,G1963,G2924,G2922,G2923);
  nand GNAME1526(G1526,G1964,G2934,G2935,G2933);
  nand GNAME1527(G1527,G1965,G2944,G2945,G2946);
  nand GNAME1528(G1528,G1966,G2954,G2955,G2953);
  nand GNAME1529(G1529,G1967,G2964,G2965,G2966);
  nand GNAME1530(G1530,G1968,G2973,G2971,G2972);
  nand GNAME1531(G1531,G1969,G2983,G2984,G2982);
  nand GNAME1532(G1532,G1970,G2993,G2991,G2992);
  nand GNAME1533(G1533,G1971,G3003,G3004,G3005);
  nand GNAME1534(G1534,G1972,G3013,G3011,G3014);
  nand GNAME1535(G1535,G1973,G3023,G3024,G3022);
  nand GNAME1536(G1536,G1974,G3033,G3031,G3034);
  nand GNAME1537(G1537,G1975,G3043,G3044,G3045);
  nand GNAME1538(G1538,G1976,G3053,G3054,G3052);
  nand GNAME1539(G1539,G1977,G3063,G3064,G3065);
  nand GNAME1540(G1540,G1978,G3073,G3071,G3072);
  nand GNAME1541(G1541,G1979,G3083,G3084,G3082);
  nand GNAME1542(G1542,G1980,G3093,G3094,G3095);
  nand GNAME1543(G1543,G1981,G3103,G3101,G3104);
  nand GNAME1544(G1544,G1982,G3113,G3111,G3112);
  nand GNAME1545(G1545,G1983,G3123,G3124,G3122);
  nand GNAME1546(G1546,G1984,G3133,G3134,G3135);
  nand GNAME1547(G1547,G1985,G3143,G3144,G3142);
  nand GNAME1548(G1548,G1986,G3153,G3154,G3155);
  nand GNAME1549(G1549,G1987,G3163,G3164,G3162);
  nor GNAME1550(G1550,G1406,G1551);
  and GNAME1551(G1551,G36215,G1988);
  not GNAME1552(G1552,G11997);
  not GNAME1553(G1553,G36002);
  not GNAME1554(G1554,G36003);
  nand GNAME1555(G1555,G3617,G1713);
  or GNAME1556(G1556,G2137,G1714);
  nand GNAME1557(G1557,G1712,G3617);
  not GNAME1558(G1558,G36185);
  nor GNAME1559(G1559,G1406,G1556);
  nand GNAME1560(G1560,G3617,G3620,G3621);
  nor GNAME1561(G1561,G3652,G1718);
  and GNAME1562(G1562,G3665,G3668);
  nand GNAME1563(G1563,G3655,G1562);
  and GNAME1564(G1564,G1994,G2144);
  and GNAME1565(G1565,G1718,G1719);
  and GNAME1566(G1566,G3643,G1565);
  and GNAME1567(G1567,G3655,G3649);
  nand GNAME1568(G1568,G3646,G1567);
  and GNAME1569(G1569,G3655,G1719);
  and GNAME1570(G1570,G3652,G1569);
  and GNAME1571(G1571,G3652,G1718,G3655);
  and GNAME1572(G1572,G2149,G2006);
  nor GNAME1573(G1573,G3655,G1720);
  and GNAME1574(G1574,G1572,G2007,G1604);
  not GNAME1575(G1575,G36101);
  not GNAME1576(G1576,G36069);
  and GNAME1577(G1577,G1717,G1565);
  and GNAME1578(G1578,G2167,G2168);
  and GNAME1579(G1579,G2016,G877);
  and GNAME1580(G1580,G2016,G876);
  and GNAME1581(G1581,G2016,G875);
  and GNAME1582(G1582,G2016,G874);
  and GNAME1583(G1583,G2016,G873);
  and GNAME1584(G1584,G2016,G872);
  and GNAME1585(G1585,G2016,G871);
  and GNAME1586(G1586,G2016,G870);
  and GNAME1587(G1587,G2016,G869);
  and GNAME1588(G1588,G2016,G868);
  and GNAME1589(G1589,G3652,G3646,G3649);
  and GNAME1590(G1590,G2016,G866);
  and GNAME1591(G1591,G2016,G865);
  and GNAME1592(G1592,G1725,G3668);
  nand GNAME1593(G1593,G3655,G1592);
  and GNAME1594(G1594,G1726,G3665);
  nand GNAME1595(G1595,G3649,G1721,G3646);
  nand GNAME1596(G1596,G2470,G1559);
  and GNAME1597(G1597,G1566,G2029);
  and GNAME1598(G1598,G1612,G2029);
  and GNAME1599(G1599,G2473,G2029);
  or GNAME1600(G1600,G1720,G1595);
  nor GNAME1601(G1601,G1596,G1600);
  and GNAME1602(G1602,G3649,G1720,G1721);
  nor GNAME1603(G1603,G2471,G1596);
  nand GNAME1604(G1604,G1718,G1720);
  and GNAME1605(G1605,G2007,G1667,G1604);
  and GNAME1606(G1606,G1719,G1721);
  and GNAME1607(G1607,G1577,G2029);
  or GNAME1608(G1608,G1720,G1568);
  or GNAME1609(G1609,G1712,G1555);
  nor GNAME1610(G1610,G1717,G1406,G2694);
  and GNAME1611(G1611,G1714,G1721);
  nand GNAME1612(G1612,G2033,G1608);
  nand GNAME1613(G1613,G2013,G2012);
  and GNAME1614(G1614,G1616,G2686);
  and GNAME1615(G1615,G1617,G2686);
  or GNAME1616(G1616,G1613,G2011,G1612);
  or GNAME1617(G1617,G4160,G1571,G1570);
  and GNAME1618(G1618,G2685,G3643);
  and GNAME1619(G1619,G1622,G1559);
  and GNAME1620(G1620,G1717,G1723);
  and GNAME1621(G1621,G2696,G36215,G1622);
  or GNAME1622(G1622,G1341,G1624);
  and GNAME1623(G1623,G1714,G1610);
  and GNAME1624(G1624,G3624,G2137);
  and GNAME1625(G1625,G36215,G1624);
  and GNAME1626(G1626,G1719,G1571);
  and GNAME1627(G1627,G1620,G1626);
  and GNAME1628(G1628,G1714,G1719);
  nand GNAME1629(G1629,G2173,G2174,G2175,G2176);
  nand GNAME1630(G1630,G2223,G2224,G2225,G2226);
  nand GNAME1631(G1631,G2145,G2146,G2147,G2148);
  nand GNAME1632(G1632,G2183,G2184,G2185,G2186);
  nand GNAME1633(G1633,G2159,G2160,G2161,G2162);
  nand GNAME1634(G1634,G2203,G2204,G2205,G2206);
  nand GNAME1635(G1635,G2213,G2214,G2215,G2216);
  nand GNAME1636(G1636,G2193,G2194,G2195,G2196);
  nand GNAME1637(G1637,G2243,G2244,G2245,G2246);
  nand GNAME1638(G1638,G2233,G2234,G2235,G2236);
  nand GNAME1639(G1639,G2383,G2384,G2385,G2386);
  nand GNAME1640(G1640,G2353,G2354,G2355,G2356);
  nand GNAME1641(G1641,G2433,G2434,G2435,G2436);
  nand GNAME1642(G1642,G2393,G2394,G2395,G2396);
  nand GNAME1643(G1643,G2373,G2374,G2375,G2376);
  nand GNAME1644(G1644,G2343,G2344,G2345,G2346);
  nand GNAME1645(G1645,G2363,G2364,G2365,G2366);
  nand GNAME1646(G1646,G2413,G2414,G2415,G2416);
  nand GNAME1647(G1647,G2423,G2424,G2425,G2426);
  nand GNAME1648(G1648,G2293,G2294,G2295,G2296);
  nand GNAME1649(G1649,G2403,G2404,G2405,G2406);
  nand GNAME1650(G1650,G2253,G2254,G2255,G2256);
  nand GNAME1651(G1651,G2283,G2284,G2285,G2286);
  nand GNAME1652(G1652,G2273,G2274,G2275,G2276);
  nand GNAME1653(G1653,G2303,G2304,G2305,G2306);
  nand GNAME1654(G1654,G2263,G2264,G2265,G2266);
  nand GNAME1655(G1655,G2313,G2314,G2315,G2316);
  nand GNAME1656(G1656,G2333,G2334,G2335,G2336);
  nand GNAME1657(G1657,G2323,G2324,G2325,G2326);
  nand GNAME1658(G1658,G2163,G2164,G2165,G2166);
  and GNAME1659(G1659,G1955,G1956,G1954,G1952,G1953);
  and GNAME1660(G1660,G1957,G1958);
  nor GNAME1661(G1661,G1721,G1998);
  and GNAME1662(G1662,G1714,G1567);
  not GNAME1663(G1663,G11853);
  nor GNAME1664(G1664,G3668,G3665);
  and GNAME1665(G1665,G1613,G1559);
  nand GNAME1666(G1666,G1564,G1664);
  nand GNAME1667(G1667,G1718,G1573);
  and GNAME1668(G1668,G1720,G1569);
  nand GNAME1669(G1669,G2874,G1608);
  nand GNAME1670(G1670,G2008,G1685,G2873,G1572);
  and GNAME1671(G1671,G2879,G2025,G2878);
  and GNAME1672(G1672,G1559,G2017);
  and GNAME1673(G1673,G1669,G1672);
  and GNAME1674(G1674,G1670,G1672);
  nor GNAME1675(G1675,G3643,G1666);
  nor GNAME1676(G1676,G1717,G1666);
  nor GNAME1677(G1677,G2137,G1275,G1406);
  and GNAME1678(G1678,G2891,G1559);
  and GNAME1679(G1679,G1609,G1570);
  nor GNAME1680(G1680,G1556,G1604);
  and GNAME1681(G1681,G1721,G1680);
  and GNAME1682(G1682,G3655,G1664);
  and GNAME1683(G1683,G1609,G1571);
  nor GNAME1684(G1684,G2137,G3646);
  or GNAME1685(G1685,G1718,G2007);
  nor GNAME1686(G1686,G2137,G1685);
  and GNAME1687(G1687,G1573,G1664);
  nand GNAME1688(G1688,G1996,G1997,G2003,G2004);
  nand GNAME1689(G1689,G2038,G2039,G2037,G2000,G2001);
  nor GNAME1690(G1690,G1695,G4159);
  and GNAME1691(G1691,G3257,G1595);
  and GNAME1692(G1692,G2006,G1568,G1667,G3253);
  nand GNAME1693(G1693,G1720,G1567);
  nor GNAME1694(G1694,G4159,G1693);
  nor GNAME1695(G1695,G1602,G1668);
  and GNAME1696(G1696,G2009,G1714);
  and GNAME1697(G1697,G2024,G2019,G2020);
  and GNAME1698(G1698,G3483,G2018,G2023);
  nand GNAME1699(G1699,G2022,G4161);
  nand GNAME1700(G1700,G1697,G1698);
  nor GNAME1701(G1701,G1699,G1700);
  and GNAME1702(G1702,G3485,G3486);
  nand GNAME1703(G1703,G1563,G2021,G1593);
  nor GNAME1704(G1704,G1682,G1703);
  and GNAME1705(G1705,G3492,G3493);
  and GNAME1706(G1706,G3608,G1609,G3660);
  and GNAME1707(G1707,G1723,G1609,G3608);
  or GNAME1708(G1708,G1628,G1611,G1662);
  nand GNAME1709(G1709,G2035,G2036,G2002,G1995,G1999);
  and GNAME1710(G1710,G3524,G3525);
  and GNAME1711(G1711,G3529,G1710,G3528,G3526,G3527);
  and GNAME1712(G1712,G3613,G3614);
  nand GNAME1713(G1713,G3618,G3619);
  nand GNAME1714(G1714,G3622,G3623);
  nand GNAME1715(G1715,G3625,G3626);
  nand GNAME1716(G1716,G3627,G3628);
  nand GNAME1717(G1717,G3641,G3642);
  nand GNAME1718(G1718,G3644,G3645);
  nand GNAME1719(G1719,G3647,G3648);
  nand GNAME1720(G1720,G3650,G3651);
  nand GNAME1721(G1721,G3653,G3654);
  nand GNAME1722(G1722,G3656,G3657);
  nand GNAME1723(G1723,G3658,G3659);
  nand GNAME1724(G1724,G3661,G3662);
  nand GNAME1725(G1725,G3663,G3664);
  nand GNAME1726(G1726,G3666,G3667);
  nand GNAME1727(G1727,G3672,G3673);
  nand GNAME1728(G1728,G3674,G3675);
  nand GNAME1729(G1729,G3676,G3677);
  nand GNAME1730(G1730,G3678,G3679);
  nand GNAME1731(G1731,G3680,G3681);
  nand GNAME1732(G1732,G3682,G3683);
  nand GNAME1733(G1733,G3684,G3685);
  nand GNAME1734(G1734,G3686,G3687);
  nand GNAME1735(G1735,G3688,G3689);
  nand GNAME1736(G1736,G3690,G3691);
  nand GNAME1737(G1737,G3692,G3693);
  nand GNAME1738(G1738,G3694,G3695);
  nand GNAME1739(G1739,G3696,G3697);
  nand GNAME1740(G1740,G3698,G3699);
  nand GNAME1741(G1741,G3700,G3701);
  nand GNAME1742(G1742,G3702,G3703);
  nand GNAME1743(G1743,G3704,G3705);
  nand GNAME1744(G1744,G3706,G3707);
  nand GNAME1745(G1745,G3708,G3709);
  nand GNAME1746(G1746,G3710,G3711);
  nand GNAME1747(G1747,G3712,G3713);
  nand GNAME1748(G1748,G3714,G3715);
  nand GNAME1749(G1749,G3716,G3717);
  nand GNAME1750(G1750,G3718,G3719);
  nand GNAME1751(G1751,G3720,G3721);
  nand GNAME1752(G1752,G3722,G3723);
  nand GNAME1753(G1753,G3724,G3725);
  nand GNAME1754(G1754,G3726,G3727);
  nand GNAME1755(G1755,G3728,G3729);
  nand GNAME1756(G1756,G3730,G3731);
  nand GNAME1757(G1757,G3732,G3733);
  nand GNAME1758(G1758,G3734,G3735);
  nand GNAME1759(G1759,G3736,G3737);
  nand GNAME1760(G1760,G3738,G3739);
  nand GNAME1761(G1761,G3740,G3741);
  nand GNAME1762(G1762,G3742,G3743);
  nand GNAME1763(G1763,G3744,G3745);
  nand GNAME1764(G1764,G3746,G3747);
  nand GNAME1765(G1765,G3748,G3749);
  nand GNAME1766(G1766,G3750,G3751);
  nand GNAME1767(G1767,G3752,G3753);
  nand GNAME1768(G1768,G3754,G3755);
  nand GNAME1769(G1769,G3756,G3757);
  nand GNAME1770(G1770,G3758,G3759);
  nand GNAME1771(G1771,G3760,G3761);
  nand GNAME1772(G1772,G3762,G3763);
  nand GNAME1773(G1773,G3764,G3765);
  nand GNAME1774(G1774,G3766,G3767);
  nand GNAME1775(G1775,G3768,G3769);
  nand GNAME1776(G1776,G3770,G3771);
  nand GNAME1777(G1777,G3772,G3773);
  nand GNAME1778(G1778,G3774,G3775);
  nand GNAME1779(G1779,G3776,G3777);
  nand GNAME1780(G1780,G3778,G3779);
  nand GNAME1781(G1781,G3780,G3781);
  nand GNAME1782(G1782,G3782,G3783);
  nand GNAME1783(G1783,G3784,G3785);
  nand GNAME1784(G1784,G3786,G3787);
  nand GNAME1785(G1785,G3788,G3789);
  nand GNAME1786(G1786,G3790,G3791);
  nand GNAME1787(G1787,G3792,G3793);
  nand GNAME1788(G1788,G3794,G3795);
  nand GNAME1789(G1789,G3796,G3797);
  nand GNAME1790(G1790,G3798,G3799);
  nand GNAME1791(G1791,G3800,G3801);
  nand GNAME1792(G1792,G3802,G3803);
  nand GNAME1793(G1793,G3804,G3805);
  nand GNAME1794(G1794,G3806,G3807);
  nand GNAME1795(G1795,G3808,G3809);
  nand GNAME1796(G1796,G3810,G3811);
  nand GNAME1797(G1797,G3812,G3813);
  nand GNAME1798(G1798,G3814,G3815);
  nand GNAME1799(G1799,G3816,G3817);
  nand GNAME1800(G1800,G3818,G3819);
  nand GNAME1801(G1801,G3820,G3821);
  nand GNAME1802(G1802,G3822,G3823);
  nand GNAME1803(G1803,G3824,G3825);
  nand GNAME1804(G1804,G3826,G3827);
  nand GNAME1805(G1805,G3828,G3829);
  nand GNAME1806(G1806,G3830,G3831);
  nand GNAME1807(G1807,G3832,G3833);
  nand GNAME1808(G1808,G3834,G3835);
  nand GNAME1809(G1809,G3836,G3837);
  nand GNAME1810(G1810,G3838,G3839);
  nand GNAME1811(G1811,G3840,G3841);
  nand GNAME1812(G1812,G3842,G3843);
  nand GNAME1813(G1813,G3844,G3845);
  nand GNAME1814(G1814,G3846,G3847);
  nand GNAME1815(G1815,G3848,G3849);
  nand GNAME1816(G1816,G3850,G3851);
  nand GNAME1817(G1817,G3852,G3853);
  nand GNAME1818(G1818,G3854,G3855);
  nand GNAME1819(G1819,G3856,G3857);
  nand GNAME1820(G1820,G3858,G3859);
  nand GNAME1821(G1821,G3860,G3861);
  nand GNAME1822(G1822,G3862,G3863);
  nand GNAME1823(G1823,G3864,G3865);
  nand GNAME1824(G1824,G3866,G3867);
  nand GNAME1825(G1825,G3868,G3869);
  nand GNAME1826(G1826,G3870,G3871);
  nand GNAME1827(G1827,G3872,G3873);
  nand GNAME1828(G1828,G3874,G3875);
  nand GNAME1829(G1829,G3882,G3883);
  nand GNAME1830(G1830,G3884,G3885);
  nand GNAME1831(G1831,G3886,G3887);
  nand GNAME1832(G1832,G3888,G3889);
  nand GNAME1833(G1833,G3890,G3891);
  nand GNAME1834(G1834,G3892,G3893);
  nand GNAME1835(G1835,G3894,G3895);
  nand GNAME1836(G1836,G3896,G3897);
  nand GNAME1837(G1837,G3898,G3899);
  nand GNAME1838(G1838,G3900,G3901);
  nand GNAME1839(G1839,G3902,G3903);
  nand GNAME1840(G1840,G3904,G3905);
  nand GNAME1841(G1841,G3906,G3907);
  nand GNAME1842(G1842,G3908,G3909);
  nand GNAME1843(G1843,G3910,G3911);
  nand GNAME1844(G1844,G3912,G3913);
  nand GNAME1845(G1845,G3914,G3915);
  nand GNAME1846(G1846,G3916,G3917);
  nand GNAME1847(G1847,G3918,G3919);
  nand GNAME1848(G1848,G3920,G3921);
  nand GNAME1849(G1849,G3922,G3923);
  nand GNAME1850(G1850,G3924,G3925);
  nand GNAME1851(G1851,G3926,G3927);
  nand GNAME1852(G1852,G3928,G3929);
  nand GNAME1853(G1853,G3930,G3931);
  nand GNAME1854(G1854,G3932,G3933);
  nand GNAME1855(G1855,G3934,G3935);
  nand GNAME1856(G1856,G3936,G3937);
  nand GNAME1857(G1857,G3938,G3939);
  nand GNAME1858(G1858,G3940,G3941);
  nand GNAME1859(G1859,G3942,G3943);
  nand GNAME1860(G1860,G3944,G3945);
  nand GNAME1861(G1861,G4049,G4050);
  nand GNAME1862(G1862,G4051,G4052);
  nand GNAME1863(G1863,G4053,G4054);
  nand GNAME1864(G1864,G4055,G4056);
  nand GNAME1865(G1865,G4057,G4058);
  nand GNAME1866(G1866,G4059,G4060);
  nand GNAME1867(G1867,G4061,G4062);
  nand GNAME1868(G1868,G4063,G4064);
  nand GNAME1869(G1869,G4065,G4066);
  nand GNAME1870(G1870,G4067,G4068);
  nand GNAME1871(G1871,G4069,G4070);
  nand GNAME1872(G1872,G4071,G4072);
  nand GNAME1873(G1873,G4073,G4074);
  nand GNAME1874(G1874,G4075,G4076);
  nand GNAME1875(G1875,G4077,G4078);
  nand GNAME1876(G1876,G4079,G4080);
  nand GNAME1877(G1877,G4081,G4082);
  nand GNAME1878(G1878,G4083,G4084);
  nand GNAME1879(G1879,G4085,G4086);
  nand GNAME1880(G1880,G4087,G4088);
  nand GNAME1881(G1881,G4089,G4090);
  nand GNAME1882(G1882,G4091,G4092);
  nand GNAME1883(G1883,G4093,G4094);
  nand GNAME1884(G1884,G4095,G4096);
  nand GNAME1885(G1885,G4097,G4098);
  nand GNAME1886(G1886,G4099,G4100);
  nand GNAME1887(G1887,G4101,G4102);
  nand GNAME1888(G1888,G4103,G4104);
  nand GNAME1889(G1889,G4105,G4106);
  nand GNAME1890(G1890,G4107,G4108);
  nand GNAME1891(G1891,G4109,G4110);
  nand GNAME1892(G1892,G4111,G4112);
  nand GNAME1893(G1893,G4113,G4114);
  nand GNAME1894(G1894,G4119,G4120);
  nand GNAME1895(G1895,G4121,G4122);
  nand GNAME1896(G1896,G4123,G4124);
  nand GNAME1897(G1897,G4125,G4126);
  nand GNAME1898(G1898,G4127,G4128);
  nand GNAME1899(G1899,G4129,G4130);
  nand GNAME1900(G1900,G4131,G4132);
  nand GNAME1901(G1901,G4133,G4134);
  nand GNAME1902(G1902,G4135,G4136);
  nand GNAME1903(G1903,G4137,G4138);
  nand GNAME1904(G1904,G4139,G4140);
  nand GNAME1905(G1905,G4141,G4142);
  nand GNAME1906(G1906,G4143,G4144);
  nand GNAME1907(G1907,G4145,G4146);
  nand GNAME1908(G1908,G4147,G4148);
  nand GNAME1909(G1909,G4149,G4150);
  nand GNAME1910(G1910,G4151,G4152);
  nand GNAME1911(G1911,G4153,G4154);
  nand GNAME1912(G1912,G4155,G4156);
  nand GNAME1913(G1913,G4157,G4158);
  or GNAME1914(G1914,G36033,G36034,G36035,G36036);
  nor GNAME1915(G1915,G1914,G36032,G36031,G36030,G36029);
  or GNAME1916(G1916,G36025,G36026,G36027,G36028);
  nor GNAME1917(G1917,G1916,G36022,G36024,G36023);
  or GNAME1918(G1918,G36018,G36019,G36020,G36021);
  nor GNAME1919(G1919,G1918,G36015,G36017,G36016);
  or GNAME1920(G1920,G36011,G36012,G36013,G36014);
  nor GNAME1921(G1921,G1920,G36008,G36010,G36009);
  and GNAME1922(G1922,G2476,G2474,G2475);
  and GNAME1923(G1923,G2486,G2487,G2488,G2489);
  and GNAME1924(G1924,G2493,G2494,G2495,G2496);
  and GNAME1925(G1925,G2500,G2501,G2502,G2506);
  and GNAME1926(G1926,G2507,G2508,G2509,G2513);
  and GNAME1927(G1927,G2514,G2515,G2516,G2520);
  and GNAME1928(G1928,G2521,G2522,G2523,G2527);
  and GNAME1929(G1929,G2528,G2529,G2530,G2534);
  and GNAME1930(G1930,G2535,G2536,G2537,G2541);
  and GNAME1931(G1931,G2542,G2543,G2544,G2548);
  and GNAME1932(G1932,G2549,G2550,G2551,G2555);
  and GNAME1933(G1933,G2556,G2557,G2558,G2562);
  and GNAME1934(G1934,G2563,G2564,G2565,G2569);
  and GNAME1935(G1935,G2570,G2571,G2572,G2576);
  and GNAME1936(G1936,G2577,G2578,G2579,G2583);
  and GNAME1937(G1937,G2584,G2585,G2586,G2590);
  and GNAME1938(G1938,G2591,G2592,G2593,G2597);
  and GNAME1939(G1939,G2598,G2599,G2600,G2604);
  and GNAME1940(G1940,G2605,G2606,G2607,G2611);
  and GNAME1941(G1941,G2612,G2613,G2614,G2618);
  and GNAME1942(G1942,G2619,G2620,G2621,G2625);
  and GNAME1943(G1943,G2626,G2627,G2628,G2632);
  and GNAME1944(G1944,G2633,G2634,G2635,G2639);
  and GNAME1945(G1945,G2640,G2641,G2642,G2646);
  and GNAME1946(G1946,G2647,G2648,G2649,G2653);
  and GNAME1947(G1947,G2654,G2655,G2656,G2660);
  and GNAME1948(G1948,G2661,G2662,G2663,G2667);
  and GNAME1949(G1949,G2668,G2669,G2670,G2674);
  and GNAME1950(G1950,G2996,G2034,G2820);
  and GNAME1951(G1951,G2927,G2034,G2836);
  and GNAME1952(G1952,G3978,G3981,G3984);
  and GNAME1953(G1953,G3987,G3990,G3993);
  and GNAME1954(G1954,G4005,G4008,G3996,G3999,G4002);
  and GNAME1955(G1955,G4020,G4023,G4011,G4014,G4017);
  and GNAME1956(G1956,G4035,G4038,G4026,G4029,G4032);
  and GNAME1957(G1957,G3957,G3960,G3948,G3951,G3954);
  and GNAME1958(G1958,G3972,G3975,G3963,G3966,G3969);
  and GNAME1959(G1959,G2885,G2881,G2884);
  and GNAME1960(G1960,G2897,G2892,G2893);
  and GNAME1961(G1961,G2907,G2902,G2906);
  and GNAME1962(G1962,G2917,G2913,G2916);
  and GNAME1963(G1963,G2927,G2925,G2926);
  and GNAME1964(G1964,G2937,G2932,G2936);
  and GNAME1965(G1965,G2947,G2942,G2943);
  and GNAME1966(G1966,G2957,G2952,G2956);
  and GNAME1967(G1967,G2967,G2962,G2963);
  and GNAME1968(G1968,G2976,G2974,G2975);
  and GNAME1969(G1969,G2986,G2981,G2985);
  and GNAME1970(G1970,G2996,G2994,G2995);
  and GNAME1971(G1971,G3006,G3001,G3002);
  and GNAME1972(G1972,G3016,G3012,G3015);
  and GNAME1973(G1973,G3026,G3021,G3025);
  and GNAME1974(G1974,G3036,G3032,G3035);
  and GNAME1975(G1975,G3046,G3041,G3042);
  and GNAME1976(G1976,G3056,G3051,G3055);
  and GNAME1977(G1977,G3066,G3061,G3062);
  and GNAME1978(G1978,G3076,G3074,G3075);
  and GNAME1979(G1979,G3086,G3081,G3085);
  and GNAME1980(G1980,G3096,G3091,G3092);
  and GNAME1981(G1981,G3106,G3102,G3105);
  and GNAME1982(G1982,G3116,G3114,G3115);
  and GNAME1983(G1983,G3126,G3121,G3125);
  and GNAME1984(G1984,G3136,G3131,G3132);
  and GNAME1985(G1985,G3146,G3141,G3145);
  and GNAME1986(G1986,G3156,G3151,G3152);
  and GNAME1987(G1987,G3166,G3161,G3165);
  not GNAME1988(G1988,G36004);
  nand GNAME1989(G1989,G1560,G1559);
  and GNAME1990(G1990,G3660,G3643);
  nand GNAME1991(G1991,G1564,G2142,G1559);
  nand GNAME1992(G1992,G1564,G2467,G1559);
  and GNAME1993(G1993,G3876,G3877);
  nand GNAME1994(G1994,G2143,G2136);
  nand GNAME1995(G1995,G1562,G1679);
  nand GNAME1996(G1996,G1664,G1686);
  nand GNAME1997(G1997,G1664,G1679);
  not GNAME1998(G1998,G1628);
  nand GNAME1999(G1999,G1664,G1681);
  nand GNAME2000(G2000,G1592,G1679);
  nand GNAME2001(G2001,G1594,G1679);
  nand GNAME2002(G2002,G1680,G1682);
  nand GNAME2003(G2003,G1664,G1683);
  nand GNAME2004(G2004,G1684,G1687);
  nand GNAME2005(G2005,G3660,G1714);
  nand GNAME2006(G2006,G3649,G1571);
  not GNAME2007(G2007,G1668);
  or GNAME2008(G2008,G1719,G1667);
  nand GNAME2009(G2009,G1720,G1606);
  not GNAME2010(G2010,G1608);
  not GNAME2011(G2011,G1600);
  or GNAME2012(G2012,G3652,G1568);
  nand GNAME2013(G2013,G3646,G1602);
  nand GNAME2014(G2014,G2468,G1565);
  nand GNAME2015(G2015,G1660,G1659,G4041);
  not GNAME2016(G2016,G1990);
  not GNAME2017(G2017,G1666);
  nand GNAME2018(G2018,G1561,G1592);
  nand GNAME2019(G2019,G1562,G1573);
  nand GNAME2020(G2020,G1573,G1592);
  nand GNAME2021(G2021,G3655,G1594);
  nand GNAME2022(G2022,G1561,G1664);
  nand GNAME2023(G2023,G1561,G1562);
  nand GNAME2024(G2024,G1573,G1594);
  not GNAME2025(G2025,G1625);
  not GNAME2026(G2026,G1989);
  not GNAME2027(G2027,G1991);
  not GNAME2028(G2028,G1992);
  not GNAME2029(G2029,G1596);
  nand GNAME2030(G2030,G1565,G2447,G1242);
  nand GNAME2031(G2031,G1559,G2011);
  nand GNAME2032(G2032,G3168,G1721);
  not GNAME2033(G2033,G1606);
  nand GNAME2034(G2034,G1893,G1625);
  nand GNAME2035(G2035,G1703,G1680);
  nand GNAME2036(G2036,G3609,G1681);
  nand GNAME2037(G2037,G3609,G1683);
  nand GNAME2038(G2038,G3167,G1684);
  nand GNAME2039(G2039,G3609,G1686);
  nand GNAME2040(G2040,G1406,G889);
  nand GNAME2041(G2041,G1550,G35973);
  nand GNAME2042(G2042,G1551,G35973);
  nand GNAME2043(G2043,G1406,G878);
  nand GNAME2044(G2044,G1550,G12017);
  nand GNAME2045(G2045,G1551,G35974);
  nand GNAME2046(G2046,G1406,G867);
  nand GNAME2047(G2047,G1550,G11998);
  nand GNAME2048(G2048,G1551,G35975);
  nand GNAME2049(G2049,G1406,G864);
  nand GNAME2050(G2050,G1550,G11999);
  nand GNAME2051(G2051,G1551,G35976);
  nand GNAME2052(G2052,G1406,G863);
  nand GNAME2053(G2053,G1550,G12022);
  nand GNAME2054(G2054,G1551,G35977);
  nand GNAME2055(G2055,G1406,G862);
  nand GNAME2056(G2056,G1550,G12021);
  nand GNAME2057(G2057,G1551,G35978);
  nand GNAME2058(G2058,G1406,G861);
  nand GNAME2059(G2059,G1550,G12000);
  nand GNAME2060(G2060,G1551,G35979);
  nand GNAME2061(G2061,G1406,G860);
  nand GNAME2062(G2062,G1550,G12001);
  nand GNAME2063(G2063,G1551,G35980);
  nand GNAME2064(G2064,G1406,G859);
  nand GNAME2065(G2065,G1550,G12020);
  nand GNAME2066(G2066,G1551,G35981);
  nand GNAME2067(G2067,G1406,G858);
  nand GNAME2068(G2068,G1550,G12019);
  nand GNAME2069(G2069,G1551,G35982);
  nand GNAME2070(G2070,G1406,G888);
  nand GNAME2071(G2071,G1550,G11987);
  nand GNAME2072(G2072,G1551,G35983);
  nand GNAME2073(G2073,G1406,G887);
  nand GNAME2074(G2074,G1550,G11988);
  nand GNAME2075(G2075,G1551,G35984);
  nand GNAME2076(G2076,G1406,G886);
  nand GNAME2077(G2077,G1550,G12034);
  nand GNAME2078(G2078,G1551,G35985);
  nand GNAME2079(G2079,G1406,G885);
  nand GNAME2080(G2080,G1550,G12033);
  nand GNAME2081(G2081,G1551,G35986);
  nand GNAME2082(G2082,G1406,G884);
  nand GNAME2083(G2083,G1550,G11989);
  nand GNAME2084(G2084,G1551,G35987);
  nand GNAME2085(G2085,G1406,G883);
  nand GNAME2086(G2086,G1550,G11990);
  nand GNAME2087(G2087,G1551,G35988);
  nand GNAME2088(G2088,G1406,G882);
  nand GNAME2089(G2089,G1550,G12032);
  nand GNAME2090(G2090,G1551,G35989);
  nand GNAME2091(G2091,G1406,G881);
  nand GNAME2092(G2092,G1550,G12031);
  nand GNAME2093(G2093,G1551,G35990);
  nand GNAME2094(G2094,G1406,G880);
  nand GNAME2095(G2095,G1550,G11991);
  nand GNAME2096(G2096,G1551,G35991);
  nand GNAME2097(G2097,G1406,G879);
  nand GNAME2098(G2098,G1550,G11992);
  nand GNAME2099(G2099,G1551,G35992);
  nand GNAME2100(G2100,G1406,G877);
  nand GNAME2101(G2101,G1550,G12029);
  nand GNAME2102(G2102,G1551,G35993);
  nand GNAME2103(G2103,G1406,G876);
  nand GNAME2104(G2104,G1550,G12028);
  nand GNAME2105(G2105,G1551,G35994);
  nand GNAME2106(G2106,G1406,G875);
  nand GNAME2107(G2107,G1550,G11993);
  nand GNAME2108(G2108,G1551,G35995);
  nand GNAME2109(G2109,G1406,G874);
  nand GNAME2110(G2110,G1550,G11994);
  nand GNAME2111(G2111,G1551,G35996);
  nand GNAME2112(G2112,G1406,G873);
  nand GNAME2113(G2113,G1550,G12027);
  nand GNAME2114(G2114,G1551,G35997);
  nand GNAME2115(G2115,G1406,G872);
  nand GNAME2116(G2116,G1550,G12026);
  nand GNAME2117(G2117,G1551,G35998);
  nand GNAME2118(G2118,G1406,G871);
  nand GNAME2119(G2119,G1550,G11995);
  nand GNAME2120(G2120,G1551,G35999);
  nand GNAME2121(G2121,G1406,G870);
  nand GNAME2122(G2122,G1550,G11996);
  nand GNAME2123(G2123,G1551,G36000);
  nand GNAME2124(G2124,G1406,G869);
  nand GNAME2125(G2125,G1550,G12025);
  nand GNAME2126(G2126,G1551,G36001);
  nand GNAME2127(G2127,G1406,G868);
  nand GNAME2128(G2128,G1550,G11997);
  nand GNAME2129(G2129,G1551,G36002);
  nand GNAME2130(G2130,G1406,G866);
  nand GNAME2131(G2131,G1550,G12024);
  nand GNAME2132(G2132,G1551,G36003);
  nand GNAME2133(G2133,G1406,G865);
  nand GNAME2134(G2134,G1550,G12018);
  nand GNAME2135(G2135,G1551,G36004);
  not GNAME2136(G2136,G1560);
  not GNAME2137(G2137,G1609);
  nand GNAME2138(G2138,G1557,G3618,G3619);
  nand GNAME2139(G2139,G1712,G1557);
  nand GNAME2140(G2140,G3671,G1562);
  or GNAME2141(G2141,G1720,G1563);
  nand GNAME2142(G2142,G2141,G2023,G2140);
  nand GNAME2143(G2143,G1915,G1917,G1919,G1921);
  nand GNAME2144(G2144,G36007,G2136);
  nand GNAME2145(G2145,G3631,G36205);
  nand GNAME2146(G2146,G3634,G36102);
  nand GNAME2147(G2147,G3637,G36070);
  nand GNAME2148(G2148,G3640,G36038);
  nand GNAME2149(G2149,G3646,G1570);
  nand GNAME2150(G2150,G3649,G1573);
  nand GNAME2151(G2151,G2150,G1574);
  nand GNAME2152(G2152,G2012,G1595);
  or GNAME2153(G2153,G1589,G1606);
  nand GNAME2154(G2154,G1631,G1566);
  nand GNAME2155(G2155,G2152,G1724);
  nand GNAME2156(G2156,G2153,G12212);
  nand GNAME2157(G2157,G2151,G11117);
  nand GNAME2158(G2158,G2154,G2155,G2156,G2157);
  nand GNAME2159(G2159,G3640,G36039);
  nand GNAME2160(G2160,G3631,G36190);
  nand GNAME2161(G2161,G3634,G36103);
  nand GNAME2162(G2162,G3637,G36071);
  nand GNAME2163(G2163,G3631,G36195);
  nand GNAME2164(G2164,G3634,G36101);
  nand GNAME2165(G2165,G3637,G36069);
  nand GNAME2166(G2166,G3640,G36037);
  nand GNAME2167(G2167,G1658,G1577);
  nand GNAME2168(G2168,G1633,G1566);
  nand GNAME2169(G2169,G2152,G1729);
  nand GNAME2170(G2170,G2153,G12275);
  nand GNAME2171(G2171,G2151,G11132);
  nand GNAME2172(G2172,G2169,G2170,G2171,G1578);
  nand GNAME2173(G2173,G3640,G36040);
  nand GNAME2174(G2174,G3631,G12085);
  nand GNAME2175(G2175,G3634,G36104);
  nand GNAME2176(G2176,G3637,G36072);
  nand GNAME2177(G2177,G1631,G1577);
  nand GNAME2178(G2178,G1629,G1566);
  nand GNAME2179(G2179,G2152,G1732);
  nand GNAME2180(G2180,G2153,G12324);
  nand GNAME2181(G2181,G2151,G11066);
  nand GNAME2182(G2182,G2180,G2181,G2179,G2177,G2178);
  nand GNAME2183(G2183,G3640,G36041);
  nand GNAME2184(G2184,G3631,G12129);
  nand GNAME2185(G2185,G3634,G36105);
  nand GNAME2186(G2186,G3637,G36073);
  nand GNAME2187(G2187,G1633,G1577);
  nand GNAME2188(G2188,G1632,G1566);
  nand GNAME2189(G2189,G2152,G1735);
  nand GNAME2190(G2190,G2153,G12319);
  nand GNAME2191(G2191,G2151,G11069);
  nand GNAME2192(G2192,G2190,G2191,G2189,G2187,G2188);
  nand GNAME2193(G2193,G3640,G36042);
  nand GNAME2194(G2194,G3631,G12128);
  nand GNAME2195(G2195,G3634,G36106);
  nand GNAME2196(G2196,G3637,G36074);
  nand GNAME2197(G2197,G1629,G1577);
  nand GNAME2198(G2198,G1636,G1566);
  nand GNAME2199(G2199,G2152,G1738);
  nand GNAME2200(G2200,G2153,G12317);
  nand GNAME2201(G2201,G2151,G11121);
  nand GNAME2202(G2202,G2200,G2201,G2199,G2197,G2198);
  nand GNAME2203(G2203,G3640,G36043);
  nand GNAME2204(G2204,G3631,G12127);
  nand GNAME2205(G2205,G3634,G36107);
  nand GNAME2206(G2206,G3637,G36075);
  nand GNAME2207(G2207,G1632,G1577);
  nand GNAME2208(G2208,G1634,G1566);
  nand GNAME2209(G2209,G2152,G1741);
  nand GNAME2210(G2210,G2153,G12315);
  nand GNAME2211(G2211,G2151,G11120);
  nand GNAME2212(G2212,G2210,G2211,G2209,G2207,G2208);
  nand GNAME2213(G2213,G3640,G36044);
  nand GNAME2214(G2214,G3631,G12126);
  nand GNAME2215(G2215,G3634,G36108);
  nand GNAME2216(G2216,G3637,G36076);
  nand GNAME2217(G2217,G1636,G1577);
  nand GNAME2218(G2218,G1635,G1566);
  nand GNAME2219(G2219,G2152,G1744);
  nand GNAME2220(G2220,G2153,G12313);
  nand GNAME2221(G2221,G2151,G11070);
  nand GNAME2222(G2222,G2220,G2221,G2219,G2217,G2218);
  nand GNAME2223(G2223,G3640,G36045);
  nand GNAME2224(G2224,G3631,G12125);
  nand GNAME2225(G2225,G3634,G36109);
  nand GNAME2226(G2226,G3637,G36077);
  nand GNAME2227(G2227,G1634,G1577);
  nand GNAME2228(G2228,G1630,G1566);
  nand GNAME2229(G2229,G2152,G1747);
  nand GNAME2230(G2230,G2153,G12311);
  nand GNAME2231(G2231,G2151,G11071);
  nand GNAME2232(G2232,G2230,G2231,G2229,G2227,G2228);
  nand GNAME2233(G2233,G3640,G36046);
  nand GNAME2234(G2234,G3631,G12124);
  nand GNAME2235(G2235,G3634,G36110);
  nand GNAME2236(G2236,G3637,G36078);
  nand GNAME2237(G2237,G1635,G1577);
  nand GNAME2238(G2238,G1638,G1566);
  nand GNAME2239(G2239,G2152,G1750);
  nand GNAME2240(G2240,G2153,G12309);
  nand GNAME2241(G2241,G2151,G11119);
  nand GNAME2242(G2242,G2240,G2241,G2239,G2237,G2238);
  nand GNAME2243(G2243,G3640,G36047);
  nand GNAME2244(G2244,G3631,G12148);
  nand GNAME2245(G2245,G3634,G36111);
  nand GNAME2246(G2246,G3637,G36079);
  nand GNAME2247(G2247,G1630,G1577);
  nand GNAME2248(G2248,G1637,G1566);
  nand GNAME2249(G2249,G2152,G1753);
  nand GNAME2250(G2250,G2153,G12307);
  nand GNAME2251(G2251,G2151,G11118);
  nand GNAME2252(G2252,G2250,G2251,G2249,G2247,G2248);
  nand GNAME2253(G2253,G3640,G36048);
  nand GNAME2254(G2254,G3631,G12147);
  nand GNAME2255(G2255,G3634,G36112);
  nand GNAME2256(G2256,G3637,G36080);
  nand GNAME2257(G2257,G1638,G1577);
  nand GNAME2258(G2258,G1650,G1566);
  nand GNAME2259(G2259,G2152,G1756);
  nand GNAME2260(G2260,G2153,G12365);
  nand GNAME2261(G2261,G2151,G11063);
  nand GNAME2262(G2262,G2260,G2261,G2259,G2257,G2258);
  nand GNAME2263(G2263,G3640,G36049);
  nand GNAME2264(G2264,G3631,G12146);
  nand GNAME2265(G2265,G3634,G36113);
  nand GNAME2266(G2266,G3637,G36081);
  nand GNAME2267(G2267,G1637,G1577);
  nand GNAME2268(G2268,G1654,G1566);
  nand GNAME2269(G2269,G2152,G1759);
  nand GNAME2270(G2270,G2153,G12363);
  nand GNAME2271(G2271,G2151,G11064);
  nand GNAME2272(G2272,G2270,G2271,G2269,G2267,G2268);
  nand GNAME2273(G2273,G3640,G36050);
  nand GNAME2274(G2274,G3631,G12145);
  nand GNAME2275(G2275,G3634,G36114);
  nand GNAME2276(G2276,G3637,G36082);
  nand GNAME2277(G2277,G1650,G1577);
  nand GNAME2278(G2278,G1652,G1566);
  nand GNAME2279(G2279,G2152,G1762);
  nand GNAME2280(G2280,G2153,G12361);
  nand GNAME2281(G2281,G2151,G11139);
  nand GNAME2282(G2282,G2280,G2281,G2279,G2277,G2278);
  nand GNAME2283(G2283,G3640,G36051);
  nand GNAME2284(G2284,G3631,G12144);
  nand GNAME2285(G2285,G3634,G36115);
  nand GNAME2286(G2286,G3637,G36083);
  nand GNAME2287(G2287,G1654,G1577);
  nand GNAME2288(G2288,G1651,G1566);
  nand GNAME2289(G2289,G2152,G1765);
  nand GNAME2290(G2290,G2153,G12359);
  nand GNAME2291(G2291,G2151,G11138);
  nand GNAME2292(G2292,G2290,G2291,G2289,G2287,G2288);
  nand GNAME2293(G2293,G3640,G36052);
  nand GNAME2294(G2294,G3631,G12143);
  nand GNAME2295(G2295,G3634,G36116);
  nand GNAME2296(G2296,G3637,G36084);
  nand GNAME2297(G2297,G1652,G1577);
  nand GNAME2298(G2298,G1648,G1566);
  nand GNAME2299(G2299,G2152,G1768);
  nand GNAME2300(G2300,G2153,G12357);
  nand GNAME2301(G2301,G2151,G11065);
  nand GNAME2302(G2302,G2300,G2301,G2299,G2297,G2298);
  nand GNAME2303(G2303,G3640,G36053);
  nand GNAME2304(G2304,G3631,G12142);
  nand GNAME2305(G2305,G3634,G36117);
  nand GNAME2306(G2306,G3637,G36085);
  nand GNAME2307(G2307,G1651,G1577);
  nand GNAME2308(G2308,G1653,G1566);
  nand GNAME2309(G2309,G2152,G1771);
  nand GNAME2310(G2310,G2153,G12355);
  nand GNAME2311(G2311,G2151,G11137);
  nand GNAME2312(G2312,G2310,G2311,G2309,G2307,G2308);
  nand GNAME2313(G2313,G3640,G36054);
  nand GNAME2314(G2314,G3631,G12141);
  nand GNAME2315(G2315,G3634,G36118);
  nand GNAME2316(G2316,G3637,G36086);
  nand GNAME2317(G2317,G1648,G1577);
  nand GNAME2318(G2318,G1655,G1566);
  nand GNAME2319(G2319,G2152,G1774);
  nand GNAME2320(G2320,G2153,G12353);
  nand GNAME2321(G2321,G2151,G11136);
  nand GNAME2322(G2322,G2320,G2321,G2319,G2317,G2318);
  nand GNAME2323(G2323,G3640,G36055);
  nand GNAME2324(G2324,G3631,G12140);
  nand GNAME2325(G2325,G3634,G36119);
  nand GNAME2326(G2326,G3637,G36087);
  nand GNAME2327(G2327,G1653,G1577);
  nand GNAME2328(G2328,G1657,G1566);
  nand GNAME2329(G2329,G2152,G1777);
  nand GNAME2330(G2330,G2153,G12351);
  nand GNAME2331(G2331,G2151,G11135);
  nand GNAME2332(G2332,G2330,G2331,G2329,G2327,G2328);
  nand GNAME2333(G2333,G3640,G36056);
  nand GNAME2334(G2334,G3631,G12139);
  nand GNAME2335(G2335,G3634,G36120);
  nand GNAME2336(G2336,G3637,G36088);
  nand GNAME2337(G2337,G1655,G1577);
  nand GNAME2338(G2338,G1656,G1566);
  nand GNAME2339(G2339,G2152,G1780);
  nand GNAME2340(G2340,G2153,G12349);
  nand GNAME2341(G2341,G2151,G11134);
  nand GNAME2342(G2342,G2340,G2341,G2339,G2337,G2338);
  nand GNAME2343(G2343,G3634,G36121);
  nand GNAME2344(G2344,G3637,G36089);
  nand GNAME2345(G2345,G3640,G36057);
  nand GNAME2346(G2346,G3631,G12138);
  nand GNAME2347(G2347,G1657,G1577);
  nand GNAME2348(G2348,G1644,G1566);
  nand GNAME2349(G2349,G2152,G1782);
  nand GNAME2350(G2350,G2153,G12347);
  nand GNAME2351(G2351,G2151,G11133);
  nand GNAME2352(G2352,G2350,G2351,G2349,G2347,G2348);
  nand GNAME2353(G2353,G3634,G36122);
  nand GNAME2354(G2354,G3637,G36090);
  nand GNAME2355(G2355,G3640,G36058);
  nand GNAME2356(G2356,G3631,G12137);
  nand GNAME2357(G2357,G1656,G1577);
  nand GNAME2358(G2358,G1640,G1566);
  nand GNAME2359(G2359,G2153,G12344);
  nand GNAME2360(G2360,G2152,G1579);
  nand GNAME2361(G2361,G2151,G11131);
  nand GNAME2362(G2362,G2360,G2361,G2359,G2357,G2358);
  nand GNAME2363(G2363,G3634,G36123);
  nand GNAME2364(G2364,G3637,G36091);
  nand GNAME2365(G2365,G3640,G36059);
  nand GNAME2366(G2366,G3631,G12136);
  nand GNAME2367(G2367,G1644,G1577);
  nand GNAME2368(G2368,G1645,G1566);
  nand GNAME2369(G2369,G2153,G12342);
  nand GNAME2370(G2370,G2152,G1580);
  nand GNAME2371(G2371,G2151,G11130);
  nand GNAME2372(G2372,G2370,G2371,G2369,G2367,G2368);
  nand GNAME2373(G2373,G3634,G36124);
  nand GNAME2374(G2374,G3637,G36092);
  nand GNAME2375(G2375,G3640,G36060);
  nand GNAME2376(G2376,G3631,G12135);
  nand GNAME2377(G2377,G1640,G1577);
  nand GNAME2378(G2378,G1643,G1566);
  nand GNAME2379(G2379,G2153,G12340);
  nand GNAME2380(G2380,G2152,G1581);
  nand GNAME2381(G2381,G2151,G11129);
  nand GNAME2382(G2382,G2380,G2381,G2379,G2377,G2378);
  nand GNAME2383(G2383,G3634,G36125);
  nand GNAME2384(G2384,G3637,G36093);
  nand GNAME2385(G2385,G3640,G36061);
  nand GNAME2386(G2386,G3631,G12134);
  nand GNAME2387(G2387,G1645,G1577);
  nand GNAME2388(G2388,G1639,G1566);
  nand GNAME2389(G2389,G2153,G12338);
  nand GNAME2390(G2390,G2152,G1582);
  nand GNAME2391(G2391,G2151,G11128);
  nand GNAME2392(G2392,G2390,G2391,G2389,G2387,G2388);
  nand GNAME2393(G2393,G3634,G36126);
  nand GNAME2394(G2394,G3637,G36094);
  nand GNAME2395(G2395,G3640,G36062);
  nand GNAME2396(G2396,G3631,G12133);
  nand GNAME2397(G2397,G1643,G1577);
  nand GNAME2398(G2398,G1642,G1566);
  nand GNAME2399(G2399,G2153,G12336);
  nand GNAME2400(G2400,G2152,G1583);
  nand GNAME2401(G2401,G2151,G11127);
  nand GNAME2402(G2402,G2400,G2401,G2399,G2397,G2398);
  nand GNAME2403(G2403,G3634,G36127);
  nand GNAME2404(G2404,G3637,G36095);
  nand GNAME2405(G2405,G3640,G36063);
  nand GNAME2406(G2406,G3631,G12132);
  nand GNAME2407(G2407,G1639,G1577);
  nand GNAME2408(G2408,G1649,G1566);
  nand GNAME2409(G2409,G2153,G12334);
  nand GNAME2410(G2410,G2152,G1584);
  nand GNAME2411(G2411,G2151,G11126);
  nand GNAME2412(G2412,G2410,G2411,G2409,G2407,G2408);
  nand GNAME2413(G2413,G3634,G36128);
  nand GNAME2414(G2414,G3637,G36096);
  nand GNAME2415(G2415,G3640,G36064);
  nand GNAME2416(G2416,G3631,G12131);
  nand GNAME2417(G2417,G1642,G1577);
  nand GNAME2418(G2418,G1646,G1566);
  nand GNAME2419(G2419,G2153,G12332);
  nand GNAME2420(G2420,G2152,G1585);
  nand GNAME2421(G2421,G2151,G11125);
  nand GNAME2422(G2422,G2420,G2421,G2419,G2417,G2418);
  nand GNAME2423(G2423,G3634,G36129);
  nand GNAME2424(G2424,G3637,G36097);
  nand GNAME2425(G2425,G3640,G36065);
  nand GNAME2426(G2426,G3631,G12130);
  nand GNAME2427(G2427,G1649,G1577);
  nand GNAME2428(G2428,G1647,G1566);
  nand GNAME2429(G2429,G2153,G12330);
  nand GNAME2430(G2430,G2152,G1586);
  nand GNAME2431(G2431,G2151,G11124);
  nand GNAME2432(G2432,G2430,G2431,G2429,G2427,G2428);
  nand GNAME2433(G2433,G3631,G12086);
  nand GNAME2434(G2434,G3634,G36130);
  nand GNAME2435(G2435,G3637,G36098);
  nand GNAME2436(G2436,G3640,G36066);
  nand GNAME2437(G2437,G1646,G1577);
  nand GNAME2438(G2438,G1641,G1566);
  nand GNAME2439(G2439,G2153,G12328);
  nand GNAME2440(G2440,G2152,G1587);
  nand GNAME2441(G2441,G2151,G11123);
  nand GNAME2442(G2442,G2440,G2441,G2439,G2437,G2438);
  nand GNAME2443(G2443,G3634,G36131);
  nand GNAME2444(G2444,G3637,G36099);
  nand GNAME2445(G2445,G3640,G36067);
  nand GNAME2446(G2446,G1558,G3643);
  nand GNAME2447(G2447,G2446,G2016);
  nand GNAME2448(G2448,G1244,G2447);
  nand GNAME2449(G2449,G1647,G1717);
  nand GNAME2450(G2450,G2448,G2449);
  nand GNAME2451(G2451,G2153,G12326);
  nand GNAME2452(G2452,G2152,G1588);
  nand GNAME2453(G2453,G2151,G11122);
  nand GNAME2454(G2454,G2450,G1565);
  nand GNAME2455(G2455,G2451,G2452,G2453,G2454);
  nand GNAME2456(G2456,G3634,G36132);
  nand GNAME2457(G2457,G3637,G36100);
  nand GNAME2458(G2458,G3640,G36068);
  nand GNAME2459(G2459,G1589,G12322);
  nand GNAME2460(G2460,G2152,G1590);
  nand GNAME2461(G2461,G2460,G2030,G2459);
  nand GNAME2462(G2462,G1589,G12211);
  nand GNAME2463(G2463,G2152,G1591);
  nand GNAME2464(G2464,G2463,G2030,G2462);
  nand GNAME2465(G2465,G3671,G1592);
  or GNAME2466(G2466,G1720,G1593);
  nand GNAME2467(G2467,G2466,G2018,G2465);
  nand GNAME2468(G2468,G3655,G3652);
  nand GNAME2469(G2469,G1594,G2014,G1564);
  nand GNAME2470(G2470,G2469,G1600);
  not GNAME2471(G2471,G1613);
  nand GNAME2472(G2472,G1718,G1721);
  nand GNAME2473(G2473,G2472,G1574);
  nand GNAME2474(G2474,G1631,G1597);
  nand GNAME2475(G2475,G12212,G1598);
  nand GNAME2476(G2476,G11117,G1599);
  nand GNAME2477(G2477,G36195,G1601);
  nand GNAME2478(G2478,G1724,G1603);
  nand GNAME2479(G2479,G1596,G36101);
  nand GNAME2480(G2480,G1572,G1605);
  nand GNAME2481(G2481,G2480,G11132);
  nand GNAME2482(G2482,G1612,G12275);
  nand GNAME2483(G2483,G1613,G1729);
  nand GNAME2484(G2484,G36205,G2011);
  nand GNAME2485(G2485,G2484,G1578,G2483,G2481,G2482);
  nand GNAME2486(G2486,G1631,G1607);
  nand GNAME2487(G2487,G1629,G1597);
  nand GNAME2488(G2488,G12324,G1598);
  nand GNAME2489(G2489,G11066,G1599);
  nand GNAME2490(G2490,G36190,G1601);
  nand GNAME2491(G2491,G1732,G1603);
  nand GNAME2492(G2492,G1596,G36103);
  nand GNAME2493(G2493,G1633,G1607);
  nand GNAME2494(G2494,G1632,G1597);
  nand GNAME2495(G2495,G12319,G1598);
  nand GNAME2496(G2496,G11069,G1599);
  nand GNAME2497(G2497,G12085,G1601);
  nand GNAME2498(G2498,G1735,G1603);
  nand GNAME2499(G2499,G1596,G36104);
  nand GNAME2500(G2500,G1629,G1607);
  nand GNAME2501(G2501,G1636,G1597);
  nand GNAME2502(G2502,G12317,G1598);
  nand GNAME2503(G2503,G11121,G1599);
  nand GNAME2504(G2504,G12129,G1601);
  nand GNAME2505(G2505,G1738,G1603);
  nand GNAME2506(G2506,G1596,G36105);
  nand GNAME2507(G2507,G1632,G1607);
  nand GNAME2508(G2508,G1634,G1597);
  nand GNAME2509(G2509,G12315,G1598);
  nand GNAME2510(G2510,G11120,G1599);
  nand GNAME2511(G2511,G12128,G1601);
  nand GNAME2512(G2512,G1741,G1603);
  nand GNAME2513(G2513,G1596,G36106);
  nand GNAME2514(G2514,G1636,G1607);
  nand GNAME2515(G2515,G1635,G1597);
  nand GNAME2516(G2516,G12313,G1598);
  nand GNAME2517(G2517,G11070,G1599);
  nand GNAME2518(G2518,G12127,G1601);
  nand GNAME2519(G2519,G1744,G1603);
  nand GNAME2520(G2520,G1596,G36107);
  nand GNAME2521(G2521,G1634,G1607);
  nand GNAME2522(G2522,G1630,G1597);
  nand GNAME2523(G2523,G12311,G1598);
  nand GNAME2524(G2524,G11071,G1599);
  nand GNAME2525(G2525,G12126,G1601);
  nand GNAME2526(G2526,G1747,G1603);
  nand GNAME2527(G2527,G1596,G36108);
  nand GNAME2528(G2528,G1635,G1607);
  nand GNAME2529(G2529,G1638,G1597);
  nand GNAME2530(G2530,G12309,G1598);
  nand GNAME2531(G2531,G11119,G1599);
  nand GNAME2532(G2532,G12125,G1601);
  nand GNAME2533(G2533,G1750,G1603);
  nand GNAME2534(G2534,G1596,G36109);
  nand GNAME2535(G2535,G1630,G1607);
  nand GNAME2536(G2536,G1637,G1597);
  nand GNAME2537(G2537,G12307,G1598);
  nand GNAME2538(G2538,G11118,G1599);
  nand GNAME2539(G2539,G12124,G1601);
  nand GNAME2540(G2540,G1753,G1603);
  nand GNAME2541(G2541,G1596,G36110);
  nand GNAME2542(G2542,G1638,G1607);
  nand GNAME2543(G2543,G1650,G1597);
  nand GNAME2544(G2544,G12365,G1598);
  nand GNAME2545(G2545,G11063,G1599);
  nand GNAME2546(G2546,G12148,G1601);
  nand GNAME2547(G2547,G1756,G1603);
  nand GNAME2548(G2548,G1596,G36111);
  nand GNAME2549(G2549,G1637,G1607);
  nand GNAME2550(G2550,G1654,G1597);
  nand GNAME2551(G2551,G12363,G1598);
  nand GNAME2552(G2552,G11064,G1599);
  nand GNAME2553(G2553,G12147,G1601);
  nand GNAME2554(G2554,G1759,G1603);
  nand GNAME2555(G2555,G1596,G36112);
  nand GNAME2556(G2556,G1650,G1607);
  nand GNAME2557(G2557,G1652,G1597);
  nand GNAME2558(G2558,G12361,G1598);
  nand GNAME2559(G2559,G11139,G1599);
  nand GNAME2560(G2560,G12146,G1601);
  nand GNAME2561(G2561,G1762,G1603);
  nand GNAME2562(G2562,G1596,G36113);
  nand GNAME2563(G2563,G1654,G1607);
  nand GNAME2564(G2564,G1651,G1597);
  nand GNAME2565(G2565,G12359,G1598);
  nand GNAME2566(G2566,G11138,G1599);
  nand GNAME2567(G2567,G12145,G1601);
  nand GNAME2568(G2568,G1765,G1603);
  nand GNAME2569(G2569,G1596,G36114);
  nand GNAME2570(G2570,G1652,G1607);
  nand GNAME2571(G2571,G1648,G1597);
  nand GNAME2572(G2572,G12357,G1598);
  nand GNAME2573(G2573,G11065,G1599);
  nand GNAME2574(G2574,G12144,G1601);
  nand GNAME2575(G2575,G1768,G1603);
  nand GNAME2576(G2576,G1596,G36115);
  nand GNAME2577(G2577,G1651,G1607);
  nand GNAME2578(G2578,G1653,G1597);
  nand GNAME2579(G2579,G12355,G1598);
  nand GNAME2580(G2580,G11137,G1599);
  nand GNAME2581(G2581,G12143,G1601);
  nand GNAME2582(G2582,G1771,G1603);
  nand GNAME2583(G2583,G1596,G36116);
  nand GNAME2584(G2584,G1648,G1607);
  nand GNAME2585(G2585,G1655,G1597);
  nand GNAME2586(G2586,G12353,G1598);
  nand GNAME2587(G2587,G11136,G1599);
  nand GNAME2588(G2588,G12142,G1601);
  nand GNAME2589(G2589,G1774,G1603);
  nand GNAME2590(G2590,G1596,G36117);
  nand GNAME2591(G2591,G1653,G1607);
  nand GNAME2592(G2592,G1657,G1597);
  nand GNAME2593(G2593,G12351,G1598);
  nand GNAME2594(G2594,G11135,G1599);
  nand GNAME2595(G2595,G12141,G1601);
  nand GNAME2596(G2596,G1777,G1603);
  nand GNAME2597(G2597,G1596,G36118);
  nand GNAME2598(G2598,G1655,G1607);
  nand GNAME2599(G2599,G1656,G1597);
  nand GNAME2600(G2600,G12349,G1598);
  nand GNAME2601(G2601,G11134,G1599);
  nand GNAME2602(G2602,G12140,G1601);
  nand GNAME2603(G2603,G1780,G1603);
  nand GNAME2604(G2604,G1596,G36119);
  nand GNAME2605(G2605,G1657,G1607);
  nand GNAME2606(G2606,G1644,G1597);
  nand GNAME2607(G2607,G12347,G1598);
  nand GNAME2608(G2608,G11133,G1599);
  nand GNAME2609(G2609,G12139,G1601);
  nand GNAME2610(G2610,G1782,G1603);
  nand GNAME2611(G2611,G1596,G36120);
  nand GNAME2612(G2612,G1656,G1607);
  nand GNAME2613(G2613,G1640,G1597);
  nand GNAME2614(G2614,G12344,G1598);
  nand GNAME2615(G2615,G11131,G1599);
  nand GNAME2616(G2616,G12138,G1601);
  nand GNAME2617(G2617,G1579,G1603);
  nand GNAME2618(G2618,G1596,G36121);
  nand GNAME2619(G2619,G1644,G1607);
  nand GNAME2620(G2620,G1645,G1597);
  nand GNAME2621(G2621,G12342,G1598);
  nand GNAME2622(G2622,G11130,G1599);
  nand GNAME2623(G2623,G12137,G1601);
  nand GNAME2624(G2624,G1580,G1603);
  nand GNAME2625(G2625,G1596,G36122);
  nand GNAME2626(G2626,G1640,G1607);
  nand GNAME2627(G2627,G1643,G1597);
  nand GNAME2628(G2628,G12340,G1598);
  nand GNAME2629(G2629,G11129,G1599);
  nand GNAME2630(G2630,G12136,G1601);
  nand GNAME2631(G2631,G1581,G1603);
  nand GNAME2632(G2632,G1596,G36123);
  nand GNAME2633(G2633,G1645,G1607);
  nand GNAME2634(G2634,G1639,G1597);
  nand GNAME2635(G2635,G12338,G1598);
  nand GNAME2636(G2636,G11128,G1599);
  nand GNAME2637(G2637,G12135,G1601);
  nand GNAME2638(G2638,G1582,G1603);
  nand GNAME2639(G2639,G1596,G36124);
  nand GNAME2640(G2640,G1643,G1607);
  nand GNAME2641(G2641,G1642,G1597);
  nand GNAME2642(G2642,G12336,G1598);
  nand GNAME2643(G2643,G11127,G1599);
  nand GNAME2644(G2644,G12134,G1601);
  nand GNAME2645(G2645,G1583,G1603);
  nand GNAME2646(G2646,G1596,G36125);
  nand GNAME2647(G2647,G1639,G1607);
  nand GNAME2648(G2648,G1649,G1597);
  nand GNAME2649(G2649,G12334,G1598);
  nand GNAME2650(G2650,G11126,G1599);
  nand GNAME2651(G2651,G12133,G1601);
  nand GNAME2652(G2652,G1584,G1603);
  nand GNAME2653(G2653,G1596,G36126);
  nand GNAME2654(G2654,G1642,G1607);
  nand GNAME2655(G2655,G1646,G1597);
  nand GNAME2656(G2656,G12332,G1598);
  nand GNAME2657(G2657,G11125,G1599);
  nand GNAME2658(G2658,G12132,G1601);
  nand GNAME2659(G2659,G1585,G1603);
  nand GNAME2660(G2660,G1596,G36127);
  nand GNAME2661(G2661,G1649,G1607);
  nand GNAME2662(G2662,G1647,G1597);
  nand GNAME2663(G2663,G12330,G1598);
  nand GNAME2664(G2664,G11124,G1599);
  nand GNAME2665(G2665,G12131,G1601);
  nand GNAME2666(G2666,G1586,G1603);
  nand GNAME2667(G2667,G1596,G36128);
  nand GNAME2668(G2668,G1646,G1607);
  nand GNAME2669(G2669,G1641,G1597);
  nand GNAME2670(G2670,G12328,G1598);
  nand GNAME2671(G2671,G11123,G1599);
  nand GNAME2672(G2672,G12130,G1601);
  nand GNAME2673(G2673,G1587,G1603);
  nand GNAME2674(G2674,G1596,G36129);
  nand GNAME2675(G2675,G12326,G1598);
  nand GNAME2676(G2676,G11122,G1599);
  nand GNAME2677(G2677,G12086,G1601);
  nand GNAME2678(G2678,G1588,G1603);
  nand GNAME2679(G2679,G12322,G2010);
  nand GNAME2680(G2680,G2679,G2030);
  nand GNAME2681(G2681,G1590,G1603);
  nand GNAME2682(G2682,G12211,G2010);
  nand GNAME2683(G2683,G2682,G2030);
  nand GNAME2684(G2684,G1591,G1603);
  or GNAME2685(G2685,G1616,G1617);
  or GNAME2686(G2686,G1620,G3660);
  nand GNAME2687(G2687,G11133,G1614);
  nand GNAME2688(G2688,G1615,G11517);
  nand GNAME2689(G2689,G1721,G1618);
  nand GNAME2690(G2690,G2689,G2687,G2688);
  or GNAME2691(G2691,G1565,G1556);
  nand GNAME2692(G2692,G2691,G3624);
  nand GNAME2693(G2693,G2016,G2692);
  not GNAME2694(G2694,G1622);
  nand GNAME2695(G2695,G1714,G1620);
  nand GNAME2696(G2696,G2695,G2005);
  nand GNAME2697(G2697,G1610,G1611);
  nand GNAME2698(G2698,G2690,G1619);
  nand GNAME2699(G2699,G11517,G1621);
  nand GNAME2700(G2700,G2694,G36133);
  nand GNAME2701(G2701,G11134,G1614);
  nand GNAME2702(G2702,G1615,G11560);
  nand GNAME2703(G2703,G1779,G1618);
  nand GNAME2704(G2704,G2703,G2701,G2702);
  nand GNAME2705(G2705,G2704,G1619);
  nand GNAME2706(G2706,G1621,G11560);
  nand GNAME2707(G2707,G1779,G1623);
  nand GNAME2708(G2708,G2694,G36134);
  nand GNAME2709(G2709,G11135,G1614);
  nand GNAME2710(G2710,G1615,G11561);
  nand GNAME2711(G2711,G1776,G1618);
  nand GNAME2712(G2712,G2711,G2709,G2710);
  nand GNAME2713(G2713,G2712,G1619);
  nand GNAME2714(G2714,G1621,G11561);
  nand GNAME2715(G2715,G1776,G1623);
  nand GNAME2716(G2716,G2694,G36135);
  nand GNAME2717(G2717,G11136,G1614);
  nand GNAME2718(G2718,G1615,G11562);
  nand GNAME2719(G2719,G1773,G1618);
  nand GNAME2720(G2720,G2719,G2717,G2718);
  nand GNAME2721(G2721,G2720,G1619);
  nand GNAME2722(G2722,G1621,G11562);
  nand GNAME2723(G2723,G1773,G1623);
  nand GNAME2724(G2724,G2694,G36136);
  nand GNAME2725(G2725,G11137,G1614);
  nand GNAME2726(G2726,G1615,G11516);
  nand GNAME2727(G2727,G1770,G1618);
  nand GNAME2728(G2728,G2727,G2725,G2726);
  nand GNAME2729(G2729,G2728,G1619);
  nand GNAME2730(G2730,G1621,G11516);
  nand GNAME2731(G2731,G1770,G1623);
  nand GNAME2732(G2732,G2694,G36137);
  nand GNAME2733(G2733,G11065,G1614);
  nand GNAME2734(G2734,G1615,G11515);
  nand GNAME2735(G2735,G1767,G1618);
  nand GNAME2736(G2736,G2735,G2733,G2734);
  nand GNAME2737(G2737,G2736,G1619);
  nand GNAME2738(G2738,G1621,G11515);
  nand GNAME2739(G2739,G1767,G1623);
  nand GNAME2740(G2740,G2694,G36138);
  nand GNAME2741(G2741,G11138,G1614);
  nand GNAME2742(G2742,G1615,G11563);
  nand GNAME2743(G2743,G1764,G1618);
  nand GNAME2744(G2744,G2743,G2741,G2742);
  nand GNAME2745(G2745,G2744,G1619);
  nand GNAME2746(G2746,G1621,G11563);
  nand GNAME2747(G2747,G1764,G1623);
  nand GNAME2748(G2748,G2694,G36139);
  nand GNAME2749(G2749,G11139,G1614);
  nand GNAME2750(G2750,G1615,G11564);
  nand GNAME2751(G2751,G1761,G1618);
  nand GNAME2752(G2752,G2751,G2749,G2750);
  nand GNAME2753(G2753,G2752,G1619);
  nand GNAME2754(G2754,G1621,G11564);
  nand GNAME2755(G2755,G1761,G1623);
  nand GNAME2756(G2756,G2694,G36140);
  nand GNAME2757(G2757,G11064,G1614);
  nand GNAME2758(G2758,G1615,G11514);
  nand GNAME2759(G2759,G1758,G1618);
  nand GNAME2760(G2760,G2759,G2757,G2758);
  nand GNAME2761(G2761,G2760,G1619);
  nand GNAME2762(G2762,G1621,G11514);
  nand GNAME2763(G2763,G1758,G1623);
  nand GNAME2764(G2764,G2694,G36141);
  nand GNAME2765(G2765,G11063,G1614);
  nand GNAME2766(G2766,G1615,G11513);
  nand GNAME2767(G2767,G1755,G1618);
  nand GNAME2768(G2768,G2767,G2765,G2766);
  nand GNAME2769(G2769,G2768,G1619);
  nand GNAME2770(G2770,G1621,G11513);
  nand GNAME2771(G2771,G1755,G1623);
  nand GNAME2772(G2772,G2694,G36142);
  nand GNAME2773(G2773,G11118,G1614);
  nand GNAME2774(G2774,G1615,G11552);
  nand GNAME2775(G2775,G1752,G1618);
  nand GNAME2776(G2776,G2775,G2773,G2774);
  nand GNAME2777(G2777,G2776,G1619);
  nand GNAME2778(G2778,G1621,G11552);
  nand GNAME2779(G2779,G1752,G1623);
  nand GNAME2780(G2780,G2694,G36143);
  nand GNAME2781(G2781,G11119,G1614);
  nand GNAME2782(G2782,G1615,G11553);
  nand GNAME2783(G2783,G1749,G1618);
  nand GNAME2784(G2784,G2783,G2781,G2782);
  nand GNAME2785(G2785,G2784,G1619);
  nand GNAME2786(G2786,G1621,G11553);
  nand GNAME2787(G2787,G1749,G1623);
  nand GNAME2788(G2788,G2694,G36144);
  nand GNAME2789(G2789,G11071,G1614);
  nand GNAME2790(G2790,G1615,G11554);
  nand GNAME2791(G2791,G1746,G1618);
  nand GNAME2792(G2792,G2791,G2789,G2790);
  nand GNAME2793(G2793,G2792,G1619);
  nand GNAME2794(G2794,G1621,G11554);
  nand GNAME2795(G2795,G1746,G1623);
  nand GNAME2796(G2796,G2694,G36145);
  nand GNAME2797(G2797,G11070,G1614);
  nand GNAME2798(G2798,G1615,G11555);
  nand GNAME2799(G2799,G1743,G1618);
  nand GNAME2800(G2800,G2799,G2797,G2798);
  nand GNAME2801(G2801,G2800,G1619);
  nand GNAME2802(G2802,G1621,G11555);
  nand GNAME2803(G2803,G1743,G1623);
  nand GNAME2804(G2804,G2694,G36146);
  nand GNAME2805(G2805,G11120,G1614);
  nand GNAME2806(G2806,G1615,G11556);
  nand GNAME2807(G2807,G1740,G1618);
  nand GNAME2808(G2808,G2807,G2805,G2806);
  nand GNAME2809(G2809,G2808,G1619);
  nand GNAME2810(G2810,G1621,G11556);
  nand GNAME2811(G2811,G1740,G1623);
  nand GNAME2812(G2812,G2694,G36147);
  nand GNAME2813(G2813,G11121,G1614);
  nand GNAME2814(G2814,G1615,G11557);
  nand GNAME2815(G2815,G1737,G1618);
  nand GNAME2816(G2816,G2815,G2813,G2814);
  nand GNAME2817(G2817,G2816,G1619);
  nand GNAME2818(G2818,G1621,G11557);
  nand GNAME2819(G2819,G1737,G1623);
  nand GNAME2820(G2820,G2694,G36148);
  nand GNAME2821(G2821,G11069,G1614);
  nand GNAME2822(G2822,G1615,G11558);
  nand GNAME2823(G2823,G1734,G1618);
  nand GNAME2824(G2824,G2823,G2821,G2822);
  nand GNAME2825(G2825,G2824,G1619);
  nand GNAME2826(G2826,G1621,G11558);
  nand GNAME2827(G2827,G1734,G1623);
  nand GNAME2828(G2828,G2694,G36149);
  nand GNAME2829(G2829,G11066,G1614);
  nand GNAME2830(G2830,G1615,G11559);
  nand GNAME2831(G2831,G1731,G1618);
  nand GNAME2832(G2832,G2831,G2829,G2830);
  nand GNAME2833(G2833,G2832,G1619);
  nand GNAME2834(G2834,G1621,G11559);
  nand GNAME2835(G2835,G1731,G1623);
  nand GNAME2836(G2836,G2694,G36150);
  nand GNAME2837(G2837,G11132,G1614);
  nand GNAME2838(G2838,G1615,G11518);
  nand GNAME2839(G2839,G1728,G1618);
  nand GNAME2840(G2840,G2839,G2837,G2838);
  nand GNAME2841(G2841,G2840,G1619);
  nand GNAME2842(G2842,G1621,G11518);
  nand GNAME2843(G2843,G1728,G1623);
  nand GNAME2844(G2844,G2694,G36151);
  nand GNAME2845(G2845,G11117,G1614);
  nand GNAME2846(G2846,G1615,G11551);
  nand GNAME2847(G2847,G1722,G1618);
  nand GNAME2848(G2848,G2847,G2845,G2846);
  nand GNAME2849(G2849,G2848,G1619);
  nand GNAME2850(G2850,G1621,G11551);
  nand GNAME2851(G2851,G1722,G1623);
  nand GNAME2852(G2852,G2694,G36152);
  nand GNAME2853(G2853,G1661,G1659,G1660);
  nand GNAME2854(G2854,G1662,G1659,G1660);
  nand GNAME2855(G2855,G2853,G2854);
  nand GNAME2856(G2856,G2015,G1611);
  nand GNAME2857(G2857,G2855,G4041);
  nand GNAME2858(G2858,G2856,G2857);
  nand GNAME2859(G2859,G3612,G4045,G4046);
  or GNAME2860(G2860,G3655,G11727,G1998,G1604);
  nand GNAME2861(G2861,G2858,G1561);
  nand GNAME2862(G2862,G2859,G3652);
  nand GNAME2863(G2863,G2860,G2861,G2862,G4047,G4048);
  nor GNAME2864(G2864,G1627,G1714);
  or GNAME2865(G2865,G1406,G1624,G1628,G2864);
  nand GNAME2866(G2866,G1627,G1663,G1559);
  nand GNAME2867(G2867,G2865,G36185);
  nand GNAME2868(G2868,G36215,G2863);
  nand GNAME2869(G2869,G1651,G1675);
  nand GNAME2870(G2870,G1653,G1676);
  nand GNAME2871(G2871,G1666,G12143);
  nand GNAME2872(G2872,G2871,G2869,G2870);
  or GNAME2873(G2873,G1604,G1719);
  nand GNAME2874(G2874,G1606,G3646);
  or GNAME2875(G2875,G1669,G1670);
  nand GNAME2876(G2876,G1666,G2875);
  nand GNAME2877(G2877,G2876,G2014);
  nand GNAME2878(G2878,G2877,G1559);
  nand GNAME2879(G2879,G36215,G1714);
  nand GNAME2880(G2880,G3611,G1771);
  nand GNAME2881(G2881,G3610,G12143);
  nand GNAME2882(G2882,G12355,G1673);
  nand GNAME2883(G2883,G11137,G1674);
  nand GNAME2884(G2884,G2872,G1677);
  nand GNAME2885(G2885,G1406,G36186);
  nand GNAME2886(G2886,G1642,G1675);
  nand GNAME2887(G2887,G1646,G1676);
  nand GNAME2888(G2888,G1666,G12132);
  nand GNAME2889(G2889,G2888,G2886,G2887);
  nand GNAME2890(G2890,G1613,G2017);
  nand GNAME2891(G2891,G2890,G1600);
  nand GNAME2892(G2892,G1585,G1678);
  nand GNAME2893(G2893,G12332,G1673);
  nand GNAME2894(G2894,G11125,G1674);
  nand GNAME2895(G2895,G2889,G1677);
  nand GNAME2896(G2896,G3610,G12132);
  nand GNAME2897(G2897,G1406,G36187);
  nand GNAME2898(G2898,G1636,G1675);
  nand GNAME2899(G2899,G1635,G1676);
  nand GNAME2900(G2900,G1666,G12127);
  nand GNAME2901(G2901,G2900,G2898,G2899);
  nand GNAME2902(G2902,G3611,G1744);
  nand GNAME2903(G2903,G3610,G12127);
  nand GNAME2904(G2904,G12313,G1673);
  nand GNAME2905(G2905,G11070,G1674);
  nand GNAME2906(G2906,G2901,G1677);
  nand GNAME2907(G2907,G1406,G36188);
  nand GNAME2908(G2908,G1655,G1675);
  nand GNAME2909(G2909,G1656,G1676);
  nand GNAME2910(G2910,G1666,G12140);
  nand GNAME2911(G2911,G2910,G2908,G2909);
  nand GNAME2912(G2912,G3611,G1780);
  nand GNAME2913(G2913,G3610,G12140);
  nand GNAME2914(G2914,G12349,G1673);
  nand GNAME2915(G2915,G11134,G1674);
  nand GNAME2916(G2916,G2911,G1677);
  nand GNAME2917(G2917,G1406,G36189);
  nand GNAME2918(G2918,G1631,G1675);
  nand GNAME2919(G2919,G1629,G1676);
  nand GNAME2920(G2920,G1666,G36190);
  nand GNAME2921(G2921,G2920,G2918,G2919);
  nand GNAME2922(G2922,G3611,G1732);
  nand GNAME2923(G2923,G3610,G36190);
  nand GNAME2924(G2924,G12324,G1673);
  nand GNAME2925(G2925,G11066,G1674);
  nand GNAME2926(G2926,G2921,G1677);
  nand GNAME2927(G2927,G1406,G36190);
  nand GNAME2928(G2928,G1637,G1675);
  nand GNAME2929(G2929,G1654,G1676);
  nand GNAME2930(G2930,G1666,G12147);
  nand GNAME2931(G2931,G2930,G2928,G2929);
  nand GNAME2932(G2932,G3611,G1759);
  nand GNAME2933(G2933,G3610,G12147);
  nand GNAME2934(G2934,G12363,G1673);
  nand GNAME2935(G2935,G11064,G1674);
  nand GNAME2936(G2936,G2931,G1677);
  nand GNAME2937(G2937,G1406,G36191);
  nand GNAME2938(G2938,G1640,G1675);
  nand GNAME2939(G2939,G1643,G1676);
  nand GNAME2940(G2940,G1666,G12136);
  nand GNAME2941(G2941,G2940,G2938,G2939);
  nand GNAME2942(G2942,G1581,G1678);
  nand GNAME2943(G2943,G12340,G1673);
  nand GNAME2944(G2944,G11129,G1674);
  nand GNAME2945(G2945,G2941,G1677);
  nand GNAME2946(G2946,G3610,G12136);
  nand GNAME2947(G2947,G1406,G36192);
  nand GNAME2948(G2948,G1654,G1675);
  nand GNAME2949(G2949,G1651,G1676);
  nand GNAME2950(G2950,G1666,G12145);
  nand GNAME2951(G2951,G2950,G2948,G2949);
  nand GNAME2952(G2952,G3611,G1765);
  nand GNAME2953(G2953,G3610,G12145);
  nand GNAME2954(G2954,G12359,G1673);
  nand GNAME2955(G2955,G11138,G1674);
  nand GNAME2956(G2956,G2951,G1677);
  nand GNAME2957(G2957,G1406,G36193);
  nand GNAME2958(G2958,G1656,G1675);
  nand GNAME2959(G2959,G1640,G1676);
  nand GNAME2960(G2960,G1666,G12138);
  nand GNAME2961(G2961,G2960,G2958,G2959);
  nand GNAME2962(G2962,G1579,G1678);
  nand GNAME2963(G2963,G12344,G1673);
  nand GNAME2964(G2964,G11131,G1674);
  nand GNAME2965(G2965,G2961,G1677);
  nand GNAME2966(G2966,G3610,G12138);
  nand GNAME2967(G2967,G1406,G36194);
  or GNAME2968(G2968,G1665,G1677);
  nand GNAME2969(G2969,G1666,G2968);
  nand GNAME2970(G2970,G2969,G1671);
  nand GNAME2971(G2971,G1677,G1631,G1676);
  nand GNAME2972(G2972,G3611,G1724);
  nand GNAME2973(G2973,G2970,G36195);
  nand GNAME2974(G2974,G12212,G1673);
  nand GNAME2975(G2975,G11117,G1674);
  nand GNAME2976(G2976,G1406,G36195);
  nand GNAME2977(G2977,G1630,G1675);
  nand GNAME2978(G2978,G1637,G1676);
  nand GNAME2979(G2979,G1666,G12124);
  nand GNAME2980(G2980,G2979,G2977,G2978);
  nand GNAME2981(G2981,G3611,G1753);
  nand GNAME2982(G2982,G3610,G12124);
  nand GNAME2983(G2983,G12307,G1673);
  nand GNAME2984(G2984,G11118,G1674);
  nand GNAME2985(G2985,G2980,G1677);
  nand GNAME2986(G2986,G1406,G36196);
  nand GNAME2987(G2987,G1629,G1675);
  nand GNAME2988(G2988,G1636,G1676);
  nand GNAME2989(G2989,G1666,G12129);
  nand GNAME2990(G2990,G2989,G2987,G2988);
  nand GNAME2991(G2991,G3611,G1738);
  nand GNAME2992(G2992,G3610,G12129);
  nand GNAME2993(G2993,G12317,G1673);
  nand GNAME2994(G2994,G11121,G1674);
  nand GNAME2995(G2995,G2990,G1677);
  nand GNAME2996(G2996,G1406,G36197);
  nand GNAME2997(G2997,G1643,G1675);
  nand GNAME2998(G2998,G1642,G1676);
  nand GNAME2999(G2999,G1666,G12134);
  nand GNAME3000(G3000,G2999,G2997,G2998);
  nand GNAME3001(G3001,G1583,G1678);
  nand GNAME3002(G3002,G12336,G1673);
  nand GNAME3003(G3003,G11127,G1674);
  nand GNAME3004(G3004,G3000,G1677);
  nand GNAME3005(G3005,G3610,G12134);
  nand GNAME3006(G3006,G1406,G36198);
  nand GNAME3007(G3007,G1653,G1675);
  nand GNAME3008(G3008,G1657,G1676);
  nand GNAME3009(G3009,G1666,G12141);
  nand GNAME3010(G3010,G3009,G3007,G3008);
  nand GNAME3011(G3011,G3611,G1777);
  nand GNAME3012(G3012,G3610,G12141);
  nand GNAME3013(G3013,G12351,G1673);
  nand GNAME3014(G3014,G11135,G1674);
  nand GNAME3015(G3015,G3010,G1677);
  nand GNAME3016(G3016,G1406,G36199);
  nand GNAME3017(G3017,G1632,G1675);
  nand GNAME3018(G3018,G1634,G1676);
  nand GNAME3019(G3019,G1666,G12128);
  nand GNAME3020(G3020,G3019,G3017,G3018);
  nand GNAME3021(G3021,G3611,G1741);
  nand GNAME3022(G3022,G3610,G12128);
  nand GNAME3023(G3023,G12315,G1673);
  nand GNAME3024(G3024,G11120,G1674);
  nand GNAME3025(G3025,G3020,G1677);
  nand GNAME3026(G3026,G1406,G36200);
  nand GNAME3027(G3027,G1648,G1675);
  nand GNAME3028(G3028,G1655,G1676);
  nand GNAME3029(G3029,G1666,G12142);
  nand GNAME3030(G3030,G3029,G3027,G3028);
  nand GNAME3031(G3031,G3611,G1774);
  nand GNAME3032(G3032,G3610,G12142);
  nand GNAME3033(G3033,G12353,G1673);
  nand GNAME3034(G3034,G11136,G1674);
  nand GNAME3035(G3035,G3030,G1677);
  nand GNAME3036(G3036,G1406,G36201);
  nand GNAME3037(G3037,G1639,G1675);
  nand GNAME3038(G3038,G1649,G1676);
  nand GNAME3039(G3039,G1666,G12133);
  nand GNAME3040(G3040,G3039,G3037,G3038);
  nand GNAME3041(G3041,G1584,G1678);
  nand GNAME3042(G3042,G12334,G1673);
  nand GNAME3043(G3043,G11126,G1674);
  nand GNAME3044(G3044,G3040,G1677);
  nand GNAME3045(G3045,G3610,G12133);
  nand GNAME3046(G3046,G1406,G36202);
  nand GNAME3047(G3047,G1650,G1675);
  nand GNAME3048(G3048,G1652,G1676);
  nand GNAME3049(G3049,G1666,G12146);
  nand GNAME3050(G3050,G3049,G3047,G3048);
  nand GNAME3051(G3051,G3611,G1762);
  nand GNAME3052(G3052,G3610,G12146);
  nand GNAME3053(G3053,G12361,G1673);
  nand GNAME3054(G3054,G11139,G1674);
  nand GNAME3055(G3055,G3050,G1677);
  nand GNAME3056(G3056,G1406,G36203);
  nand GNAME3057(G3057,G1644,G1675);
  nand GNAME3058(G3058,G1645,G1676);
  nand GNAME3059(G3059,G1666,G12137);
  nand GNAME3060(G3060,G3059,G3057,G3058);
  nand GNAME3061(G3061,G1580,G1678);
  nand GNAME3062(G3062,G12342,G1673);
  nand GNAME3063(G3063,G11130,G1674);
  nand GNAME3064(G3064,G3060,G1677);
  nand GNAME3065(G3065,G3610,G12137);
  nand GNAME3066(G3066,G1406,G36204);
  nand GNAME3067(G3067,G1658,G1675);
  nand GNAME3068(G3068,G1633,G1676);
  nand GNAME3069(G3069,G1666,G36205);
  nand GNAME3070(G3070,G3069,G3067,G3068);
  nand GNAME3071(G3071,G3611,G1729);
  nand GNAME3072(G3072,G3610,G36205);
  nand GNAME3073(G3073,G12275,G1673);
  nand GNAME3074(G3074,G11132,G1674);
  nand GNAME3075(G3075,G3070,G1677);
  nand GNAME3076(G3076,G1406,G36205);
  nand GNAME3077(G3077,G1635,G1675);
  nand GNAME3078(G3078,G1638,G1676);
  nand GNAME3079(G3079,G1666,G12125);
  nand GNAME3080(G3080,G3079,G3077,G3078);
  nand GNAME3081(G3081,G3611,G1750);
  nand GNAME3082(G3082,G3610,G12125);
  nand GNAME3083(G3083,G12309,G1673);
  nand GNAME3084(G3084,G11119,G1674);
  nand GNAME3085(G3085,G3080,G1677);
  nand GNAME3086(G3086,G1406,G36206);
  nand GNAME3087(G3087,G1646,G1675);
  nand GNAME3088(G3088,G1641,G1676);
  nand GNAME3089(G3089,G1666,G12130);
  nand GNAME3090(G3090,G3089,G3087,G3088);
  nand GNAME3091(G3091,G1587,G1678);
  nand GNAME3092(G3092,G12328,G1673);
  nand GNAME3093(G3093,G11123,G1674);
  nand GNAME3094(G3094,G3090,G1677);
  nand GNAME3095(G3095,G3610,G12130);
  nand GNAME3096(G3096,G1406,G36207);
  nand GNAME3097(G3097,G1657,G1675);
  nand GNAME3098(G3098,G1644,G1676);
  nand GNAME3099(G3099,G1666,G12139);
  nand GNAME3100(G3100,G3099,G3097,G3098);
  nand GNAME3101(G3101,G3611,G1782);
  nand GNAME3102(G3102,G3610,G12139);
  nand GNAME3103(G3103,G12347,G1673);
  nand GNAME3104(G3104,G11133,G1674);
  nand GNAME3105(G3105,G3100,G1677);
  nand GNAME3106(G3106,G1406,G36208);
  nand GNAME3107(G3107,G1633,G1675);
  nand GNAME3108(G3108,G1632,G1676);
  nand GNAME3109(G3109,G1666,G12085);
  nand GNAME3110(G3110,G3109,G3107,G3108);
  nand GNAME3111(G3111,G3611,G1735);
  nand GNAME3112(G3112,G3610,G12085);
  nand GNAME3113(G3113,G12319,G1673);
  nand GNAME3114(G3114,G11069,G1674);
  nand GNAME3115(G3115,G3110,G1677);
  nand GNAME3116(G3116,G1406,G36209);
  nand GNAME3117(G3117,G1638,G1675);
  nand GNAME3118(G3118,G1650,G1676);
  nand GNAME3119(G3119,G1666,G12148);
  nand GNAME3120(G3120,G3119,G3117,G3118);
  nand GNAME3121(G3121,G3611,G1756);
  nand GNAME3122(G3122,G3610,G12148);
  nand GNAME3123(G3123,G12365,G1673);
  nand GNAME3124(G3124,G11063,G1674);
  nand GNAME3125(G3125,G3120,G1677);
  nand GNAME3126(G3126,G1406,G36210);
  nand GNAME3127(G3127,G1645,G1675);
  nand GNAME3128(G3128,G1639,G1676);
  nand GNAME3129(G3129,G1666,G12135);
  nand GNAME3130(G3130,G3129,G3127,G3128);
  nand GNAME3131(G3131,G1582,G1678);
  nand GNAME3132(G3132,G12338,G1673);
  nand GNAME3133(G3133,G11128,G1674);
  nand GNAME3134(G3134,G3130,G1677);
  nand GNAME3135(G3135,G3610,G12135);
  nand GNAME3136(G3136,G1406,G36211);
  nand GNAME3137(G3137,G1652,G1675);
  nand GNAME3138(G3138,G1648,G1676);
  nand GNAME3139(G3139,G1666,G12144);
  nand GNAME3140(G3140,G3139,G3137,G3138);
  nand GNAME3141(G3141,G3611,G1768);
  nand GNAME3142(G3142,G3610,G12144);
  nand GNAME3143(G3143,G12357,G1673);
  nand GNAME3144(G3144,G11065,G1674);
  nand GNAME3145(G3145,G3140,G1677);
  nand GNAME3146(G3146,G1406,G36212);
  nand GNAME3147(G3147,G1649,G1675);
  nand GNAME3148(G3148,G1647,G1676);
  nand GNAME3149(G3149,G1666,G12131);
  nand GNAME3150(G3150,G3149,G3147,G3148);
  nand GNAME3151(G3151,G1586,G1678);
  nand GNAME3152(G3152,G12330,G1673);
  nand GNAME3153(G3153,G11124,G1674);
  nand GNAME3154(G3154,G3150,G1677);
  nand GNAME3155(G3155,G3610,G12131);
  nand GNAME3156(G3156,G1406,G36213);
  nand GNAME3157(G3157,G1634,G1675);
  nand GNAME3158(G3158,G1630,G1676);
  nand GNAME3159(G3159,G1666,G12126);
  nand GNAME3160(G3160,G3159,G3157,G3158);
  nand GNAME3161(G3161,G3611,G1747);
  nand GNAME3162(G3162,G3610,G12126);
  nand GNAME3163(G3163,G12311,G1673);
  nand GNAME3164(G3164,G11071,G1674);
  nand GNAME3165(G3165,G3160,G1677);
  nand GNAME3166(G3166,G1406,G36214);
  nand GNAME3167(G3167,G2024,G2019,G2020);
  or GNAME3168(G3168,G1706,G1707);
  nand GNAME3169(G3169,G1709,G1753);
  nand GNAME3170(G3170,G3168,G1752);
  nand GNAME3171(G3171,G1638,G3499);
  nand GNAME3172(G3172,G1709,G1750);
  nand GNAME3173(G3173,G3168,G1749);
  nand GNAME3174(G3174,G1630,G3499);
  nand GNAME3175(G3175,G1709,G1747);
  nand GNAME3176(G3176,G3168,G1746);
  nand GNAME3177(G3177,G1635,G3499);
  nand GNAME3178(G3178,G1709,G1744);
  nand GNAME3179(G3179,G3168,G1743);
  nand GNAME3180(G3180,G1634,G3499);
  nand GNAME3181(G3181,G1709,G1741);
  nand GNAME3182(G3182,G3168,G1740);
  nand GNAME3183(G3183,G1636,G3499);
  nand GNAME3184(G3184,G1709,G1738);
  nand GNAME3185(G3185,G3168,G1737);
  nand GNAME3186(G3186,G1632,G3499);
  nand GNAME3187(G3187,G2036,G1995,G2035);
  nand GNAME3188(G3188,G2002,G1999);
  nand GNAME3189(G3189,G3188,G1587);
  nand GNAME3190(G3190,G1647,G1688);
  nand GNAME3191(G3191,G3187,G1588);
  nand GNAME3192(G3192,G1641,G1689);
  nand GNAME3193(G3193,G1709,G1735);
  nand GNAME3194(G3194,G3168,G1734);
  nand GNAME3195(G3195,G1629,G3499);
  nand GNAME3196(G3196,G1709,G1587);
  nand GNAME3197(G3197,G1647,G3499);
  nand GNAME3198(G3198,G1709,G1586);
  nand GNAME3199(G3199,G1646,G3499);
  nand GNAME3200(G3200,G1709,G1585);
  nand GNAME3201(G3201,G1649,G3499);
  nand GNAME3202(G3202,G1709,G1584);
  nand GNAME3203(G3203,G1642,G3499);
  nand GNAME3204(G3204,G1709,G1583);
  nand GNAME3205(G3205,G1639,G3499);
  nand GNAME3206(G3206,G1709,G1582);
  nand GNAME3207(G3207,G1643,G3499);
  nand GNAME3208(G3208,G1709,G1581);
  nand GNAME3209(G3209,G1645,G3499);
  nand GNAME3210(G3210,G1709,G1580);
  nand GNAME3211(G3211,G1640,G3499);
  nand GNAME3212(G3212,G1709,G1579);
  nand GNAME3213(G3213,G1644,G3499);
  nand GNAME3214(G3214,G1709,G1732);
  nand GNAME3215(G3215,G3168,G1731);
  nand GNAME3216(G3216,G1633,G3499);
  nand GNAME3217(G3217,G1709,G1782);
  nand GNAME3218(G3218,G1656,G3499);
  nand GNAME3219(G3219,G1709,G1780);
  nand GNAME3220(G3220,G3168,G1779);
  nand GNAME3221(G3221,G1657,G3499);
  nand GNAME3222(G3222,G1709,G1777);
  nand GNAME3223(G3223,G3168,G1776);
  nand GNAME3224(G3224,G1655,G3499);
  nand GNAME3225(G3225,G1709,G1774);
  nand GNAME3226(G3226,G3168,G1773);
  nand GNAME3227(G3227,G1653,G3499);
  nand GNAME3228(G3228,G1709,G1771);
  nand GNAME3229(G3229,G3168,G1770);
  nand GNAME3230(G3230,G1648,G3499);
  nand GNAME3231(G3231,G1709,G1768);
  nand GNAME3232(G3232,G3168,G1767);
  nand GNAME3233(G3233,G1651,G3499);
  nand GNAME3234(G3234,G1709,G1765);
  nand GNAME3235(G3235,G3168,G1764);
  nand GNAME3236(G3236,G1652,G3499);
  nand GNAME3237(G3237,G1709,G1762);
  nand GNAME3238(G3238,G3168,G1761);
  nand GNAME3239(G3239,G1654,G3499);
  nand GNAME3240(G3240,G1709,G1759);
  nand GNAME3241(G3241,G3168,G1758);
  nand GNAME3242(G3242,G1650,G3499);
  nand GNAME3243(G3243,G1709,G1756);
  nand GNAME3244(G3244,G3168,G1755);
  nand GNAME3245(G3245,G1637,G3499);
  nand GNAME3246(G3246,G1709,G1729);
  nand GNAME3247(G3247,G3168,G1728);
  nand GNAME3248(G3248,G1631,G3499);
  nand GNAME3249(G3249,G1624,G4115,G4116);
  nand GNAME3250(G3250,G1709,G1724);
  nand GNAME3251(G3251,G3168,G1722);
  nand GNAME3252(G3252,G1658,G3499);
  nand GNAME3253(G3253,G1714,G1626);
  or GNAME3254(G3254,G12083,G1695);
  nand GNAME3255(G3255,G1692,G2009,G3254);
  or GNAME3256(G3256,G1569,G1606);
  nand GNAME3257(G3257,G3256,G3646);
  nand GNAME3258(G3258,G1693,G1691);
  nand GNAME3259(G3259,G11118,G1690);
  nand GNAME3260(G3260,G3258,G1753);
  nand GNAME3261(G3261,G1638,G3255);
  nand GNAME3262(G3262,G1630,G3624);
  nand GNAME3263(G3263,G11119,G1690);
  nand GNAME3264(G3264,G3258,G1750);
  nand GNAME3265(G3265,G1630,G3255);
  nand GNAME3266(G3266,G1635,G3624);
  nand GNAME3267(G3267,G11071,G1690);
  nand GNAME3268(G3268,G3258,G1747);
  nand GNAME3269(G3269,G1635,G3255);
  nand GNAME3270(G3270,G1634,G3624);
  nand GNAME3271(G3271,G11070,G1690);
  nand GNAME3272(G3272,G3258,G1744);
  nand GNAME3273(G3273,G1634,G3255);
  nand GNAME3274(G3274,G1636,G3624);
  nand GNAME3275(G3275,G11120,G1690);
  nand GNAME3276(G3276,G3258,G1741);
  nand GNAME3277(G3277,G1636,G3255);
  nand GNAME3278(G3278,G1632,G3624);
  nand GNAME3279(G3279,G11121,G1690);
  nand GNAME3280(G3280,G3258,G1738);
  nand GNAME3281(G3281,G1632,G3255);
  nand GNAME3282(G3282,G1629,G3624);
  nand GNAME3283(G3283,G1690,G11068);
  nand GNAME3284(G3284,G3258,G1591);
  nand GNAME3285(G3285,G1242,G3255);
  nand GNAME3286(G3286,G1690,G11067);
  nand GNAME3287(G3287,G3258,G1590);
  nand GNAME3288(G3288,G1244,G3255);
  nand GNAME3289(G3289,G11069,G1690);
  nand GNAME3290(G3290,G3258,G1735);
  nand GNAME3291(G3291,G1629,G3255);
  nand GNAME3292(G3292,G1633,G3624);
  nand GNAME3293(G3293,G11122,G1690);
  nand GNAME3294(G3294,G3258,G1588);
  nand GNAME3295(G3295,G1641,G3255);
  nand GNAME3296(G3296,G1647,G3624);
  nand GNAME3297(G3297,G11123,G1690);
  nand GNAME3298(G3298,G3258,G1587);
  nand GNAME3299(G3299,G1647,G3255);
  nand GNAME3300(G3300,G1646,G3624);
  nand GNAME3301(G3301,G11124,G1690);
  nand GNAME3302(G3302,G3258,G1586);
  nand GNAME3303(G3303,G1646,G3255);
  nand GNAME3304(G3304,G1649,G3624);
  nand GNAME3305(G3305,G11125,G1690);
  nand GNAME3306(G3306,G3258,G1585);
  nand GNAME3307(G3307,G1649,G3255);
  nand GNAME3308(G3308,G1642,G3624);
  nand GNAME3309(G3309,G11126,G1690);
  nand GNAME3310(G3310,G3258,G1584);
  nand GNAME3311(G3311,G1642,G3255);
  nand GNAME3312(G3312,G1639,G3624);
  nand GNAME3313(G3313,G11127,G1690);
  nand GNAME3314(G3314,G3258,G1583);
  nand GNAME3315(G3315,G1639,G3255);
  nand GNAME3316(G3316,G1643,G3624);
  nand GNAME3317(G3317,G11128,G1690);
  nand GNAME3318(G3318,G3258,G1582);
  nand GNAME3319(G3319,G1643,G3255);
  nand GNAME3320(G3320,G1645,G3624);
  nand GNAME3321(G3321,G11129,G1690);
  nand GNAME3322(G3322,G3258,G1581);
  nand GNAME3323(G3323,G1645,G3255);
  nand GNAME3324(G3324,G1640,G3624);
  nand GNAME3325(G3325,G11130,G1690);
  nand GNAME3326(G3326,G3258,G1580);
  nand GNAME3327(G3327,G1640,G3255);
  nand GNAME3328(G3328,G1644,G3624);
  nand GNAME3329(G3329,G11131,G1690);
  nand GNAME3330(G3330,G3258,G1579);
  nand GNAME3331(G3331,G1644,G3255);
  nand GNAME3332(G3332,G1656,G3624);
  nand GNAME3333(G3333,G11066,G1690);
  nand GNAME3334(G3334,G3258,G1732);
  nand GNAME3335(G3335,G1633,G3255);
  nand GNAME3336(G3336,G1631,G3624);
  nand GNAME3337(G3337,G11133,G1690);
  nand GNAME3338(G3338,G3258,G1782);
  nand GNAME3339(G3339,G1656,G3255);
  nand GNAME3340(G3340,G1657,G3624);
  nand GNAME3341(G3341,G11134,G1690);
  nand GNAME3342(G3342,G3258,G1780);
  nand GNAME3343(G3343,G1657,G3255);
  nand GNAME3344(G3344,G1655,G3624);
  nand GNAME3345(G3345,G11135,G1690);
  nand GNAME3346(G3346,G3258,G1777);
  nand GNAME3347(G3347,G1655,G3255);
  nand GNAME3348(G3348,G1653,G3624);
  nand GNAME3349(G3349,G11136,G1690);
  nand GNAME3350(G3350,G3258,G1774);
  nand GNAME3351(G3351,G1653,G3255);
  nand GNAME3352(G3352,G1648,G3624);
  nand GNAME3353(G3353,G11137,G1690);
  nand GNAME3354(G3354,G3258,G1771);
  nand GNAME3355(G3355,G1648,G3255);
  nand GNAME3356(G3356,G1651,G3624);
  nand GNAME3357(G3357,G11065,G1690);
  nand GNAME3358(G3358,G3258,G1768);
  nand GNAME3359(G3359,G1651,G3255);
  nand GNAME3360(G3360,G1652,G3624);
  nand GNAME3361(G3361,G11138,G1690);
  nand GNAME3362(G3362,G3258,G1765);
  nand GNAME3363(G3363,G1652,G3255);
  nand GNAME3364(G3364,G1654,G3624);
  nand GNAME3365(G3365,G11139,G1690);
  nand GNAME3366(G3366,G3258,G1762);
  nand GNAME3367(G3367,G1654,G3255);
  nand GNAME3368(G3368,G1650,G3624);
  nand GNAME3369(G3369,G11064,G1690);
  nand GNAME3370(G3370,G3258,G1759);
  nand GNAME3371(G3371,G1650,G3255);
  nand GNAME3372(G3372,G1637,G3624);
  nand GNAME3373(G3373,G11063,G1690);
  nand GNAME3374(G3374,G3258,G1756);
  nand GNAME3375(G3375,G1637,G3255);
  nand GNAME3376(G3376,G1638,G3624);
  nand GNAME3377(G3377,G11132,G1690);
  nand GNAME3378(G3378,G3258,G1729);
  nand GNAME3379(G3379,G1631,G3255);
  nand GNAME3380(G3380,G1658,G3624);
  nand GNAME3381(G3381,G11117,G1690);
  nand GNAME3382(G3382,G3258,G1724);
  nand GNAME3383(G3383,G1658,G3255);
  or GNAME3384(G3384,G12083,G1693);
  nand GNAME3385(G3385,G3384,G1691);
  nand GNAME3386(G3386,G1692,G1695);
  nand GNAME3387(G3387,G11118,G1694);
  nand GNAME3388(G3388,G3386,G1753);
  nand GNAME3389(G3389,G1638,G3385);
  nand GNAME3390(G3390,G11119,G1694);
  nand GNAME3391(G3391,G3386,G1750);
  nand GNAME3392(G3392,G1630,G3385);
  nand GNAME3393(G3393,G11071,G1694);
  nand GNAME3394(G3394,G3386,G1747);
  nand GNAME3395(G3395,G1635,G3385);
  nand GNAME3396(G3396,G11070,G1694);
  nand GNAME3397(G3397,G3386,G1744);
  nand GNAME3398(G3398,G1634,G3385);
  nand GNAME3399(G3399,G11120,G1694);
  nand GNAME3400(G3400,G3386,G1741);
  nand GNAME3401(G3401,G1636,G3385);
  nand GNAME3402(G3402,G11121,G1694);
  nand GNAME3403(G3403,G3386,G1738);
  nand GNAME3404(G3404,G1632,G3385);
  nand GNAME3405(G3405,G11068,G1694);
  nand GNAME3406(G3406,G3386,G1591);
  nand GNAME3407(G3407,G1242,G3385);
  nand GNAME3408(G3408,G11067,G1694);
  nand GNAME3409(G3409,G3386,G1590);
  nand GNAME3410(G3410,G1244,G3385);
  nand GNAME3411(G3411,G11069,G1694);
  nand GNAME3412(G3412,G3386,G1735);
  nand GNAME3413(G3413,G1629,G3385);
  nand GNAME3414(G3414,G11122,G1694);
  nand GNAME3415(G3415,G3386,G1588);
  nand GNAME3416(G3416,G1641,G3385);
  nand GNAME3417(G3417,G11123,G1694);
  nand GNAME3418(G3418,G3386,G1587);
  nand GNAME3419(G3419,G1647,G3385);
  nand GNAME3420(G3420,G11124,G1694);
  nand GNAME3421(G3421,G3386,G1586);
  nand GNAME3422(G3422,G1646,G3385);
  nand GNAME3423(G3423,G11125,G1694);
  nand GNAME3424(G3424,G3386,G1585);
  nand GNAME3425(G3425,G1649,G3385);
  nand GNAME3426(G3426,G11126,G1694);
  nand GNAME3427(G3427,G3386,G1584);
  nand GNAME3428(G3428,G1642,G3385);
  nand GNAME3429(G3429,G11127,G1694);
  nand GNAME3430(G3430,G3386,G1583);
  nand GNAME3431(G3431,G1639,G3385);
  nand GNAME3432(G3432,G11128,G1694);
  nand GNAME3433(G3433,G3386,G1582);
  nand GNAME3434(G3434,G1643,G3385);
  nand GNAME3435(G3435,G11129,G1694);
  nand GNAME3436(G3436,G3386,G1581);
  nand GNAME3437(G3437,G1645,G3385);
  nand GNAME3438(G3438,G11130,G1694);
  nand GNAME3439(G3439,G3386,G1580);
  nand GNAME3440(G3440,G1640,G3385);
  nand GNAME3441(G3441,G11131,G1694);
  nand GNAME3442(G3442,G3386,G1579);
  nand GNAME3443(G3443,G1644,G3385);
  nand GNAME3444(G3444,G11066,G1694);
  nand GNAME3445(G3445,G3386,G1732);
  nand GNAME3446(G3446,G1633,G3385);
  nand GNAME3447(G3447,G11133,G1694);
  nand GNAME3448(G3448,G3386,G1782);
  nand GNAME3449(G3449,G1656,G3385);
  nand GNAME3450(G3450,G11134,G1694);
  nand GNAME3451(G3451,G3386,G1780);
  nand GNAME3452(G3452,G1657,G3385);
  nand GNAME3453(G3453,G11135,G1694);
  nand GNAME3454(G3454,G3386,G1777);
  nand GNAME3455(G3455,G1655,G3385);
  nand GNAME3456(G3456,G11136,G1694);
  nand GNAME3457(G3457,G3386,G1774);
  nand GNAME3458(G3458,G1653,G3385);
  nand GNAME3459(G3459,G11137,G1694);
  nand GNAME3460(G3460,G3386,G1771);
  nand GNAME3461(G3461,G1648,G3385);
  nand GNAME3462(G3462,G11065,G1694);
  nand GNAME3463(G3463,G3386,G1768);
  nand GNAME3464(G3464,G1651,G3385);
  nand GNAME3465(G3465,G11138,G1694);
  nand GNAME3466(G3466,G3386,G1765);
  nand GNAME3467(G3467,G1652,G3385);
  nand GNAME3468(G3468,G11139,G1694);
  nand GNAME3469(G3469,G3386,G1762);
  nand GNAME3470(G3470,G1654,G3385);
  nand GNAME3471(G3471,G11064,G1694);
  nand GNAME3472(G3472,G3386,G1759);
  nand GNAME3473(G3473,G1650,G3385);
  nand GNAME3474(G3474,G11063,G1694);
  nand GNAME3475(G3475,G3386,G1756);
  nand GNAME3476(G3476,G1637,G3385);
  nand GNAME3477(G3477,G11132,G1694);
  nand GNAME3478(G3478,G3386,G1729);
  nand GNAME3479(G3479,G1631,G3385);
  nand GNAME3480(G3480,G11117,G1694);
  nand GNAME3481(G3481,G3386,G1724);
  nand GNAME3482(G3482,G1658,G3385);
  nand GNAME3483(G3483,G1561,G1594);
  nand GNAME3484(G3484,G3646,G1701);
  nand GNAME3485(G3485,G1647,G1699);
  nand GNAME3486(G3486,G1641,G1700);
  nand GNAME3487(G3487,G1242,G1718);
  nand GNAME3488(G3488,G1244,G1718);
  nand GNAME3489(G3489,G1641,G1718);
  nand GNAME3490(G3490,G1698,G1704,G1697,G4161,G2022);
  or GNAME3491(G3491,G1682,G1699);
  nand GNAME3492(G3492,G3491,G1587);
  nand GNAME3493(G3493,G1700,G1588);
  nand GNAME3494(G3494,G1703,G1591);
  nand GNAME3495(G3495,G1703,G1590);
  nand GNAME3496(G3496,G1703,G1588);
  nand GNAME3497(G3497,G1701,G1704);
  or GNAME3498(G3498,G1708,G1709);
  or GNAME3499(G3499,G1688,G1689);
  nand GNAME3500(G3500,G3499,G1753);
  nand GNAME3501(G3501,G36078,G1706);
  nand GNAME3502(G3502,G36110,G1707);
  nand GNAME3503(G3503,G1638,G3498);
  nand GNAME3504(G3504,G3499,G1750);
  nand GNAME3505(G3505,G36077,G1706);
  nand GNAME3506(G3506,G36109,G1707);
  nand GNAME3507(G3507,G1630,G3498);
  nand GNAME3508(G3508,G3499,G1747);
  nand GNAME3509(G3509,G36076,G1706);
  nand GNAME3510(G3510,G36108,G1707);
  nand GNAME3511(G3511,G1635,G3498);
  nand GNAME3512(G3512,G3499,G1744);
  nand GNAME3513(G3513,G36075,G1706);
  nand GNAME3514(G3514,G36107,G1707);
  nand GNAME3515(G3515,G1634,G3498);
  nand GNAME3516(G3516,G3499,G1741);
  nand GNAME3517(G3517,G36074,G1706);
  nand GNAME3518(G3518,G36106,G1707);
  nand GNAME3519(G3519,G1636,G3498);
  nand GNAME3520(G3520,G3499,G1738);
  nand GNAME3521(G3521,G36073,G1706);
  nand GNAME3522(G3522,G36105,G1707);
  nand GNAME3523(G3523,G1632,G3498);
  nand GNAME3524(G3524,G36088,G1706);
  nand GNAME3525(G3525,G36120,G1707);
  nand GNAME3526(G3526,G1647,G3188);
  nand GNAME3527(G3527,G1688,G1587);
  nand GNAME3528(G3528,G1641,G3187);
  nand GNAME3529(G3529,G1689,G1588);
  nand GNAME3530(G3530,G1242,G1708);
  nand GNAME3531(G3531,G1244,G1708);
  nand GNAME3532(G3532,G3499,G1735);
  nand GNAME3533(G3533,G36072,G1706);
  nand GNAME3534(G3534,G36104,G1707);
  nand GNAME3535(G3535,G1629,G3498);
  nand GNAME3536(G3536,G1641,G1708);
  nand GNAME3537(G3537,G1647,G3498);
  nand GNAME3538(G3538,G3499,G1587);
  nand GNAME3539(G3539,G1646,G3498);
  nand GNAME3540(G3540,G3499,G1586);
  nand GNAME3541(G3541,G1649,G3498);
  nand GNAME3542(G3542,G3499,G1585);
  nand GNAME3543(G3543,G1642,G3498);
  nand GNAME3544(G3544,G3499,G1584);
  nand GNAME3545(G3545,G1639,G3498);
  nand GNAME3546(G3546,G3499,G1583);
  nand GNAME3547(G3547,G1643,G3498);
  nand GNAME3548(G3548,G3499,G1582);
  nand GNAME3549(G3549,G1645,G3498);
  nand GNAME3550(G3550,G3499,G1581);
  nand GNAME3551(G3551,G1640,G3498);
  nand GNAME3552(G3552,G3499,G1580);
  nand GNAME3553(G3553,G1644,G3498);
  nand GNAME3554(G3554,G3499,G1579);
  nand GNAME3555(G3555,G3499,G1732);
  nand GNAME3556(G3556,G36071,G1706);
  nand GNAME3557(G3557,G36103,G1707);
  nand GNAME3558(G3558,G1633,G3498);
  nand GNAME3559(G3559,G3499,G1782);
  nand GNAME3560(G3560,G1656,G3498);
  nand GNAME3561(G3561,G3499,G1780);
  nand GNAME3562(G3562,G36087,G1706);
  nand GNAME3563(G3563,G36119,G1707);
  nand GNAME3564(G3564,G1657,G3498);
  nand GNAME3565(G3565,G3499,G1777);
  nand GNAME3566(G3566,G36086,G1706);
  nand GNAME3567(G3567,G36118,G1707);
  nand GNAME3568(G3568,G1655,G3498);
  nand GNAME3569(G3569,G3499,G1774);
  nand GNAME3570(G3570,G36085,G1706);
  nand GNAME3571(G3571,G36117,G1707);
  nand GNAME3572(G3572,G1653,G3498);
  nand GNAME3573(G3573,G3499,G1771);
  nand GNAME3574(G3574,G36084,G1706);
  nand GNAME3575(G3575,G36116,G1707);
  nand GNAME3576(G3576,G1648,G3498);
  nand GNAME3577(G3577,G3499,G1768);
  nand GNAME3578(G3578,G36083,G1706);
  nand GNAME3579(G3579,G36115,G1707);
  nand GNAME3580(G3580,G1651,G3498);
  nand GNAME3581(G3581,G3499,G1765);
  nand GNAME3582(G3582,G36082,G1706);
  nand GNAME3583(G3583,G36114,G1707);
  nand GNAME3584(G3584,G1652,G3498);
  nand GNAME3585(G3585,G3499,G1762);
  nand GNAME3586(G3586,G36081,G1706);
  nand GNAME3587(G3587,G36113,G1707);
  nand GNAME3588(G3588,G1654,G3498);
  nand GNAME3589(G3589,G3499,G1759);
  nand GNAME3590(G3590,G36080,G1706);
  nand GNAME3591(G3591,G36112,G1707);
  nand GNAME3592(G3592,G1650,G3498);
  nand GNAME3593(G3593,G3499,G1756);
  nand GNAME3594(G3594,G36079,G1706);
  nand GNAME3595(G3595,G36111,G1707);
  nand GNAME3596(G3596,G1637,G3498);
  nand GNAME3597(G3597,G3499,G1729);
  nand GNAME3598(G3598,G36070,G1706);
  nand GNAME3599(G3599,G36102,G1707);
  nand GNAME3600(G3600,G1631,G3498);
  nand GNAME3601(G3601,G1722,G1624);
  nand GNAME3602(G3602,G3499,G1724);
  nand GNAME3603(G3603,G36069,G1706);
  nand GNAME3604(G3604,G36101,G1707);
  nand GNAME3605(G3605,G1658,G3498);
  nand GNAME3606(G3606,G1666,G1665);
  nand GNAME3607(G3607,G1665,G2017);
  nand GNAME3608(G3608,G2012,G2013,G1600,G1608,G2033);
  or GNAME3609(G3609,G1562,G1594,G1592);
  nand GNAME3610(G3610,G3606,G1671);
  nand GNAME3611(G3611,G2031,G3607);
  nand GNAME3612(G3612,G1662,G11853);
  nand GNAME3613(G3613,G1988,G35998);
  nand GNAME3614(G3614,G12026,G36004);
  nand GNAME3615(G3615,G1988,G35999);
  nand GNAME3616(G3616,G11995,G36004);
  nand GNAME3617(G3617,G3615,G3616);
  nand GNAME3618(G3618,G1988,G35997);
  nand GNAME3619(G3619,G12027,G36004);
  or GNAME3620(G3620,G36185,G4162,G1555);
  or GNAME3621(G3621,G1558,G1713,G1557);
  nand GNAME3622(G3622,G1988,G35996);
  nand GNAME3623(G3623,G11994,G36004);
  not GNAME3624(G3624,G1714);
  nand GNAME3625(G3625,G1989,G36005);
  nand GNAME3626(G3626,G2138,G2026);
  nand GNAME3627(G3627,G1989,G36006);
  nand GNAME3628(G3628,G2139,G2026);
  nand GNAME3629(G3629,G1988,G36002,G36003);
  nand GNAME3630(G3630,G36004,G11997,G12024);
  nand GNAME3631(G3631,G3629,G3630);
  nand GNAME3632(G3632,G1988,G1553,G36003);
  nand GNAME3633(G3633,G36004,G1552,G12024);
  nand GNAME3634(G3634,G3632,G3633);
  nand GNAME3635(G3635,G1988,G1554,G36002);
  or GNAME3636(G3636,G1988,G12024,G1552);
  nand GNAME3637(G3637,G3635,G3636);
  or GNAME3638(G3638,G36004,G36003,G36002);
  or GNAME3639(G3639,G1988,G11997,G12024);
  nand GNAME3640(G3640,G3638,G3639);
  nand GNAME3641(G3641,G1988,G36001);
  nand GNAME3642(G3642,G12025,G36004);
  not GNAME3643(G3643,G1717);
  nand GNAME3644(G3644,G1988,G35994);
  nand GNAME3645(G3645,G12028,G36004);
  not GNAME3646(G3646,G1718);
  nand GNAME3647(G3647,G1988,G35995);
  nand GNAME3648(G3648,G11993,G36004);
  not GNAME3649(G3649,G1719);
  nand GNAME3650(G3650,G1988,G35993);
  nand GNAME3651(G3651,G12029,G36004);
  not GNAME3652(G3652,G1720);
  nand GNAME3653(G3653,G1988,G35992);
  nand GNAME3654(G3654,G11992,G36004);
  not GNAME3655(G3655,G1721);
  nand GNAME3656(G3656,G1988,G35973);
  nand GNAME3657(G3657,G35973,G36004);
  nand GNAME3658(G3658,G1988,G36000);
  nand GNAME3659(G3659,G11996,G36004);
  not GNAME3660(G3660,G1723);
  nand GNAME3661(G3661,G2016,G889);
  nand GNAME3662(G3662,G1722,G1990);
  nand GNAME3663(G3663,G2136,G36005);
  nand GNAME3664(G3664,G1560,G2138);
  not GNAME3665(G3665,G1725);
  nand GNAME3666(G3666,G2136,G36006);
  nand GNAME3667(G3667,G1560,G2139);
  not GNAME3668(G3668,G1726);
  nand GNAME3669(G3669,G3649,G1718);
  nand GNAME3670(G3670,G3646,G1719);
  nand GNAME3671(G3671,G3669,G3670);
  nand GNAME3672(G3672,G1991,G36037);
  nand GNAME3673(G3673,G2158,G2027);
  nand GNAME3674(G3674,G1988,G35974);
  nand GNAME3675(G3675,G12017,G36004);
  nand GNAME3676(G3676,G2016,G878);
  nand GNAME3677(G3677,G1990,G1728);
  nand GNAME3678(G3678,G1991,G36038);
  nand GNAME3679(G3679,G2172,G2027);
  nand GNAME3680(G3680,G1988,G35975);
  nand GNAME3681(G3681,G11998,G36004);
  nand GNAME3682(G3682,G2016,G867);
  nand GNAME3683(G3683,G1990,G1731);
  nand GNAME3684(G3684,G1991,G36039);
  nand GNAME3685(G3685,G2182,G2027);
  nand GNAME3686(G3686,G1988,G35976);
  nand GNAME3687(G3687,G11999,G36004);
  nand GNAME3688(G3688,G2016,G864);
  nand GNAME3689(G3689,G1990,G1734);
  nand GNAME3690(G3690,G1991,G36040);
  nand GNAME3691(G3691,G2192,G2027);
  nand GNAME3692(G3692,G1988,G35977);
  nand GNAME3693(G3693,G12022,G36004);
  nand GNAME3694(G3694,G2016,G863);
  nand GNAME3695(G3695,G1990,G1737);
  nand GNAME3696(G3696,G1991,G36041);
  nand GNAME3697(G3697,G2202,G2027);
  nand GNAME3698(G3698,G1988,G35978);
  nand GNAME3699(G3699,G12021,G36004);
  nand GNAME3700(G3700,G2016,G862);
  nand GNAME3701(G3701,G1990,G1740);
  nand GNAME3702(G3702,G1991,G36042);
  nand GNAME3703(G3703,G2212,G2027);
  nand GNAME3704(G3704,G1988,G35979);
  nand GNAME3705(G3705,G12000,G36004);
  nand GNAME3706(G3706,G2016,G861);
  nand GNAME3707(G3707,G1990,G1743);
  nand GNAME3708(G3708,G1991,G36043);
  nand GNAME3709(G3709,G2222,G2027);
  nand GNAME3710(G3710,G1988,G35980);
  nand GNAME3711(G3711,G12001,G36004);
  nand GNAME3712(G3712,G2016,G860);
  nand GNAME3713(G3713,G1990,G1746);
  nand GNAME3714(G3714,G1991,G36044);
  nand GNAME3715(G3715,G2232,G2027);
  nand GNAME3716(G3716,G1988,G35981);
  nand GNAME3717(G3717,G12020,G36004);
  nand GNAME3718(G3718,G2016,G859);
  nand GNAME3719(G3719,G1990,G1749);
  nand GNAME3720(G3720,G1991,G36045);
  nand GNAME3721(G3721,G2242,G2027);
  nand GNAME3722(G3722,G1988,G35982);
  nand GNAME3723(G3723,G12019,G36004);
  nand GNAME3724(G3724,G2016,G858);
  nand GNAME3725(G3725,G1990,G1752);
  nand GNAME3726(G3726,G1991,G36046);
  nand GNAME3727(G3727,G2252,G2027);
  nand GNAME3728(G3728,G1988,G35983);
  nand GNAME3729(G3729,G11987,G36004);
  nand GNAME3730(G3730,G2016,G888);
  nand GNAME3731(G3731,G1990,G1755);
  nand GNAME3732(G3732,G1991,G36047);
  nand GNAME3733(G3733,G2262,G2027);
  nand GNAME3734(G3734,G1988,G35984);
  nand GNAME3735(G3735,G11988,G36004);
  nand GNAME3736(G3736,G2016,G887);
  nand GNAME3737(G3737,G1990,G1758);
  nand GNAME3738(G3738,G1991,G36048);
  nand GNAME3739(G3739,G2272,G2027);
  nand GNAME3740(G3740,G1988,G35985);
  nand GNAME3741(G3741,G12034,G36004);
  nand GNAME3742(G3742,G2016,G886);
  nand GNAME3743(G3743,G1990,G1761);
  nand GNAME3744(G3744,G1991,G36049);
  nand GNAME3745(G3745,G2282,G2027);
  nand GNAME3746(G3746,G1988,G35986);
  nand GNAME3747(G3747,G12033,G36004);
  nand GNAME3748(G3748,G2016,G885);
  nand GNAME3749(G3749,G1990,G1764);
  nand GNAME3750(G3750,G1991,G36050);
  nand GNAME3751(G3751,G2292,G2027);
  nand GNAME3752(G3752,G1988,G35987);
  nand GNAME3753(G3753,G11989,G36004);
  nand GNAME3754(G3754,G2016,G884);
  nand GNAME3755(G3755,G1990,G1767);
  nand GNAME3756(G3756,G1991,G36051);
  nand GNAME3757(G3757,G2302,G2027);
  nand GNAME3758(G3758,G1988,G35988);
  nand GNAME3759(G3759,G11990,G36004);
  nand GNAME3760(G3760,G2016,G883);
  nand GNAME3761(G3761,G1990,G1770);
  nand GNAME3762(G3762,G1991,G36052);
  nand GNAME3763(G3763,G2312,G2027);
  nand GNAME3764(G3764,G1988,G35989);
  nand GNAME3765(G3765,G12032,G36004);
  nand GNAME3766(G3766,G2016,G882);
  nand GNAME3767(G3767,G1990,G1773);
  nand GNAME3768(G3768,G1991,G36053);
  nand GNAME3769(G3769,G2322,G2027);
  nand GNAME3770(G3770,G1988,G35990);
  nand GNAME3771(G3771,G12031,G36004);
  nand GNAME3772(G3772,G2016,G881);
  nand GNAME3773(G3773,G1990,G1776);
  nand GNAME3774(G3774,G1991,G36054);
  nand GNAME3775(G3775,G2332,G2027);
  nand GNAME3776(G3776,G1988,G35991);
  nand GNAME3777(G3777,G11991,G36004);
  nand GNAME3778(G3778,G2016,G880);
  nand GNAME3779(G3779,G1990,G1779);
  nand GNAME3780(G3780,G1991,G36055);
  nand GNAME3781(G3781,G2342,G2027);
  nand GNAME3782(G3782,G2016,G879);
  nand GNAME3783(G3783,G1721,G1990);
  nand GNAME3784(G3784,G1991,G36056);
  nand GNAME3785(G3785,G2352,G2027);
  nand GNAME3786(G3786,G1991,G36057);
  nand GNAME3787(G3787,G2362,G2027);
  nand GNAME3788(G3788,G1991,G36058);
  nand GNAME3789(G3789,G2372,G2027);
  nand GNAME3790(G3790,G1991,G36059);
  nand GNAME3791(G3791,G2382,G2027);
  nand GNAME3792(G3792,G1991,G36060);
  nand GNAME3793(G3793,G2392,G2027);
  nand GNAME3794(G3794,G1991,G36061);
  nand GNAME3795(G3795,G2402,G2027);
  nand GNAME3796(G3796,G1991,G36062);
  nand GNAME3797(G3797,G2412,G2027);
  nand GNAME3798(G3798,G1991,G36063);
  nand GNAME3799(G3799,G2422,G2027);
  nand GNAME3800(G3800,G1991,G36064);
  nand GNAME3801(G3801,G2432,G2027);
  nand GNAME3802(G3802,G1991,G36065);
  nand GNAME3803(G3803,G2442,G2027);
  nand GNAME3804(G3804,G1991,G36066);
  nand GNAME3805(G3805,G2455,G2027);
  nand GNAME3806(G3806,G1991,G36067);
  nand GNAME3807(G3807,G2461,G2027);
  nand GNAME3808(G3808,G1991,G36068);
  nand GNAME3809(G3809,G2464,G2027);
  nand GNAME3810(G3810,G1992,G36069);
  nand GNAME3811(G3811,G2158,G2028);
  nand GNAME3812(G3812,G1992,G36070);
  nand GNAME3813(G3813,G2172,G2028);
  nand GNAME3814(G3814,G1992,G36071);
  nand GNAME3815(G3815,G2182,G2028);
  nand GNAME3816(G3816,G1992,G36072);
  nand GNAME3817(G3817,G2192,G2028);
  nand GNAME3818(G3818,G1992,G36073);
  nand GNAME3819(G3819,G2202,G2028);
  nand GNAME3820(G3820,G1992,G36074);
  nand GNAME3821(G3821,G2212,G2028);
  nand GNAME3822(G3822,G1992,G36075);
  nand GNAME3823(G3823,G2222,G2028);
  nand GNAME3824(G3824,G1992,G36076);
  nand GNAME3825(G3825,G2232,G2028);
  nand GNAME3826(G3826,G1992,G36077);
  nand GNAME3827(G3827,G2242,G2028);
  nand GNAME3828(G3828,G1992,G36078);
  nand GNAME3829(G3829,G2252,G2028);
  nand GNAME3830(G3830,G1992,G36079);
  nand GNAME3831(G3831,G2262,G2028);
  nand GNAME3832(G3832,G1992,G36080);
  nand GNAME3833(G3833,G2272,G2028);
  nand GNAME3834(G3834,G1992,G36081);
  nand GNAME3835(G3835,G2282,G2028);
  nand GNAME3836(G3836,G1992,G36082);
  nand GNAME3837(G3837,G2292,G2028);
  nand GNAME3838(G3838,G1992,G36083);
  nand GNAME3839(G3839,G2302,G2028);
  nand GNAME3840(G3840,G1992,G36084);
  nand GNAME3841(G3841,G2312,G2028);
  nand GNAME3842(G3842,G1992,G36085);
  nand GNAME3843(G3843,G2322,G2028);
  nand GNAME3844(G3844,G1992,G36086);
  nand GNAME3845(G3845,G2332,G2028);
  nand GNAME3846(G3846,G1992,G36087);
  nand GNAME3847(G3847,G2342,G2028);
  nand GNAME3848(G3848,G1992,G36088);
  nand GNAME3849(G3849,G2352,G2028);
  nand GNAME3850(G3850,G1992,G36089);
  nand GNAME3851(G3851,G2362,G2028);
  nand GNAME3852(G3852,G1992,G36090);
  nand GNAME3853(G3853,G2372,G2028);
  nand GNAME3854(G3854,G1992,G36091);
  nand GNAME3855(G3855,G2382,G2028);
  nand GNAME3856(G3856,G1992,G36092);
  nand GNAME3857(G3857,G2392,G2028);
  nand GNAME3858(G3858,G1992,G36093);
  nand GNAME3859(G3859,G2402,G2028);
  nand GNAME3860(G3860,G1992,G36094);
  nand GNAME3861(G3861,G2412,G2028);
  nand GNAME3862(G3862,G1992,G36095);
  nand GNAME3863(G3863,G2422,G2028);
  nand GNAME3864(G3864,G1992,G36096);
  nand GNAME3865(G3865,G2432,G2028);
  nand GNAME3866(G3866,G1992,G36097);
  nand GNAME3867(G3867,G2442,G2028);
  nand GNAME3868(G3868,G1992,G36098);
  nand GNAME3869(G3869,G2455,G2028);
  nand GNAME3870(G3870,G1992,G36099);
  nand GNAME3871(G3871,G2461,G2028);
  nand GNAME3872(G3872,G1992,G36100);
  nand GNAME3873(G3873,G2464,G2028);
  nand GNAME3874(G3874,G1596,G36102);
  nand GNAME3875(G3875,G2485,G2029);
  nand GNAME3876(G3876,G1596,G36130);
  nand GNAME3877(G3877,G2029,G2450,G1565);
  nand GNAME3878(G3878,G1596,G36131);
  nand GNAME3879(G3879,G2680,G2029);
  nand GNAME3880(G3880,G1596,G36132);
  nand GNAME3881(G3881,G2683,G2029);
  nand GNAME3882(G3882,G2025,G36153);
  nand GNAME3883(G3883,G1658,G1625);
  nand GNAME3884(G3884,G2025,G36154);
  nand GNAME3885(G3885,G1631,G1625);
  nand GNAME3886(G3886,G2025,G36155);
  nand GNAME3887(G3887,G1633,G1625);
  nand GNAME3888(G3888,G2025,G36156);
  nand GNAME3889(G3889,G1629,G1625);
  nand GNAME3890(G3890,G2025,G36157);
  nand GNAME3891(G3891,G1632,G1625);
  nand GNAME3892(G3892,G2025,G36158);
  nand GNAME3893(G3893,G1636,G1625);
  nand GNAME3894(G3894,G2025,G36159);
  nand GNAME3895(G3895,G1634,G1625);
  nand GNAME3896(G3896,G2025,G36160);
  nand GNAME3897(G3897,G1635,G1625);
  nand GNAME3898(G3898,G2025,G36161);
  nand GNAME3899(G3899,G1630,G1625);
  nand GNAME3900(G3900,G2025,G36162);
  nand GNAME3901(G3901,G1638,G1625);
  nand GNAME3902(G3902,G2025,G36163);
  nand GNAME3903(G3903,G1637,G1625);
  nand GNAME3904(G3904,G2025,G36164);
  nand GNAME3905(G3905,G1650,G1625);
  nand GNAME3906(G3906,G2025,G36165);
  nand GNAME3907(G3907,G1654,G1625);
  nand GNAME3908(G3908,G2025,G36166);
  nand GNAME3909(G3909,G1652,G1625);
  nand GNAME3910(G3910,G2025,G36167);
  nand GNAME3911(G3911,G1651,G1625);
  nand GNAME3912(G3912,G2025,G36168);
  nand GNAME3913(G3913,G1648,G1625);
  nand GNAME3914(G3914,G2025,G36169);
  nand GNAME3915(G3915,G1653,G1625);
  nand GNAME3916(G3916,G2025,G36170);
  nand GNAME3917(G3917,G1655,G1625);
  nand GNAME3918(G3918,G2025,G36171);
  nand GNAME3919(G3919,G1657,G1625);
  nand GNAME3920(G3920,G2025,G36172);
  nand GNAME3921(G3921,G1656,G1625);
  nand GNAME3922(G3922,G2025,G36173);
  nand GNAME3923(G3923,G1644,G1625);
  nand GNAME3924(G3924,G2025,G36174);
  nand GNAME3925(G3925,G1640,G1625);
  nand GNAME3926(G3926,G2025,G36175);
  nand GNAME3927(G3927,G1645,G1625);
  nand GNAME3928(G3928,G2025,G36176);
  nand GNAME3929(G3929,G1643,G1625);
  nand GNAME3930(G3930,G2025,G36177);
  nand GNAME3931(G3931,G1639,G1625);
  nand GNAME3932(G3932,G2025,G36178);
  nand GNAME3933(G3933,G1642,G1625);
  nand GNAME3934(G3934,G2025,G36179);
  nand GNAME3935(G3935,G1649,G1625);
  nand GNAME3936(G3936,G2025,G36180);
  nand GNAME3937(G3937,G1646,G1625);
  nand GNAME3938(G3938,G2025,G36181);
  nand GNAME3939(G3939,G1647,G1625);
  nand GNAME3940(G3940,G2025,G36182);
  nand GNAME3941(G3941,G1641,G1625);
  nand GNAME3942(G3942,G2025,G36183);
  nand GNAME3943(G3943,G1244,G1625);
  nand GNAME3944(G3944,G2025,G36184);
  nand GNAME3945(G3945,G1242,G1625);
  or GNAME3946(G3946,G1631,G1729);
  nand GNAME3947(G3947,G1631,G1729);
  nand GNAME3948(G3948,G3946,G3947);
  or GNAME3949(G3949,G1629,G1735);
  nand GNAME3950(G3950,G1629,G1735);
  nand GNAME3951(G3951,G3949,G3950);
  or GNAME3952(G3952,G1630,G1750);
  nand GNAME3953(G3953,G1630,G1750);
  nand GNAME3954(G3954,G3952,G3953);
  or GNAME3955(G3955,G1632,G1738);
  nand GNAME3956(G3956,G1632,G1738);
  nand GNAME3957(G3957,G3955,G3956);
  or GNAME3958(G3958,G1633,G1732);
  nand GNAME3959(G3959,G1633,G1732);
  nand GNAME3960(G3960,G3958,G3959);
  or GNAME3961(G3961,G1636,G1741);
  nand GNAME3962(G3962,G1636,G1741);
  nand GNAME3963(G3963,G3961,G3962);
  or GNAME3964(G3964,G1634,G1744);
  nand GNAME3965(G3965,G1634,G1744);
  nand GNAME3966(G3966,G3964,G3965);
  or GNAME3967(G3967,G1635,G1747);
  nand GNAME3968(G3968,G1635,G1747);
  nand GNAME3969(G3969,G3967,G3968);
  or GNAME3970(G3970,G1637,G1756);
  nand GNAME3971(G3971,G1637,G1756);
  nand GNAME3972(G3972,G3970,G3971);
  or GNAME3973(G3973,G1638,G1753);
  nand GNAME3974(G3974,G1638,G1753);
  nand GNAME3975(G3975,G3973,G3974);
  nand GNAME3976(G3976,G1640,G1580);
  or GNAME3977(G3977,G1580,G1640);
  nand GNAME3978(G3978,G3976,G3977);
  nand GNAME3979(G3979,G1639,G1583);
  or GNAME3980(G3980,G1583,G1639);
  nand GNAME3981(G3981,G3979,G3980);
  nand GNAME3982(G3982,G1244,G1590);
  or GNAME3983(G3983,G1244,G1590);
  nand GNAME3984(G3984,G3982,G3983);
  nand GNAME3985(G3985,G1643,G1582);
  or GNAME3986(G3986,G1582,G1643);
  nand GNAME3987(G3987,G3985,G3986);
  nand GNAME3988(G3988,G1641,G1588);
  or GNAME3989(G3989,G1588,G1641);
  nand GNAME3990(G3990,G3988,G3989);
  nand GNAME3991(G3991,G1642,G1584);
  or GNAME3992(G3992,G1584,G1642);
  nand GNAME3993(G3993,G3991,G3992);
  nand GNAME3994(G3994,G1646,G1586);
  or GNAME3995(G3995,G1586,G1646);
  nand GNAME3996(G3996,G3994,G3995);
  nand GNAME3997(G3997,G1644,G1579);
  or GNAME3998(G3998,G1579,G1644);
  nand GNAME3999(G3999,G3997,G3998);
  nand GNAME4000(G4000,G1645,G1581);
  or GNAME4001(G4001,G1581,G1645);
  nand GNAME4002(G4002,G4000,G4001);
  nand GNAME4003(G4003,G1242,G1591);
  or GNAME4004(G4004,G1242,G1591);
  nand GNAME4005(G4005,G4003,G4004);
  nand GNAME4006(G4006,G1647,G1587);
  or GNAME4007(G4007,G1587,G1647);
  nand GNAME4008(G4008,G4006,G4007);
  or GNAME4009(G4009,G1650,G1759);
  nand GNAME4010(G4010,G1650,G1759);
  nand GNAME4011(G4011,G4009,G4010);
  nand GNAME4012(G4012,G1649,G1585);
  or GNAME4013(G4013,G1585,G1649);
  nand GNAME4014(G4014,G4012,G4013);
  or GNAME4015(G4015,G1648,G1771);
  nand GNAME4016(G4016,G1648,G1771);
  nand GNAME4017(G4017,G4015,G4016);
  or GNAME4018(G4018,G1651,G1768);
  nand GNAME4019(G4019,G1651,G1768);
  nand GNAME4020(G4020,G4018,G4019);
  or GNAME4021(G4021,G1652,G1765);
  nand GNAME4022(G4022,G1652,G1765);
  nand GNAME4023(G4023,G4021,G4022);
  or GNAME4024(G4024,G1655,G1777);
  nand GNAME4025(G4025,G1655,G1777);
  nand GNAME4026(G4026,G4024,G4025);
  or GNAME4027(G4027,G1653,G1774);
  nand GNAME4028(G4028,G1653,G1774);
  nand GNAME4029(G4029,G4027,G4028);
  or GNAME4030(G4030,G1654,G1762);
  nand GNAME4031(G4031,G1654,G1762);
  nand GNAME4032(G4032,G4030,G4031);
  or GNAME4033(G4033,G1656,G1782);
  nand GNAME4034(G4034,G1656,G1782);
  nand GNAME4035(G4035,G4033,G4034);
  or GNAME4036(G4036,G1657,G1780);
  nand GNAME4037(G4037,G1657,G1780);
  nand GNAME4038(G4038,G4036,G4037);
  or GNAME4039(G4039,G1658,G1724);
  nand GNAME4040(G4040,G1658,G1724);
  nand GNAME4041(G4041,G4039,G4040);
  nand GNAME4042(G4042,G1611,G11853);
  nand GNAME4043(G4043,G1663,G1661);
  nand GNAME4044(G4044,G4042,G4043);
  nand GNAME4045(G4045,G1718,G1663,G1611);
  nand GNAME4046(G4046,G3646,G4044);
  or GNAME4047(G4047,G11853,G1604,G3624,G1719);
  nand GNAME4048(G4048,G11853,G1718,G1661);
  nand GNAME4049(G4049,G1663,G12307);
  nand GNAME4050(G4050,G1638,G11853);
  nand GNAME4051(G4051,G1663,G12309);
  nand GNAME4052(G4052,G1630,G11853);
  nand GNAME4053(G4053,G1663,G12311);
  nand GNAME4054(G4054,G1635,G11853);
  nand GNAME4055(G4055,G1663,G12313);
  nand GNAME4056(G4056,G1634,G11853);
  nand GNAME4057(G4057,G1663,G12315);
  nand GNAME4058(G4058,G1636,G11853);
  nand GNAME4059(G4059,G1663,G12317);
  nand GNAME4060(G4060,G1632,G11853);
  nand GNAME4061(G4061,G1663,G12319);
  nand GNAME4062(G4062,G1629,G11853);
  nand GNAME4063(G4063,G1663,G12211);
  nand GNAME4064(G4064,G1242,G11853);
  nand GNAME4065(G4065,G1663,G12322);
  nand GNAME4066(G4066,G1244,G11853);
  nand GNAME4067(G4067,G1663,G12324);
  nand GNAME4068(G4068,G1633,G11853);
  nand GNAME4069(G4069,G1663,G12326);
  nand GNAME4070(G4070,G1641,G11853);
  nand GNAME4071(G4071,G1663,G12328);
  nand GNAME4072(G4072,G1647,G11853);
  nand GNAME4073(G4073,G1663,G12330);
  nand GNAME4074(G4074,G1646,G11853);
  nand GNAME4075(G4075,G1663,G12332);
  nand GNAME4076(G4076,G1649,G11853);
  nand GNAME4077(G4077,G1663,G12334);
  nand GNAME4078(G4078,G1642,G11853);
  nand GNAME4079(G4079,G1663,G12336);
  nand GNAME4080(G4080,G1639,G11853);
  nand GNAME4081(G4081,G1663,G12338);
  nand GNAME4082(G4082,G1643,G11853);
  nand GNAME4083(G4083,G1663,G12340);
  nand GNAME4084(G4084,G1645,G11853);
  nand GNAME4085(G4085,G1663,G12342);
  nand GNAME4086(G4086,G1640,G11853);
  nand GNAME4087(G4087,G1663,G12344);
  nand GNAME4088(G4088,G1644,G11853);
  nand GNAME4089(G4089,G1663,G12275);
  nand GNAME4090(G4090,G1631,G11853);
  nand GNAME4091(G4091,G1663,G12347);
  nand GNAME4092(G4092,G1656,G11853);
  nand GNAME4093(G4093,G1663,G12349);
  nand GNAME4094(G4094,G1657,G11853);
  nand GNAME4095(G4095,G1663,G12351);
  nand GNAME4096(G4096,G1655,G11853);
  nand GNAME4097(G4097,G1663,G12353);
  nand GNAME4098(G4098,G1653,G11853);
  nand GNAME4099(G4099,G1663,G12355);
  nand GNAME4100(G4100,G1648,G11853);
  nand GNAME4101(G4101,G1663,G12357);
  nand GNAME4102(G4102,G1651,G11853);
  nand GNAME4103(G4103,G1663,G12359);
  nand GNAME4104(G4104,G1652,G11853);
  nand GNAME4105(G4105,G1663,G12361);
  nand GNAME4106(G4106,G1654,G11853);
  nand GNAME4107(G4107,G1663,G12363);
  nand GNAME4108(G4108,G1650,G11853);
  nand GNAME4109(G4109,G1663,G12365);
  nand GNAME4110(G4110,G1637,G11853);
  nand GNAME4111(G4111,G1663,G12212);
  nand GNAME4112(G4112,G1658,G11853);
  nand GNAME4113(G4113,G3643,G1722);
  nand GNAME4114(G4114,G11117,G1717);
  nand GNAME4115(G4115,G1575,G1723);
  nand GNAME4116(G4116,G1576,G3660);
  or GNAME4117(G4117,G1567,G1718);
  nand GNAME4118(G4118,G3652,G1718);
  nand GNAME4119(G4119,G36110,G1723);
  nand GNAME4120(G4120,G36078,G3660);
  nand GNAME4121(G4121,G36109,G1723);
  nand GNAME4122(G4122,G36077,G3660);
  nand GNAME4123(G4123,G36108,G1723);
  nand GNAME4124(G4124,G36076,G3660);
  nand GNAME4125(G4125,G36107,G1723);
  nand GNAME4126(G4126,G36075,G3660);
  nand GNAME4127(G4127,G36106,G1723);
  nand GNAME4128(G4128,G36074,G3660);
  nand GNAME4129(G4129,G36105,G1723);
  nand GNAME4130(G4130,G36073,G3660);
  nand GNAME4131(G4131,G36104,G1723);
  nand GNAME4132(G4132,G36072,G3660);
  nand GNAME4133(G4133,G36103,G1723);
  nand GNAME4134(G4134,G36071,G3660);
  nand GNAME4135(G4135,G36120,G1723);
  nand GNAME4136(G4136,G36088,G3660);
  nand GNAME4137(G4137,G36119,G1723);
  nand GNAME4138(G4138,G36087,G3660);
  nand GNAME4139(G4139,G36118,G1723);
  nand GNAME4140(G4140,G36086,G3660);
  nand GNAME4141(G4141,G36117,G1723);
  nand GNAME4142(G4142,G36085,G3660);
  nand GNAME4143(G4143,G36116,G1723);
  nand GNAME4144(G4144,G36084,G3660);
  nand GNAME4145(G4145,G36115,G1723);
  nand GNAME4146(G4146,G36083,G3660);
  nand GNAME4147(G4147,G36114,G1723);
  nand GNAME4148(G4148,G36082,G3660);
  nand GNAME4149(G4149,G36113,G1723);
  nand GNAME4150(G4150,G36081,G3660);
  nand GNAME4151(G4151,G36112,G1723);
  nand GNAME4152(G4152,G36080,G3660);
  nand GNAME4153(G4153,G36111,G1723);
  nand GNAME4154(G4154,G36079,G3660);
  nand GNAME4155(G4155,G36102,G1723);
  nand GNAME4156(G4156,G36070,G3660);
  nand GNAME4157(G4157,G36101,G1723);
  nand GNAME4158(G4158,G36069,G3660);
  not GNAME4159(G4159,G12083);
  not GNAME4160(G4160,G1605);
  not GNAME4161(G4161,G1687);
  not GNAME4162(G4162,G1712);
  or GNAME4163(G4163,G7754,G15018);
  nand GNAME4164(G4164,G4165,G4167,G4166);
  nand GNAME4165(G4165,G15018,G7754);
  or GNAME4166(G4166,G7570,G15017);
  nand GNAME4167(G4167,G4168,G4170,G4169);
  nand GNAME4168(G4168,G15017,G7570);
  or GNAME4169(G4169,G7756,G15016);
  nand GNAME4170(G4170,G4171,G4173,G4172);
  nand GNAME4171(G4171,G15016,G7756);
  or GNAME4172(G4172,G7568,G15015);
  nand GNAME4173(G4173,G7126,G7128,G7127);
  or GNAME4174(G4174,G4661,G4691,G4665,G6248);
  or GNAME4175(G4175,G4176,G4691);
  nand GNAME4176(G4176,G6159,G6160,G6158,G4974,G6157);
  nand GNAME4177(G4177,G6167,G4974,G6166);
  nand GNAME4178(G4178,G6169,G4974,G6168);
  nand GNAME4179(G4179,G6171,G4974,G6170);
  nand GNAME4180(G4180,G6173,G4974,G6172);
  nand GNAME4181(G4181,G6175,G4974,G6174);
  nand GNAME4182(G4182,G6177,G4974,G6176);
  nand GNAME4183(G4183,G6179,G4974,G6178);
  nand GNAME4184(G4184,G6181,G4974,G6180);
  nand GNAME4185(G4185,G6183,G4974,G6182);
  nand GNAME4186(G4186,G6191,G6192,G6190,G4974,G6189);
  nand GNAME4187(G4187,G6196,G6197,G6195,G6193,G6194);
  nand GNAME4188(G4188,G6201,G6202,G6200,G6198,G6199);
  nand GNAME4189(G4189,G6206,G6207,G6205,G6203,G6204);
  nand GNAME4190(G4190,G6211,G6212,G6210,G6208,G6209);
  nand GNAME4191(G4191,G6216,G6217,G6215,G6213,G6214);
  nand GNAME4192(G4192,G6221,G6222,G6220,G6218,G6219);
  nand GNAME4193(G4193,G6226,G6227,G6225,G6223,G6224);
  nand GNAME4194(G4194,G6231,G6232,G6230,G6228,G6229);
  nand GNAME4195(G4195,G6236,G6237,G6235,G6233,G6234);
  nand GNAME4196(G4196,G6128,G6129,G6127,G6125,G6126);
  nand GNAME4197(G4197,G6133,G6134,G6132,G6130,G6131);
  nand GNAME4198(G4198,G6138,G6139,G6137,G6135,G6136);
  nand GNAME4199(G4199,G6143,G6144,G6142,G6140,G6141);
  nand GNAME4200(G4200,G6148,G6149,G6147,G6145,G6146);
  nand GNAME4201(G4201,G6153,G6154,G6152,G6150,G6151);
  nand GNAME4202(G4202,G6164,G6165,G6163,G6161,G6162);
  nand GNAME4203(G4203,G6187,G6188,G6186,G6184,G6185);
  nand GNAME4204(G4204,G6241,G6242,G6240,G6238,G6239);
  nand GNAME4205(G4205,G6246,G6247,G6245,G6243,G6244);
  nand GNAME4206(G4206,G6592,G4688);
  nand GNAME4207(G4207,G5399,G5397,G5398);
  nand GNAME4208(G4208,G6593,G4688);
  nand GNAME4209(G4209,G5386,G5384,G5385);
  nand GNAME4210(G4210,G6599,G4688);
  nand GNAME4211(G4211,G4687,G6600,G6601);
  nand GNAME4212(G4212,G4687,G6602,G6603);
  nand GNAME4213(G4213,G4687,G6604,G6605);
  nand GNAME4214(G4214,G4687,G6606,G6607);
  nand GNAME4215(G4215,G4687,G6608,G6609);
  nand GNAME4216(G4216,G4687,G6610,G6611);
  nand GNAME4217(G4217,G4687,G6612,G6613);
  nand GNAME4218(G4218,G4687,G6614,G6615);
  nand GNAME4219(G4219,G4687,G6616,G6617);
  nand GNAME4220(G4220,G6623,G6624,G6625,G4687);
  nand GNAME4221(G4221,G6629,G6630,G6628,G6626,G6627);
  nand GNAME4222(G4222,G6634,G6635,G6633,G6631,G6632);
  nand GNAME4223(G4223,G6639,G6640,G6638,G6636,G6637);
  nand GNAME4224(G4224,G6644,G6645,G6643,G6641,G6642);
  nand GNAME4225(G4225,G6649,G6650,G6648,G6646,G6647);
  nand GNAME4226(G4226,G6654,G6655,G6653,G6651,G6652);
  nand GNAME4227(G4227,G6659,G6660,G6658,G6656,G6657);
  nand GNAME4228(G4228,G6664,G6665,G6663,G6661,G6662);
  nand GNAME4229(G4229,G6669,G6670,G6668,G6666,G6667);
  nand GNAME4230(G4230,G6559,G6560,G6558,G6556,G6557);
  nand GNAME4231(G4231,G6564,G6565,G6563,G6561,G6562);
  nand GNAME4232(G4232,G6569,G6570,G6568,G6566,G6567);
  nand GNAME4233(G4233,G6574,G6575,G6573,G6571,G6572);
  nand GNAME4234(G4234,G6579,G6580,G6578,G6576,G6577);
  nand GNAME4235(G4235,G6584,G6585,G6583,G6581,G6582);
  nand GNAME4236(G4236,G6597,G6598,G6596,G6594,G6595);
  nand GNAME4237(G4237,G6621,G6622,G6620,G6618,G6619);
  nand GNAME4238(G4238,G6674,G6675,G6673,G6671,G6672);
  nand GNAME4239(G4239,G6679,G6680,G6678,G6676,G6677);
  nand GNAME4240(G4240,G6700,G4604);
  nand GNAME4241(G4241,G4551,G4555,G4691,G4645);
  nand GNAME4242(G4242,G6478,G6476,G6477);
  nand GNAME4243(G4243,G6481,G6479,G6480);
  nand GNAME4244(G4244,G6485,G6486,G6487,G4691);
  nand GNAME4245(G4245,G6488,G6489,G6490,G4691);
  nand GNAME4246(G4246,G6491,G6492,G6493,G4691);
  nand GNAME4247(G4247,G6494,G6495,G6496,G4691);
  nand GNAME4248(G4248,G6497,G6498,G6499,G4691);
  nand GNAME4249(G4249,G6500,G6501,G6502,G4691);
  nand GNAME4250(G4250,G6503,G6504,G6505,G4691);
  nand GNAME4251(G4251,G6506,G6507,G6508,G4691);
  nand GNAME4252(G4252,G6509,G6510,G6511,G4691);
  nand GNAME4253(G4253,G6512,G6513,G6514,G4691);
  nand GNAME4254(G4254,G6518,G6519,G6520,G4691);
  nand GNAME4255(G4255,G6521,G6522,G6523,G4691);
  nand GNAME4256(G4256,G6524,G6525,G6526,G4691);
  nand GNAME4257(G4257,G6527,G6528,G6529,G4691);
  nand GNAME4258(G4258,G6530,G6531,G6532,G4691);
  nand GNAME4259(G4259,G6533,G6534,G6535,G4691);
  nand GNAME4260(G4260,G6536,G6537,G6538,G4691);
  nand GNAME4261(G4261,G6539,G6540,G6541,G4691);
  nand GNAME4262(G4262,G6542,G6543,G6544,G4691);
  nand GNAME4263(G4263,G6545,G6546,G6547,G4691);
  nand GNAME4264(G4264,G6458,G6459,G6460,G4691);
  nand GNAME4265(G4265,G6461,G6462,G6463,G4691);
  nand GNAME4266(G4266,G6464,G6465,G6466,G4691);
  nand GNAME4267(G4267,G6467,G6468,G6469,G4691);
  nand GNAME4268(G4268,G6470,G6471,G6472,G4691);
  nand GNAME4269(G4269,G6473,G6474,G6475,G4691);
  nand GNAME4270(G4270,G6482,G6483,G6484,G4691);
  nand GNAME4271(G4271,G6515,G6516,G6517,G4691);
  nand GNAME4272(G4272,G6548,G6549,G6550,G4691);
  nand GNAME4273(G4273,G6551,G6552,G6553,G4691);
  nand GNAME4274(G4274,G6381,G6382);
  nand GNAME4275(G4275,G6383,G6384);
  nand GNAME4276(G4276,G6390,G6388,G6389);
  nand GNAME4277(G4277,G6393,G6391,G6392);
  nand GNAME4278(G4278,G6396,G6394,G6395);
  nand GNAME4279(G4279,G6399,G6397,G6398);
  nand GNAME4280(G4280,G6402,G6400,G6401);
  nand GNAME4281(G4281,G6405,G6403,G6404);
  nand GNAME4282(G4282,G6408,G6406,G6407);
  nand GNAME4283(G4283,G6411,G6409,G6410);
  nand GNAME4284(G4284,G6414,G6412,G6413);
  nand GNAME4285(G4285,G6417,G6415,G6416);
  nand GNAME4286(G4286,G6423,G6421,G6422);
  nand GNAME4287(G4287,G6426,G6424,G6425);
  nand GNAME4288(G4288,G6429,G6427,G6428);
  nand GNAME4289(G4289,G6432,G6430,G6431);
  nand GNAME4290(G4290,G6435,G6433,G6434);
  nand GNAME4291(G4291,G6438,G6436,G6437);
  nand GNAME4292(G4292,G6441,G6439,G6440);
  nand GNAME4293(G4293,G6444,G6442,G6443);
  nand GNAME4294(G4294,G6447,G6445,G6446);
  nand GNAME4295(G4295,G6450,G6448,G6449);
  nand GNAME4296(G4296,G6365,G6363,G6364);
  nand GNAME4297(G4297,G6368,G6366,G6367);
  nand GNAME4298(G4298,G6371,G6369,G6370);
  nand GNAME4299(G4299,G6374,G6372,G6373);
  nand GNAME4300(G4300,G6377,G6375,G6376);
  nand GNAME4301(G4301,G6380,G6378,G6379);
  nand GNAME4302(G4302,G6387,G6385,G6386);
  nand GNAME4303(G4303,G6420,G6418,G6419);
  nand GNAME4304(G4304,G6453,G6451,G6452);
  nand GNAME4305(G4305,G6454,G6455);
  nand GNAME4306(G4306,G6335,G6336);
  nand GNAME4307(G4307,G6337,G6338);
  nand GNAME4308(G4308,G6339,G6340);
  nand GNAME4309(G4309,G6341,G6342);
  nand GNAME4310(G4310,G6343,G6344);
  nand GNAME4311(G4311,G6345,G6346);
  nand GNAME4312(G4312,G6347,G6348);
  nand GNAME4313(G4313,G6349,G6350);
  nand GNAME4314(G4314,G6351,G6352);
  nand GNAME4315(G4315,G6353,G6354);
  nand GNAME4316(G4316,G6319,G6320);
  nand GNAME4317(G4317,G6321,G6322);
  nand GNAME4318(G4318,G6323,G6324);
  nand GNAME4319(G4319,G6325,G6326);
  nand GNAME4320(G4320,G6327,G6328);
  nand GNAME4321(G4321,G6329,G6330);
  nand GNAME4322(G4322,G6331,G6332);
  nand GNAME4323(G4323,G6333,G6334);
  nand GNAME4324(G4324,G6355,G6356);
  nand GNAME4325(G4325,G6357,G6358);
  nand GNAME4326(G4326,G6269,G4680);
  nand GNAME4327(G4327,G6270,G4680);
  nand GNAME4328(G4328,G6273,G4680);
  nand GNAME4329(G4329,G6274,G6275);
  nand GNAME4330(G4330,G6276,G6277);
  nand GNAME4331(G4331,G6278,G6279);
  nand GNAME4332(G4332,G6280,G6281);
  nand GNAME4333(G4333,G6282,G6283);
  nand GNAME4334(G4334,G6284,G6285);
  nand GNAME4335(G4335,G6286,G6287);
  nand GNAME4336(G4336,G6288,G6289);
  nand GNAME4337(G4337,G6290,G6291);
  nand GNAME4338(G4338,G6294,G6295);
  nand GNAME4339(G4339,G6296,G6297);
  nand GNAME4340(G4340,G6298,G6299);
  nand GNAME4341(G4341,G6300,G6301);
  nand GNAME4342(G4342,G6302,G6303);
  nand GNAME4343(G4343,G6304,G6305);
  nand GNAME4344(G4344,G6306,G6307);
  nand GNAME4345(G4345,G6308,G6309);
  nand GNAME4346(G4346,G6310,G6311);
  nand GNAME4347(G4347,G6312,G6313);
  nand GNAME4348(G4348,G6254,G6255);
  nand GNAME4349(G4349,G6256,G6257);
  nand GNAME4350(G4350,G6258,G6259);
  nand GNAME4351(G4351,G6260,G6261);
  nand GNAME4352(G4352,G6262,G6263);
  nand GNAME4353(G4353,G6264,G6265);
  nand GNAME4354(G4354,G6271,G6272);
  nand GNAME4355(G4355,G6292,G6293);
  nand GNAME4356(G4356,G6314,G6315);
  nand GNAME4357(G4357,G6316,G6317);
  nand GNAME4358(G4358,G6250,G6251);
  and GNAME4359(G4359,G6252,G4567);
  and GNAME4360(G4360,G6252,G4566);
  and GNAME4361(G4361,G6252,G4565);
  and GNAME4362(G4362,G6252,G4564);
  and GNAME4363(G4363,G6252,G4563);
  and GNAME4364(G4364,G6252,G4562);
  and GNAME4365(G4365,G6252,G4561);
  and GNAME4366(G4366,G6252,G4560);
  and GNAME4367(G4367,G6252,G4559);
  and GNAME4368(G4368,G6249,G4759);
  and GNAME4369(G4369,G6249,G4757);
  and GNAME4370(G4370,G6249,G4754);
  and GNAME4371(G4371,G6249,G4751);
  and GNAME4372(G4372,G6249,G4748);
  and GNAME4373(G4373,G6249,G4745);
  and GNAME4374(G4374,G6249,G4742);
  and GNAME4375(G4375,G6249,G4739);
  and GNAME4376(G4376,G6249,G4736);
  and GNAME4377(G4377,G6249,G4733);
  and GNAME4378(G4378,G6249,G4730);
  and GNAME4379(G4379,G6249,G4727);
  and GNAME4380(G4380,G6249,G4724);
  and GNAME4381(G4381,G6249,G4721);
  and GNAME4382(G4382,G6249,G4718);
  and GNAME4383(G4383,G6249,G4715);
  and GNAME4384(G4384,G6249,G4712);
  and GNAME4385(G4385,G6249,G4709);
  and GNAME4386(G4386,G6249,G4706);
  and GNAME4387(G4387,G6249,G4701);
  nand GNAME4388(G4388,G36460,G5631);
  not GNAME4389(G4389,G36460);
  nand GNAME4390(G4390,G4987,G4985,G4986);
  nand GNAME4391(G4391,G4990,G4988,G4989);
  nand GNAME4392(G4392,G4993,G4991,G4992);
  nand GNAME4393(G4393,G4996,G4994,G4995);
  nand GNAME4394(G4394,G4999,G4997,G4998);
  nand GNAME4395(G4395,G5002,G5000,G5001);
  nand GNAME4396(G4396,G5005,G5003,G5004);
  nand GNAME4397(G4397,G5008,G5006,G5007);
  nand GNAME4398(G4398,G5011,G5009,G5010);
  nand GNAME4399(G4399,G5014,G5012,G5013);
  nand GNAME4400(G4400,G5017,G5015,G5016);
  nand GNAME4401(G4401,G5020,G5018,G5019);
  nand GNAME4402(G4402,G5023,G5021,G5022);
  nand GNAME4403(G4403,G5026,G5024,G5025);
  nand GNAME4404(G4404,G5029,G5027,G5028);
  nand GNAME4405(G4405,G5032,G5030,G5031);
  nand GNAME4406(G4406,G5035,G5033,G5034);
  nand GNAME4407(G4407,G5038,G5036,G5037);
  nand GNAME4408(G4408,G5041,G5039,G5040);
  nand GNAME4409(G4409,G5044,G5042,G5043);
  nand GNAME4410(G4410,G5047,G5045,G5046);
  nand GNAME4411(G4411,G5050,G5048,G5049);
  nand GNAME4412(G4412,G5053,G5051,G5052);
  nand GNAME4413(G4413,G5056,G5054,G5055);
  nand GNAME4414(G4414,G5059,G5057,G5058);
  nand GNAME4415(G4415,G5062,G5060,G5061);
  nand GNAME4416(G4416,G5065,G5063,G5064);
  nand GNAME4417(G4417,G5068,G5066,G5067);
  nand GNAME4418(G4418,G5071,G5069,G5070);
  nand GNAME4419(G4419,G5074,G5072,G5073);
  nand GNAME4420(G4420,G5077,G5075,G5076);
  nand GNAME4421(G4421,G5080,G5078,G5079);
  and GNAME4422(G4422,G4933,G36252);
  and GNAME4423(G4423,G4933,G36253);
  and GNAME4424(G4424,G4933,G36254);
  and GNAME4425(G4425,G4933,G36255);
  and GNAME4426(G4426,G4933,G36256);
  and GNAME4427(G4427,G4933,G36257);
  and GNAME4428(G4428,G4933,G36258);
  and GNAME4429(G4429,G4933,G36259);
  and GNAME4430(G4430,G4933,G36260);
  and GNAME4431(G4431,G4933,G36261);
  and GNAME4432(G4432,G4933,G36262);
  and GNAME4433(G4433,G4933,G36263);
  and GNAME4434(G4434,G4933,G36264);
  and GNAME4435(G4435,G4933,G36265);
  and GNAME4436(G4436,G4933,G36266);
  and GNAME4437(G4437,G4933,G36267);
  and GNAME4438(G4438,G4933,G36268);
  and GNAME4439(G4439,G4933,G36269);
  and GNAME4440(G4440,G4933,G36270);
  and GNAME4441(G4441,G4933,G36271);
  and GNAME4442(G4442,G4933,G36272);
  and GNAME4443(G4443,G4933,G36273);
  and GNAME4444(G4444,G4933,G36274);
  and GNAME4445(G4445,G4933,G36275);
  and GNAME4446(G4446,G4933,G36276);
  and GNAME4447(G4447,G4933,G36277);
  and GNAME4448(G4448,G4933,G36278);
  and GNAME4449(G4449,G4933,G36279);
  and GNAME4450(G4450,G4933,G36280);
  and GNAME4451(G4451,G4933,G36281);
  nand GNAME4452(G4452,G4845,G5417,G5415,G5416);
  nand GNAME4453(G4453,G4846,G5421,G5419,G5420);
  nand GNAME4454(G4454,G4847,G5430,G5428,G5429);
  nand GNAME4455(G4455,G4848,G5437,G5435,G5436);
  nand GNAME4456(G4456,G4849,G5444,G5442,G5443);
  nand GNAME4457(G4457,G4850,G5451,G5449,G5450);
  nand GNAME4458(G4458,G4851,G5458,G5456,G5457);
  nand GNAME4459(G4459,G4852,G5465,G5463,G5464);
  nand GNAME4460(G4460,G4853,G5472,G5470,G5471);
  nand GNAME4461(G4461,G4854,G5479,G5477,G5478);
  nand GNAME4462(G4462,G4855,G5486,G5484,G5485);
  nand GNAME4463(G4463,G4856,G5493,G5491,G5492);
  nand GNAME4464(G4464,G4857,G5500,G5498,G5499);
  nand GNAME4465(G4465,G4858,G5507,G5505,G5506);
  nand GNAME4466(G4466,G4859,G5514,G5512,G5513);
  nand GNAME4467(G4467,G4860,G5521,G5519,G5520);
  nand GNAME4468(G4468,G4861,G5528,G5526,G5527);
  nand GNAME4469(G4469,G4862,G5535,G5533,G5534);
  nand GNAME4470(G4470,G4863,G5542,G5540,G5541);
  nand GNAME4471(G4471,G4864,G5549,G5547,G5548);
  nand GNAME4472(G4472,G4865,G5556,G5554,G5555);
  nand GNAME4473(G4473,G4866,G5563,G5561,G5562);
  nand GNAME4474(G4474,G4867,G5570,G5568,G5569);
  nand GNAME4475(G4475,G4868,G5577,G5575,G5576);
  nand GNAME4476(G4476,G4869,G5584,G5582,G5583);
  nand GNAME4477(G4477,G4870,G5591,G5589,G5590);
  nand GNAME4478(G4478,G4871,G5598,G5596,G5597);
  nand GNAME4479(G4479,G4872,G5605,G5603,G5604);
  nand GNAME4480(G4480,G4873,G5612,G5610,G5611);
  nand GNAME4481(G4481,G5616,G4937,G5615,G5613,G5614);
  nand GNAME4482(G4482,G5619,G6953,G6954);
  nand GNAME4483(G4483,G5622,G6955,G6956);
  nand GNAME4484(G4484,G4874,G5637,G5635,G5636);
  nand GNAME4485(G4485,G4875,G5646,G5644,G5645);
  nand GNAME4486(G4486,G4876,G5655,G5653,G5654);
  nand GNAME4487(G4487,G4877,G5664,G5662,G5663);
  nand GNAME4488(G4488,G4878,G5673,G5671,G5672);
  nand GNAME4489(G4489,G4879,G5682,G5680,G5681);
  nand GNAME4490(G4490,G4880,G5691,G5689,G5690);
  nand GNAME4491(G4491,G4881,G5700,G5698,G5699);
  nand GNAME4492(G4492,G4882,G5709,G5707,G5708);
  nand GNAME4493(G4493,G4883,G5718,G5716,G5717);
  nand GNAME4494(G4494,G4884,G5727,G5725,G5726);
  nand GNAME4495(G4495,G4885,G5736,G5734,G5735);
  nand GNAME4496(G4496,G4886,G5745,G5743,G5744);
  nand GNAME4497(G4497,G4887,G5754,G5752,G5753);
  nand GNAME4498(G4498,G4888,G5763,G5761,G5762);
  nand GNAME4499(G4499,G4889,G5772,G5770,G5771);
  nand GNAME4500(G4500,G4890,G5781,G5779,G5780);
  nand GNAME4501(G4501,G4891,G5790,G5788,G5789);
  nand GNAME4502(G4502,G4892,G5799,G5800,G5798);
  nand GNAME4503(G4503,G4893,G5808,G5809,G5807);
  nand GNAME4504(G4504,G5825,G5823,G5824);
  nand GNAME4505(G4505,G4901,G5838,G5836,G5839);
  nand GNAME4506(G4506,G4902,G5853,G5851,G5852);
  nand GNAME4507(G4507,G4903,G5860,G5861,G5859);
  nand GNAME4508(G4508,G4904,G5870,G5868,G5871);
  nand GNAME4509(G4509,G4905,G5880,G5878,G5879);
  nand GNAME4510(G4510,G4906,G5890,G5891,G5889);
  nand GNAME4511(G4511,G4907,G5903,G5901,G5902);
  nand GNAME4512(G4512,G4908,G5910,G5911,G5909);
  nand GNAME4513(G4513,G4909,G5923,G5921,G5922);
  nand GNAME4514(G4514,G4910,G5929,G5927,G5928);
  nand GNAME4515(G4515,G4911,G5939,G5940,G5938);
  nand GNAME4516(G4516,G4912,G5949,G5950,G5948);
  nand GNAME4517(G4517,G4913,G5962,G5960,G5961);
  nand GNAME4518(G4518,G4914,G5969,G5967,G5970);
  nand GNAME4519(G4519,G4915,G5979,G5980,G5978);
  nand GNAME4520(G4520,G4916,G5989,G5987,G5990);
  nand GNAME4521(G4521,G4917,G6002,G6000,G6001);
  nand GNAME4522(G4522,G4918,G6009,G6010,G6008);
  nand GNAME4523(G4523,G4919,G6022,G6020,G6021);
  nand GNAME4524(G4524,G4920,G6029,G6027,G6028);
  nand GNAME4525(G4525,G4921,G6039,G6040,G6038);
  nand GNAME4526(G4526,G4922,G6052,G6050,G6051);
  nand GNAME4527(G4527,G4923,G6059,G6057,G6060);
  nand GNAME4528(G4528,G4924,G6069,G6067,G6068);
  nand GNAME4529(G4529,G4925,G6079,G6080,G6078);
  nand GNAME4530(G4530,G4926,G6092,G6090,G6091);
  nand GNAME4531(G4531,G4927,G6099,G6100,G6098);
  nand GNAME4532(G4532,G4928,G6112,G6110,G6111);
  nand GNAME4533(G4533,G4929,G6119,G6120,G6118);
  nor GNAME4534(G4534,G4389,G4535);
  and GNAME4535(G4535,G36460,G4932);
  not GNAME4536(G4536,G13813);
  not GNAME4537(G4537,G36247);
  not GNAME4538(G4538,G36248);
  nand GNAME4539(G4539,G6693,G4690);
  nor GNAME4540(G4540,G4691,G5082);
  nand GNAME4541(G4541,G4689,G6693);
  not GNAME4542(G4542,G36430);
  and GNAME4543(G4543,G36460,G4540);
  nand GNAME4544(G4544,G6693,G6696,G6697);
  and GNAME4545(G4545,G4940,G5087);
  and GNAME4546(G4546,G6743,G6746);
  and GNAME4547(G4547,G4695,G4696);
  nor GNAME4548(G4548,G4694,G4970);
  nor GNAME4549(G4549,G4697,G6731);
  nand GNAME4550(G4550,G6725,G4549);
  nand GNAME4551(G4551,G6725,G4697);
  and GNAME4552(G4552,G6728,G6731);
  and GNAME4553(G4553,G4695,G4552);
  and GNAME4554(G4554,G6731,G6722);
  nand GNAME4555(G4555,G6728,G4696);
  or GNAME4556(G4556,G4695,G4555);
  or GNAME4557(G4557,G4586,G4961,G4584);
  nor GNAME4558(G4558,G6719,G4970);
  and GNAME4559(G4559,G4959,G845);
  and GNAME4560(G4560,G4959,G844);
  and GNAME4561(G4561,G4959,G843);
  and GNAME4562(G4562,G4959,G842);
  and GNAME4563(G4563,G4959,G841);
  and GNAME4564(G4564,G4959,G840);
  and GNAME4565(G4565,G4959,G839);
  and GNAME4566(G4566,G4959,G838);
  and GNAME4567(G4567,G4959,G837);
  and GNAME4568(G4568,G4959,G836);
  and GNAME4569(G4569,G6725,G4554);
  and GNAME4570(G4570,G4959,G834);
  and GNAME4571(G4571,G4959,G833);
  and GNAME4572(G4572,G4702,G6746);
  and GNAME4573(G4573,G4703,G6743);
  or GNAME4574(G4574,G4695,G4551);
  nand GNAME4575(G4575,G5407,G4543);
  and GNAME4576(G4576,G4548,G4969);
  and GNAME4577(G4577,G5411,G4969);
  nand GNAME4578(G4578,G6722,G6725,G6728);
  and GNAME4579(G4579,G5409,G4969);
  or GNAME4580(G4580,G4698,G4574);
  nor GNAME4581(G4581,G4575,G4580);
  nor GNAME4582(G4582,G5408,G4575);
  and GNAME4583(G4583,G4558,G4969);
  and GNAME4584(G4584,G4697,G4696);
  and GNAME4585(G4585,G4697,G6731);
  and GNAME4586(G4586,G4698,G4695);
  nand GNAME4587(G4587,G4958,G4664,G4957,G4948,G4649);
  nor GNAME4588(G4588,G4698,G4578);
  or GNAME4589(G4589,G4689,G4539);
  and GNAME4590(G4590,G6700,G5082);
  and GNAME4591(G4591,G36460,G4590);
  nor GNAME4592(G4592,G6719,G4965);
  and GNAME4593(G4593,G36460,G4691);
  or GNAME4594(G4594,G4642,G4639);
  and GNAME4595(G4595,G4597,G5624);
  and GNAME4596(G4596,G4598,G5624);
  or GNAME4597(G4597,G4960,G4594,G4588,G4949,G4553);
  or GNAME4598(G4598,G4668,G4587);
  and GNAME4599(G4599,G5623,G6719);
  and GNAME4600(G4600,G4603,G4543);
  and GNAME4601(G4601,G4694,G4700);
  and GNAME4602(G4602,G5634,G36460,G4603);
  or GNAME4603(G4603,G4388,G4590);
  and GNAME4604(G4604,G4696,G4553);
  and GNAME4605(G4605,G4601,G4604);
  nand GNAME4606(G4606,G5114,G5115,G5116,G5117);
  nand GNAME4607(G4607,G5164,G5165,G5166,G5167);
  nand GNAME4608(G4608,G5088,G5089,G5090,G5091);
  nand GNAME4609(G4609,G5124,G5125,G5126,G5127);
  nand GNAME4610(G4610,G5100,G5101,G5102,G5103);
  nand GNAME4611(G4611,G5144,G5145,G5146,G5147);
  nand GNAME4612(G4612,G5154,G5155,G5156,G5157);
  nand GNAME4613(G4613,G5134,G5135,G5136,G5137);
  nand GNAME4614(G4614,G5184,G5185,G5186,G5187);
  nand GNAME4615(G4615,G5174,G5175,G5176,G5177);
  nand GNAME4616(G4616,G5324,G5325,G5326,G5327);
  nand GNAME4617(G4617,G5294,G5295,G5296,G5297);
  nand GNAME4618(G4618,G5374,G5375,G5376,G5377);
  nand GNAME4619(G4619,G5334,G5335,G5336,G5337);
  nand GNAME4620(G4620,G5314,G5315,G5316,G5317);
  nand GNAME4621(G4621,G5284,G5285,G5286,G5287);
  nand GNAME4622(G4622,G5304,G5305,G5306,G5307);
  nand GNAME4623(G4623,G5354,G5355,G5356,G5357);
  nand GNAME4624(G4624,G5364,G5365,G5366,G5367);
  nand GNAME4625(G4625,G5234,G5235,G5236,G5237);
  nand GNAME4626(G4626,G5344,G5345,G5346,G5347);
  nand GNAME4627(G4627,G5194,G5195,G5196,G5197);
  nand GNAME4628(G4628,G5224,G5225,G5226,G5227);
  nand GNAME4629(G4629,G5214,G5215,G5216,G5217);
  nand GNAME4630(G4630,G5244,G5245,G5246,G5247);
  nand GNAME4631(G4631,G5204,G5205,G5206,G5207);
  nand GNAME4632(G4632,G5254,G5255,G5256,G5257);
  nand GNAME4633(G4633,G5274,G5275,G5276,G5277);
  nand GNAME4634(G4634,G5264,G5265,G5266,G5267);
  and GNAME4635(G4635,G4897,G4898,G4896,G4894,G4895);
  and GNAME4636(G4636,G4899,G4900);
  nand GNAME4637(G4637,G5104,G5105,G5106,G5107);
  and GNAME4638(G4638,G4635,G4636);
  nor GNAME4639(G4639,G4695,G4550);
  nand GNAME4640(G4640,G4696,G4549);
  and GNAME4641(G4641,G6722,G4949);
  nor GNAME4642(G4642,G6731,G4574);
  nand GNAME4643(G4643,G6722,G4584);
  nor GNAME4644(G4644,G6731,G4643);
  nor GNAME4645(G4645,G6722,G4698);
  nor GNAME4646(G4646,G6746,G6743);
  and GNAME4647(G4647,G4594,G4543);
  nand GNAME4648(G4648,G4545,G4646);
  nand GNAME4649(G4649,G4695,G4585);
  or GNAME4650(G4650,G4641,G4950,G4588);
  nand GNAME4651(G4651,G4951,G7121,G4643,G5831);
  nor GNAME4652(G4652,G5835,G4591,G4593);
  and GNAME4653(G4653,G4543,G4964);
  and GNAME4654(G4654,G4650,G4653);
  and GNAME4655(G4655,G4651,G4653);
  nor GNAME4656(G4656,G6719,G4648);
  nor GNAME4657(G4657,G4694,G4648);
  nor GNAME4658(G4658,G5082,G4240,G4389);
  and GNAME4659(G4659,G5847,G4543);
  and GNAME4660(G4660,G4589,G4644);
  and GNAME4661(G4661,G4540,G4586);
  and GNAME4662(G4662,G4697,G4661);
  and GNAME4663(G4663,G6728,G4661);
  nand GNAME4664(G4664,G4696,G4585);
  nor GNAME4665(G4665,G5082,G4664);
  nand GNAME4666(G4666,G4941,G4943,G4945,G4946);
  nand GNAME4667(G4667,G4977,G4978,G4979,G4980);
  and GNAME4668(G4668,G4696,G4552);
  and GNAME4669(G4669,G4589,G4668);
  nand GNAME4670(G4670,G4589,G4585);
  nand GNAME4671(G4671,G4695,G4646);
  nand GNAME4672(G4672,G6700,G6736);
  nor GNAME4673(G4673,G4589,G4672);
  and GNAME4674(G4674,G5082,G4700,G6700);
  and GNAME4675(G4675,G4956,G4953,G4955);
  nand GNAME4676(G4676,G4671,G4954);
  nand GNAME4677(G4677,G4981,G4675);
  and GNAME4678(G4678,G4554,G4646);
  and GNAME4679(G4679,G6684,G4554);
  and GNAME4680(G4680,G6268,G6266,G6267);
  and GNAME4681(G4681,G4931,G4574,G7122,G4578);
  nand GNAME4682(G4682,G4947,G4550,G4948,G4640);
  and GNAME4683(G4683,G4682,G13899);
  or GNAME4684(G4684,G4666,G4667);
  and GNAME4685(G4685,G6685,G4589,G6736);
  and GNAME4686(G4686,G4700,G4589,G6685);
  and GNAME4687(G4687,G6586,G6587);
  and GNAME4688(G4688,G6591,G4687,G6590,G6588,G6589);
  and GNAME4689(G4689,G6689,G6690);
  nand GNAME4690(G4690,G6694,G6695);
  nand GNAME4691(G4691,G6698,G6699);
  nand GNAME4692(G4692,G6701,G6702);
  nand GNAME4693(G4693,G6703,G6704);
  nand GNAME4694(G4694,G6717,G6718);
  nand GNAME4695(G4695,G6720,G6721);
  nand GNAME4696(G4696,G6723,G6724);
  nand GNAME4697(G4697,G6726,G6727);
  nand GNAME4698(G4698,G6729,G6730);
  nand GNAME4699(G4699,G6732,G6733);
  nand GNAME4700(G4700,G6734,G6735);
  nand GNAME4701(G4701,G6737,G6738);
  nand GNAME4702(G4702,G6741,G6742);
  nand GNAME4703(G4703,G6744,G6745);
  nand GNAME4704(G4704,G6747,G6748);
  nand GNAME4705(G4705,G6749,G6750);
  nand GNAME4706(G4706,G6751,G6752);
  nand GNAME4707(G4707,G6753,G6754);
  nand GNAME4708(G4708,G6755,G6756);
  nand GNAME4709(G4709,G6757,G6758);
  nand GNAME4710(G4710,G6759,G6760);
  nand GNAME4711(G4711,G6761,G6762);
  nand GNAME4712(G4712,G6763,G6764);
  nand GNAME4713(G4713,G6765,G6766);
  nand GNAME4714(G4714,G6767,G6768);
  nand GNAME4715(G4715,G6769,G6770);
  nand GNAME4716(G4716,G6771,G6772);
  nand GNAME4717(G4717,G6773,G6774);
  nand GNAME4718(G4718,G6775,G6776);
  nand GNAME4719(G4719,G6777,G6778);
  nand GNAME4720(G4720,G6779,G6780);
  nand GNAME4721(G4721,G6781,G6782);
  nand GNAME4722(G4722,G6783,G6784);
  nand GNAME4723(G4723,G6785,G6786);
  nand GNAME4724(G4724,G6787,G6788);
  nand GNAME4725(G4725,G6789,G6790);
  nand GNAME4726(G4726,G6791,G6792);
  nand GNAME4727(G4727,G6793,G6794);
  nand GNAME4728(G4728,G6795,G6796);
  nand GNAME4729(G4729,G6797,G6798);
  nand GNAME4730(G4730,G6799,G6800);
  nand GNAME4731(G4731,G6801,G6802);
  nand GNAME4732(G4732,G6803,G6804);
  nand GNAME4733(G4733,G6805,G6806);
  nand GNAME4734(G4734,G6807,G6808);
  nand GNAME4735(G4735,G6809,G6810);
  nand GNAME4736(G4736,G6811,G6812);
  nand GNAME4737(G4737,G6813,G6814);
  nand GNAME4738(G4738,G6815,G6816);
  nand GNAME4739(G4739,G6817,G6818);
  nand GNAME4740(G4740,G6819,G6820);
  nand GNAME4741(G4741,G6821,G6822);
  nand GNAME4742(G4742,G6823,G6824);
  nand GNAME4743(G4743,G6825,G6826);
  nand GNAME4744(G4744,G6827,G6828);
  nand GNAME4745(G4745,G6829,G6830);
  nand GNAME4746(G4746,G6831,G6832);
  nand GNAME4747(G4747,G6833,G6834);
  nand GNAME4748(G4748,G6835,G6836);
  nand GNAME4749(G4749,G6837,G6838);
  nand GNAME4750(G4750,G6839,G6840);
  nand GNAME4751(G4751,G6841,G6842);
  nand GNAME4752(G4752,G6843,G6844);
  nand GNAME4753(G4753,G6845,G6846);
  nand GNAME4754(G4754,G6847,G6848);
  nand GNAME4755(G4755,G6849,G6850);
  nand GNAME4756(G4756,G6851,G6852);
  nand GNAME4757(G4757,G6853,G6854);
  nand GNAME4758(G4758,G6855,G6856);
  nand GNAME4759(G4759,G6857,G6858);
  nand GNAME4760(G4760,G6859,G6860);
  nand GNAME4761(G4761,G6861,G6862);
  nand GNAME4762(G4762,G6863,G6864);
  nand GNAME4763(G4763,G6865,G6866);
  nand GNAME4764(G4764,G6867,G6868);
  nand GNAME4765(G4765,G6869,G6870);
  nand GNAME4766(G4766,G6871,G6872);
  nand GNAME4767(G4767,G6873,G6874);
  nand GNAME4768(G4768,G6875,G6876);
  nand GNAME4769(G4769,G6877,G6878);
  nand GNAME4770(G4770,G6879,G6880);
  nand GNAME4771(G4771,G6881,G6882);
  nand GNAME4772(G4772,G6883,G6884);
  nand GNAME4773(G4773,G6885,G6886);
  nand GNAME4774(G4774,G6887,G6888);
  nand GNAME4775(G4775,G6889,G6890);
  nand GNAME4776(G4776,G6891,G6892);
  nand GNAME4777(G4777,G6893,G6894);
  nand GNAME4778(G4778,G6895,G6896);
  nand GNAME4779(G4779,G6897,G6898);
  nand GNAME4780(G4780,G6899,G6900);
  nand GNAME4781(G4781,G6901,G6902);
  nand GNAME4782(G4782,G6903,G6904);
  nand GNAME4783(G4783,G6905,G6906);
  nand GNAME4784(G4784,G6907,G6908);
  nand GNAME4785(G4785,G6909,G6910);
  nand GNAME4786(G4786,G6911,G6912);
  nand GNAME4787(G4787,G6913,G6914);
  nand GNAME4788(G4788,G6915,G6916);
  nand GNAME4789(G4789,G6917,G6918);
  nand GNAME4790(G4790,G6919,G6920);
  nand GNAME4791(G4791,G6921,G6922);
  nand GNAME4792(G4792,G6923,G6924);
  nand GNAME4793(G4793,G6925,G6926);
  nand GNAME4794(G4794,G6927,G6928);
  nand GNAME4795(G4795,G6929,G6930);
  nand GNAME4796(G4796,G6931,G6932);
  nand GNAME4797(G4797,G6933,G6934);
  nand GNAME4798(G4798,G6935,G6936);
  nand GNAME4799(G4799,G6937,G6938);
  nand GNAME4800(G4800,G6939,G6940);
  nand GNAME4801(G4801,G6941,G6942);
  nand GNAME4802(G4802,G6943,G6944);
  nand GNAME4803(G4803,G6945,G6946);
  nand GNAME4804(G4804,G6947,G6948);
  nand GNAME4805(G4805,G6957,G6958);
  nand GNAME4806(G4806,G6959,G6960);
  nand GNAME4807(G4807,G6961,G6962);
  nand GNAME4808(G4808,G6963,G6964);
  nand GNAME4809(G4809,G6965,G6966);
  nand GNAME4810(G4810,G6967,G6968);
  nand GNAME4811(G4811,G6969,G6970);
  nand GNAME4812(G4812,G6971,G6972);
  nand GNAME4813(G4813,G6973,G6974);
  nand GNAME4814(G4814,G6975,G6976);
  nand GNAME4815(G4815,G6977,G6978);
  nand GNAME4816(G4816,G6979,G6980);
  nand GNAME4817(G4817,G6981,G6982);
  nand GNAME4818(G4818,G6983,G6984);
  nand GNAME4819(G4819,G6985,G6986);
  nand GNAME4820(G4820,G6987,G6988);
  nand GNAME4821(G4821,G6989,G6990);
  nand GNAME4822(G4822,G6991,G6992);
  nand GNAME4823(G4823,G6993,G6994);
  nand GNAME4824(G4824,G6995,G6996);
  nand GNAME4825(G4825,G6997,G6998);
  nand GNAME4826(G4826,G6999,G7000);
  nand GNAME4827(G4827,G7001,G7002);
  nand GNAME4828(G4828,G7003,G7004);
  nand GNAME4829(G4829,G7005,G7006);
  nand GNAME4830(G4830,G7007,G7008);
  nand GNAME4831(G4831,G7009,G7010);
  nand GNAME4832(G4832,G7011,G7012);
  nand GNAME4833(G4833,G7013,G7014);
  nand GNAME4834(G4834,G7015,G7016);
  nand GNAME4835(G4835,G7017,G7018);
  nand GNAME4836(G4836,G7019,G7020);
  or GNAME4837(G4837,G36278,G36279,G36280,G36281);
  nor GNAME4838(G4838,G4837,G36277,G36276,G36275,G36274);
  or GNAME4839(G4839,G36270,G36271,G36272,G36273);
  nor GNAME4840(G4840,G4839,G36267,G36269,G36268);
  or GNAME4841(G4841,G36263,G36264,G36265,G36266);
  nor GNAME4842(G4842,G4841,G36260,G36262,G36261);
  or GNAME4843(G4843,G36256,G36257,G36258,G36259);
  nor GNAME4844(G4844,G4843,G36253,G36255,G36254);
  and GNAME4845(G4845,G5414,G5412,G5413);
  and GNAME4846(G4846,G6949,G6950,G5422,G5423);
  and GNAME4847(G4847,G5424,G5425,G5426,G5427);
  and GNAME4848(G4848,G5431,G5432,G5433,G5434);
  and GNAME4849(G4849,G5438,G5439,G5440,G5441);
  and GNAME4850(G4850,G5445,G5446,G5447,G5448);
  and GNAME4851(G4851,G5452,G5453,G5454,G5455);
  and GNAME4852(G4852,G5459,G5460,G5461,G5462);
  and GNAME4853(G4853,G5466,G5467,G5468,G5469);
  and GNAME4854(G4854,G5473,G5474,G5475,G5476);
  and GNAME4855(G4855,G5480,G5481,G5482,G5483);
  and GNAME4856(G4856,G5487,G5488,G5489,G5490);
  and GNAME4857(G4857,G5494,G5495,G5496,G5497);
  and GNAME4858(G4858,G5501,G5502,G5503,G5504);
  and GNAME4859(G4859,G5508,G5509,G5510,G5511);
  and GNAME4860(G4860,G5515,G5516,G5517,G5518);
  and GNAME4861(G4861,G5522,G5523,G5524,G5525);
  and GNAME4862(G4862,G5529,G5530,G5531,G5532);
  and GNAME4863(G4863,G5536,G5537,G5538,G5539);
  and GNAME4864(G4864,G5543,G5544,G5545,G5546);
  and GNAME4865(G4865,G5550,G5551,G5552,G5553);
  and GNAME4866(G4866,G5557,G5558,G5559,G5560);
  and GNAME4867(G4867,G5564,G5565,G5566,G5567);
  and GNAME4868(G4868,G5571,G5572,G5573,G5574);
  and GNAME4869(G4869,G5578,G5579,G5580,G5581);
  and GNAME4870(G4870,G5585,G5586,G5587,G5588);
  and GNAME4871(G4871,G5592,G5593,G5594,G5595);
  and GNAME4872(G4872,G5599,G5600,G5601,G5602);
  and GNAME4873(G4873,G5606,G5607,G5608,G5609);
  and GNAME4874(G4874,G5639,G6062,G5638);
  and GNAME4875(G4875,G5648,G5873,G5647);
  and GNAME4876(G4876,G5657,G5972,G5656);
  and GNAME4877(G4877,G5666,G5992,G5665);
  and GNAME4878(G4878,G5675,G5841,G5674);
  and GNAME4879(G4879,G5684,G6102,G5683);
  and GNAME4880(G4880,G5693,G5913,G5692);
  and GNAME4881(G4881,G5702,G6012,G5701);
  and GNAME4882(G4882,G5711,G5893,G5710);
  and GNAME4883(G4883,G5720,G6082,G5719);
  and GNAME4884(G4884,G5729,G5942,G5728);
  and GNAME4885(G4885,G5738,G6042,G5737);
  and GNAME4886(G4886,G5747,G6122,G5746);
  and GNAME4887(G4887,G5756,G5863,G5755);
  and GNAME4888(G4888,G5765,G5982,G5764);
  and GNAME4889(G4889,G5774,G5952,G5773);
  and GNAME4890(G4890,G5783,G6072,G5782);
  and GNAME4891(G4891,G5792,G5883,G5791);
  and GNAME4892(G4892,G5801,G6032,G5797);
  and GNAME4893(G4893,G5810,G5932,G5806);
  and GNAME4894(G4894,G7055,G7058,G7061);
  and GNAME4895(G4895,G7064,G7067,G7070);
  and GNAME4896(G4896,G7082,G7085,G7073,G7076,G7079);
  and GNAME4897(G4897,G7097,G7100,G7088,G7091,G7094);
  and GNAME4898(G4898,G7112,G7115,G7103,G7106,G7109);
  and GNAME4899(G4899,G7034,G7037,G7025,G7028,G7031);
  and GNAME4900(G4900,G7049,G7052,G7040,G7043,G7046);
  and GNAME4901(G4901,G5841,G5837,G5840);
  and GNAME4902(G4902,G5850,G5848,G5849);
  and GNAME4903(G4903,G5863,G5858,G5862);
  and GNAME4904(G4904,G5873,G5869,G5872);
  and GNAME4905(G4905,G5883,G5881,G5882);
  and GNAME4906(G4906,G5893,G5888,G5892);
  and GNAME4907(G4907,G5900,G5898,G5899);
  and GNAME4908(G4908,G5913,G5908,G5912);
  and GNAME4909(G4909,G5920,G5918,G5919);
  and GNAME4910(G4910,G5932,G5930,G5931);
  and GNAME4911(G4911,G5942,G5937,G5941);
  and GNAME4912(G4912,G5952,G5947,G5951);
  and GNAME4913(G4913,G5959,G5957,G5958);
  and GNAME4914(G4914,G5972,G5968,G5971);
  and GNAME4915(G4915,G5982,G5977,G5981);
  and GNAME4916(G4916,G5992,G5988,G5991);
  and GNAME4917(G4917,G5999,G5997,G5998);
  and GNAME4918(G4918,G6012,G6007,G6011);
  and GNAME4919(G4919,G6019,G6017,G6018);
  and GNAME4920(G4920,G6032,G6030,G6031);
  and GNAME4921(G4921,G6042,G6037,G6041);
  and GNAME4922(G4922,G6049,G6047,G6048);
  and GNAME4923(G4923,G6062,G6058,G6061);
  and GNAME4924(G4924,G6072,G6070,G6071);
  and GNAME4925(G4925,G6082,G6077,G6081);
  and GNAME4926(G4926,G6089,G6087,G6088);
  and GNAME4927(G4927,G6102,G6097,G6101);
  and GNAME4928(G4928,G6109,G6107,G6108);
  and GNAME4929(G4929,G6122,G6117,G6121);
  or GNAME4930(G4930,G4553,G4588);
  and GNAME4931(G4931,G4556,G6361,G4643);
  not GNAME4932(G4932,G36249);
  nand GNAME4933(G4933,G4544,G4543);
  and GNAME4934(G4934,G6719,G6736);
  nand GNAME4935(G4935,G5085,G4543,G4545,G4546);
  nand GNAME4936(G4936,G5085,G4543,G4545,G4572);
  and GNAME4937(G4937,G6951,G6952);
  not GNAME4938(G4938,G13005);
  and GNAME4939(G4939,G7119,G5818);
  nand GNAME4940(G4940,G5086,G5081);
  nand GNAME4941(G4941,G4646,G4665);
  nand GNAME4942(G4942,G4646,G4669);
  nand GNAME4943(G4943,G4646,G4662);
  or GNAME4944(G4944,G4670,G4671);
  nand GNAME4945(G4945,G4646,G4660);
  nand GNAME4946(G4946,G4646,G4663);
  or GNAME4947(G4947,G6731,G4551);
  nand GNAME4948(G4948,G4698,G4584);
  not GNAME4949(G4949,G4640);
  and GNAME4950(G4950,G6725,G4553);
  or GNAME4951(G4951,G4696,G4649);
  nand GNAME4952(G4952,G6736,G4691);
  nand GNAME4953(G4953,G4695,G4573);
  nand GNAME4954(G4954,G4698,G4646);
  nand GNAME4955(G4955,G4695,G4572);
  nand GNAME4956(G4956,G4695,G4546);
  nand GNAME4957(G4957,G4695,G4549);
  nand GNAME4958(G4958,G4697,G4586);
  not GNAME4959(G4959,G4934);
  not GNAME4960(G4960,G4580);
  nor GNAME4961(G4961,G4698,G4556);
  nand GNAME4962(G4962,G4982,G4547);
  nand GNAME4963(G4963,G4636,G4635,G7118);
  not GNAME4964(G4964,G4648);
  not GNAME4965(G4965,G4591);
  not GNAME4966(G4966,G4933);
  not GNAME4967(G4967,G4935);
  not GNAME4968(G4968,G4936);
  not GNAME4969(G4969,G4575);
  not GNAME4970(G4970,G4547);
  nand GNAME4971(G4971,G4547,G5388,G4207);
  nand GNAME4972(G4972,G4593,G4603,G6719);
  nand GNAME4973(G4973,G4543,G4960);
  nand GNAME4974(G4974,G6123,G4697);
  or GNAME4975(G4975,G4675,G4670);
  nand GNAME4976(G4976,G6684,G4669);
  nand GNAME4977(G4977,G6684,G4660);
  nand GNAME4978(G4978,G6684,G4662);
  nand GNAME4979(G4979,G6684,G4663);
  nand GNAME4980(G4980,G6684,G4665);
  nand GNAME4981(G4981,G6684,G4698);
  not GNAME4982(G4982,G4552);
  not GNAME4983(G4983,G4590);
  nand GNAME4984(G4984,G4697,G4554);
  nand GNAME4985(G4985,G4389,G857);
  nand GNAME4986(G4986,G4534,G36218);
  nand GNAME4987(G4987,G4535,G36218);
  nand GNAME4988(G4988,G4389,G846);
  nand GNAME4989(G4989,G4534,G13833);
  nand GNAME4990(G4990,G4535,G36219);
  nand GNAME4991(G4991,G4389,G835);
  nand GNAME4992(G4992,G4534,G13814);
  nand GNAME4993(G4993,G4535,G36220);
  nand GNAME4994(G4994,G4389,G832);
  nand GNAME4995(G4995,G4534,G13815);
  nand GNAME4996(G4996,G4535,G36221);
  nand GNAME4997(G4997,G4389,G831);
  nand GNAME4998(G4998,G4534,G13838);
  nand GNAME4999(G4999,G4535,G36222);
  nand GNAME5000(G5000,G4389,G830);
  nand GNAME5001(G5001,G4534,G13837);
  nand GNAME5002(G5002,G4535,G36223);
  nand GNAME5003(G5003,G4389,G829);
  nand GNAME5004(G5004,G4534,G13816);
  nand GNAME5005(G5005,G4535,G36224);
  nand GNAME5006(G5006,G4389,G828);
  nand GNAME5007(G5007,G4534,G13817);
  nand GNAME5008(G5008,G4535,G36225);
  nand GNAME5009(G5009,G4389,G827);
  nand GNAME5010(G5010,G4534,G13836);
  nand GNAME5011(G5011,G4535,G36226);
  nand GNAME5012(G5012,G4389,G826);
  nand GNAME5013(G5013,G4534,G13835);
  nand GNAME5014(G5014,G4535,G36227);
  nand GNAME5015(G5015,G4389,G856);
  nand GNAME5016(G5016,G4534,G13803);
  nand GNAME5017(G5017,G4535,G36228);
  nand GNAME5018(G5018,G4389,G855);
  nand GNAME5019(G5019,G4534,G13804);
  nand GNAME5020(G5020,G4535,G36229);
  nand GNAME5021(G5021,G4389,G854);
  nand GNAME5022(G5022,G4534,G13850);
  nand GNAME5023(G5023,G4535,G36230);
  nand GNAME5024(G5024,G4389,G853);
  nand GNAME5025(G5025,G4534,G13849);
  nand GNAME5026(G5026,G4535,G36231);
  nand GNAME5027(G5027,G4389,G852);
  nand GNAME5028(G5028,G4534,G13805);
  nand GNAME5029(G5029,G4535,G36232);
  nand GNAME5030(G5030,G4389,G851);
  nand GNAME5031(G5031,G4534,G13806);
  nand GNAME5032(G5032,G4535,G36233);
  nand GNAME5033(G5033,G4389,G850);
  nand GNAME5034(G5034,G4534,G13848);
  nand GNAME5035(G5035,G4535,G36234);
  nand GNAME5036(G5036,G4389,G849);
  nand GNAME5037(G5037,G4534,G13847);
  nand GNAME5038(G5038,G4535,G36235);
  nand GNAME5039(G5039,G4389,G848);
  nand GNAME5040(G5040,G4534,G13807);
  nand GNAME5041(G5041,G4535,G36236);
  nand GNAME5042(G5042,G4389,G847);
  nand GNAME5043(G5043,G4534,G13808);
  nand GNAME5044(G5044,G4535,G36237);
  nand GNAME5045(G5045,G4389,G845);
  nand GNAME5046(G5046,G4534,G13845);
  nand GNAME5047(G5047,G4535,G36238);
  nand GNAME5048(G5048,G4389,G844);
  nand GNAME5049(G5049,G4534,G13844);
  nand GNAME5050(G5050,G4535,G36239);
  nand GNAME5051(G5051,G4389,G843);
  nand GNAME5052(G5052,G4534,G13809);
  nand GNAME5053(G5053,G4535,G36240);
  nand GNAME5054(G5054,G4389,G842);
  nand GNAME5055(G5055,G4534,G13810);
  nand GNAME5056(G5056,G4535,G36241);
  nand GNAME5057(G5057,G4389,G841);
  nand GNAME5058(G5058,G4534,G13843);
  nand GNAME5059(G5059,G4535,G36242);
  nand GNAME5060(G5060,G4389,G840);
  nand GNAME5061(G5061,G4534,G13842);
  nand GNAME5062(G5062,G4535,G36243);
  nand GNAME5063(G5063,G4389,G839);
  nand GNAME5064(G5064,G4534,G13811);
  nand GNAME5065(G5065,G4535,G36244);
  nand GNAME5066(G5066,G4389,G838);
  nand GNAME5067(G5067,G4534,G13812);
  nand GNAME5068(G5068,G4535,G36245);
  nand GNAME5069(G5069,G4389,G837);
  nand GNAME5070(G5070,G4534,G13841);
  nand GNAME5071(G5071,G4535,G36246);
  nand GNAME5072(G5072,G4389,G836);
  nand GNAME5073(G5073,G4534,G13813);
  nand GNAME5074(G5074,G4535,G36247);
  nand GNAME5075(G5075,G4389,G834);
  nand GNAME5076(G5076,G4534,G13840);
  nand GNAME5077(G5077,G4535,G36248);
  nand GNAME5078(G5078,G4389,G833);
  nand GNAME5079(G5079,G4534,G13834);
  nand GNAME5080(G5080,G4535,G36249);
  not GNAME5081(G5081,G4544);
  not GNAME5082(G5082,G4589);
  nand GNAME5083(G5083,G4541,G6694,G6695);
  nand GNAME5084(G5084,G4689,G4541);
  nand GNAME5085(G5085,G4982,G6739,G6740);
  nand GNAME5086(G5086,G4838,G4840,G4842,G4844);
  nand GNAME5087(G5087,G36252,G5081);
  nand GNAME5088(G5088,G6707,G36450);
  nand GNAME5089(G5089,G6710,G36347);
  nand GNAME5090(G5090,G6713,G36315);
  nand GNAME5091(G5091,G6716,G36283);
  or GNAME5092(G5092,G4585,G4557);
  or GNAME5093(G5093,G4569,G4949,G4950);
  nand GNAME5094(G5094,G7125,G4574);
  nand GNAME5095(G5095,G4608,G4548);
  nand GNAME5096(G5096,G5094,G4701);
  nand GNAME5097(G5097,G5093,G13406);
  nand GNAME5098(G5098,G5092,G12609);
  nand GNAME5099(G5099,G5095,G5096,G5097,G5098);
  nand GNAME5100(G5100,G6716,G36284);
  nand GNAME5101(G5101,G6707,G36435);
  nand GNAME5102(G5102,G6710,G36348);
  nand GNAME5103(G5103,G6713,G36316);
  nand GNAME5104(G5104,G6707,G36440);
  nand GNAME5105(G5105,G6710,G36346);
  nand GNAME5106(G5106,G6713,G36314);
  nand GNAME5107(G5107,G6716,G36282);
  nand GNAME5108(G5108,G4637,G4558);
  nand GNAME5109(G5109,G4610,G4548);
  nand GNAME5110(G5110,G5094,G4706);
  nand GNAME5111(G5111,G5093,G13421);
  nand GNAME5112(G5112,G5092,G12624);
  nand GNAME5113(G5113,G5111,G5112,G5110,G5108,G5109);
  nand GNAME5114(G5114,G6716,G36285);
  nand GNAME5115(G5115,G6707,G13901);
  nand GNAME5116(G5116,G6710,G36349);
  nand GNAME5117(G5117,G6713,G36317);
  nand GNAME5118(G5118,G4608,G4558);
  nand GNAME5119(G5119,G4606,G4548);
  nand GNAME5120(G5120,G5094,G4709);
  nand GNAME5121(G5121,G5093,G13356);
  nand GNAME5122(G5122,G5092,G12558);
  nand GNAME5123(G5123,G5121,G5122,G5120,G5118,G5119);
  nand GNAME5124(G5124,G6716,G36286);
  nand GNAME5125(G5125,G6707,G13945);
  nand GNAME5126(G5126,G6710,G36350);
  nand GNAME5127(G5127,G6713,G36318);
  nand GNAME5128(G5128,G4610,G4558);
  nand GNAME5129(G5129,G4609,G4548);
  nand GNAME5130(G5130,G5094,G4712);
  nand GNAME5131(G5131,G5093,G13359);
  nand GNAME5132(G5132,G5092,G12561);
  nand GNAME5133(G5133,G5131,G5132,G5130,G5128,G5129);
  nand GNAME5134(G5134,G6716,G36287);
  nand GNAME5135(G5135,G6707,G13944);
  nand GNAME5136(G5136,G6710,G36351);
  nand GNAME5137(G5137,G6713,G36319);
  nand GNAME5138(G5138,G4606,G4558);
  nand GNAME5139(G5139,G4613,G4548);
  nand GNAME5140(G5140,G5094,G4715);
  nand GNAME5141(G5141,G5093,G13410);
  nand GNAME5142(G5142,G5092,G12613);
  nand GNAME5143(G5143,G5141,G5142,G5140,G5138,G5139);
  nand GNAME5144(G5144,G6716,G36288);
  nand GNAME5145(G5145,G6707,G13943);
  nand GNAME5146(G5146,G6710,G36352);
  nand GNAME5147(G5147,G6713,G36320);
  nand GNAME5148(G5148,G4609,G4558);
  nand GNAME5149(G5149,G4611,G4548);
  nand GNAME5150(G5150,G5094,G4718);
  nand GNAME5151(G5151,G5093,G13409);
  nand GNAME5152(G5152,G5092,G12612);
  nand GNAME5153(G5153,G5151,G5152,G5150,G5148,G5149);
  nand GNAME5154(G5154,G6716,G36289);
  nand GNAME5155(G5155,G6707,G13942);
  nand GNAME5156(G5156,G6710,G36353);
  nand GNAME5157(G5157,G6713,G36321);
  nand GNAME5158(G5158,G4613,G4558);
  nand GNAME5159(G5159,G4612,G4548);
  nand GNAME5160(G5160,G5094,G4721);
  nand GNAME5161(G5161,G5093,G13360);
  nand GNAME5162(G5162,G5092,G12562);
  nand GNAME5163(G5163,G5161,G5162,G5160,G5158,G5159);
  nand GNAME5164(G5164,G6716,G36290);
  nand GNAME5165(G5165,G6707,G13941);
  nand GNAME5166(G5166,G6710,G36354);
  nand GNAME5167(G5167,G6713,G36322);
  nand GNAME5168(G5168,G4611,G4558);
  nand GNAME5169(G5169,G4607,G4548);
  nand GNAME5170(G5170,G5094,G4724);
  nand GNAME5171(G5171,G5093,G13361);
  nand GNAME5172(G5172,G5092,G12563);
  nand GNAME5173(G5173,G5171,G5172,G5170,G5168,G5169);
  nand GNAME5174(G5174,G6716,G36291);
  nand GNAME5175(G5175,G6707,G13940);
  nand GNAME5176(G5176,G6710,G36355);
  nand GNAME5177(G5177,G6713,G36323);
  nand GNAME5178(G5178,G4612,G4558);
  nand GNAME5179(G5179,G4615,G4548);
  nand GNAME5180(G5180,G5094,G4727);
  nand GNAME5181(G5181,G5093,G13408);
  nand GNAME5182(G5182,G5092,G12611);
  nand GNAME5183(G5183,G5181,G5182,G5180,G5178,G5179);
  nand GNAME5184(G5184,G6716,G36292);
  nand GNAME5185(G5185,G6707,G13964);
  nand GNAME5186(G5186,G6710,G36356);
  nand GNAME5187(G5187,G6713,G36324);
  nand GNAME5188(G5188,G4607,G4558);
  nand GNAME5189(G5189,G4614,G4548);
  nand GNAME5190(G5190,G5094,G4730);
  nand GNAME5191(G5191,G5093,G13407);
  nand GNAME5192(G5192,G5092,G12610);
  nand GNAME5193(G5193,G5191,G5192,G5190,G5188,G5189);
  nand GNAME5194(G5194,G6716,G36293);
  nand GNAME5195(G5195,G6707,G13963);
  nand GNAME5196(G5196,G6710,G36357);
  nand GNAME5197(G5197,G6713,G36325);
  nand GNAME5198(G5198,G4615,G4558);
  nand GNAME5199(G5199,G4627,G4548);
  nand GNAME5200(G5200,G5094,G4733);
  nand GNAME5201(G5201,G5093,G13353);
  nand GNAME5202(G5202,G5092,G12555);
  nand GNAME5203(G5203,G5201,G5202,G5200,G5198,G5199);
  nand GNAME5204(G5204,G6716,G36294);
  nand GNAME5205(G5205,G6707,G13962);
  nand GNAME5206(G5206,G6710,G36358);
  nand GNAME5207(G5207,G6713,G36326);
  nand GNAME5208(G5208,G4614,G4558);
  nand GNAME5209(G5209,G4631,G4548);
  nand GNAME5210(G5210,G5094,G4736);
  nand GNAME5211(G5211,G5093,G13354);
  nand GNAME5212(G5212,G5092,G12556);
  nand GNAME5213(G5213,G5211,G5212,G5210,G5208,G5209);
  nand GNAME5214(G5214,G6716,G36295);
  nand GNAME5215(G5215,G6707,G13961);
  nand GNAME5216(G5216,G6710,G36359);
  nand GNAME5217(G5217,G6713,G36327);
  nand GNAME5218(G5218,G4627,G4558);
  nand GNAME5219(G5219,G4629,G4548);
  nand GNAME5220(G5220,G5094,G4739);
  nand GNAME5221(G5221,G5093,G13428);
  nand GNAME5222(G5222,G5092,G12631);
  nand GNAME5223(G5223,G5221,G5222,G5220,G5218,G5219);
  nand GNAME5224(G5224,G6716,G36296);
  nand GNAME5225(G5225,G6707,G13960);
  nand GNAME5226(G5226,G6710,G36360);
  nand GNAME5227(G5227,G6713,G36328);
  nand GNAME5228(G5228,G4631,G4558);
  nand GNAME5229(G5229,G4628,G4548);
  nand GNAME5230(G5230,G5094,G4742);
  nand GNAME5231(G5231,G5093,G13427);
  nand GNAME5232(G5232,G5092,G12630);
  nand GNAME5233(G5233,G5231,G5232,G5230,G5228,G5229);
  nand GNAME5234(G5234,G6716,G36297);
  nand GNAME5235(G5235,G6707,G13959);
  nand GNAME5236(G5236,G6710,G36361);
  nand GNAME5237(G5237,G6713,G36329);
  nand GNAME5238(G5238,G4629,G4558);
  nand GNAME5239(G5239,G4625,G4548);
  nand GNAME5240(G5240,G5094,G4745);
  nand GNAME5241(G5241,G5093,G13355);
  nand GNAME5242(G5242,G5092,G12557);
  nand GNAME5243(G5243,G5241,G5242,G5240,G5238,G5239);
  nand GNAME5244(G5244,G6716,G36298);
  nand GNAME5245(G5245,G6707,G13958);
  nand GNAME5246(G5246,G6710,G36362);
  nand GNAME5247(G5247,G6713,G36330);
  nand GNAME5248(G5248,G4628,G4558);
  nand GNAME5249(G5249,G4630,G4548);
  nand GNAME5250(G5250,G5094,G4748);
  nand GNAME5251(G5251,G5093,G13426);
  nand GNAME5252(G5252,G5092,G12629);
  nand GNAME5253(G5253,G5251,G5252,G5250,G5248,G5249);
  nand GNAME5254(G5254,G6716,G36299);
  nand GNAME5255(G5255,G6707,G13957);
  nand GNAME5256(G5256,G6710,G36363);
  nand GNAME5257(G5257,G6713,G36331);
  nand GNAME5258(G5258,G4625,G4558);
  nand GNAME5259(G5259,G4632,G4548);
  nand GNAME5260(G5260,G5094,G4751);
  nand GNAME5261(G5261,G5093,G13425);
  nand GNAME5262(G5262,G5092,G12628);
  nand GNAME5263(G5263,G5261,G5262,G5260,G5258,G5259);
  nand GNAME5264(G5264,G6716,G36300);
  nand GNAME5265(G5265,G6707,G13956);
  nand GNAME5266(G5266,G6710,G36364);
  nand GNAME5267(G5267,G6713,G36332);
  nand GNAME5268(G5268,G4630,G4558);
  nand GNAME5269(G5269,G4634,G4548);
  nand GNAME5270(G5270,G5094,G4754);
  nand GNAME5271(G5271,G5093,G13424);
  nand GNAME5272(G5272,G5092,G12627);
  nand GNAME5273(G5273,G5271,G5272,G5270,G5268,G5269);
  nand GNAME5274(G5274,G6716,G36301);
  nand GNAME5275(G5275,G6707,G13955);
  nand GNAME5276(G5276,G6710,G36365);
  nand GNAME5277(G5277,G6713,G36333);
  nand GNAME5278(G5278,G4632,G4558);
  nand GNAME5279(G5279,G4633,G4548);
  nand GNAME5280(G5280,G5094,G4757);
  nand GNAME5281(G5281,G5093,G13423);
  nand GNAME5282(G5282,G5092,G12626);
  nand GNAME5283(G5283,G5281,G5282,G5280,G5278,G5279);
  nand GNAME5284(G5284,G6710,G36366);
  nand GNAME5285(G5285,G6713,G36334);
  nand GNAME5286(G5286,G6716,G36302);
  nand GNAME5287(G5287,G6707,G13954);
  nand GNAME5288(G5288,G4634,G4558);
  nand GNAME5289(G5289,G4621,G4548);
  nand GNAME5290(G5290,G5094,G4759);
  nand GNAME5291(G5291,G5093,G13422);
  nand GNAME5292(G5292,G5092,G12625);
  nand GNAME5293(G5293,G5291,G5292,G5290,G5288,G5289);
  nand GNAME5294(G5294,G6710,G36367);
  nand GNAME5295(G5295,G6713,G36335);
  nand GNAME5296(G5296,G6716,G36303);
  nand GNAME5297(G5297,G6707,G13953);
  nand GNAME5298(G5298,G4633,G4558);
  nand GNAME5299(G5299,G4617,G4548);
  nand GNAME5300(G5300,G5094,G4559);
  nand GNAME5301(G5301,G5093,G13420);
  nand GNAME5302(G5302,G5092,G12623);
  nand GNAME5303(G5303,G5301,G5302,G5300,G5298,G5299);
  nand GNAME5304(G5304,G6710,G36368);
  nand GNAME5305(G5305,G6713,G36336);
  nand GNAME5306(G5306,G6716,G36304);
  nand GNAME5307(G5307,G6707,G13952);
  nand GNAME5308(G5308,G4621,G4558);
  nand GNAME5309(G5309,G4622,G4548);
  nand GNAME5310(G5310,G5094,G4560);
  nand GNAME5311(G5311,G5093,G13419);
  nand GNAME5312(G5312,G5092,G12622);
  nand GNAME5313(G5313,G5311,G5312,G5310,G5308,G5309);
  nand GNAME5314(G5314,G6710,G36369);
  nand GNAME5315(G5315,G6713,G36337);
  nand GNAME5316(G5316,G6716,G36305);
  nand GNAME5317(G5317,G6707,G13951);
  nand GNAME5318(G5318,G4617,G4558);
  nand GNAME5319(G5319,G4620,G4548);
  nand GNAME5320(G5320,G5094,G4561);
  nand GNAME5321(G5321,G5093,G13418);
  nand GNAME5322(G5322,G5092,G12621);
  nand GNAME5323(G5323,G5321,G5322,G5320,G5318,G5319);
  nand GNAME5324(G5324,G6710,G36370);
  nand GNAME5325(G5325,G6713,G36338);
  nand GNAME5326(G5326,G6716,G36306);
  nand GNAME5327(G5327,G6707,G13950);
  nand GNAME5328(G5328,G4622,G4558);
  nand GNAME5329(G5329,G4616,G4548);
  nand GNAME5330(G5330,G5094,G4562);
  nand GNAME5331(G5331,G5093,G13417);
  nand GNAME5332(G5332,G5092,G12620);
  nand GNAME5333(G5333,G5331,G5332,G5330,G5328,G5329);
  nand GNAME5334(G5334,G6710,G36371);
  nand GNAME5335(G5335,G6713,G36339);
  nand GNAME5336(G5336,G6716,G36307);
  nand GNAME5337(G5337,G6707,G13949);
  nand GNAME5338(G5338,G4620,G4558);
  nand GNAME5339(G5339,G4619,G4548);
  nand GNAME5340(G5340,G5094,G4563);
  nand GNAME5341(G5341,G5093,G13416);
  nand GNAME5342(G5342,G5092,G12619);
  nand GNAME5343(G5343,G5341,G5342,G5340,G5338,G5339);
  nand GNAME5344(G5344,G6710,G36372);
  nand GNAME5345(G5345,G6713,G36340);
  nand GNAME5346(G5346,G6716,G36308);
  nand GNAME5347(G5347,G6707,G13948);
  nand GNAME5348(G5348,G4616,G4558);
  nand GNAME5349(G5349,G4626,G4548);
  nand GNAME5350(G5350,G5094,G4564);
  nand GNAME5351(G5351,G5093,G13415);
  nand GNAME5352(G5352,G5092,G12618);
  nand GNAME5353(G5353,G5351,G5352,G5350,G5348,G5349);
  nand GNAME5354(G5354,G6710,G36373);
  nand GNAME5355(G5355,G6713,G36341);
  nand GNAME5356(G5356,G6716,G36309);
  nand GNAME5357(G5357,G6707,G13947);
  nand GNAME5358(G5358,G4619,G4558);
  nand GNAME5359(G5359,G4623,G4548);
  nand GNAME5360(G5360,G5094,G4565);
  nand GNAME5361(G5361,G5093,G13414);
  nand GNAME5362(G5362,G5092,G12617);
  nand GNAME5363(G5363,G5361,G5362,G5360,G5358,G5359);
  nand GNAME5364(G5364,G6710,G36374);
  nand GNAME5365(G5365,G6713,G36342);
  nand GNAME5366(G5366,G6716,G36310);
  nand GNAME5367(G5367,G6707,G13946);
  nand GNAME5368(G5368,G4626,G4558);
  nand GNAME5369(G5369,G4624,G4548);
  nand GNAME5370(G5370,G5094,G4566);
  nand GNAME5371(G5371,G5093,G13413);
  nand GNAME5372(G5372,G5092,G12616);
  nand GNAME5373(G5373,G5371,G5372,G5370,G5368,G5369);
  nand GNAME5374(G5374,G6707,G13902);
  nand GNAME5375(G5375,G6710,G36375);
  nand GNAME5376(G5376,G6713,G36343);
  nand GNAME5377(G5377,G6716,G36311);
  nand GNAME5378(G5378,G4623,G4558);
  nand GNAME5379(G5379,G4618,G4548);
  nand GNAME5380(G5380,G5094,G4567);
  nand GNAME5381(G5381,G5093,G13412);
  nand GNAME5382(G5382,G5092,G12615);
  nand GNAME5383(G5383,G5381,G5382,G5380,G5378,G5379);
  nand GNAME5384(G5384,G6710,G36376);
  nand GNAME5385(G5385,G6713,G36344);
  nand GNAME5386(G5386,G6716,G36312);
  nand GNAME5387(G5387,G4542,G6719);
  nand GNAME5388(G5388,G5387,G4959);
  nand GNAME5389(G5389,G4209,G5388);
  nand GNAME5390(G5390,G4624,G4694);
  nand GNAME5391(G5391,G5389,G5390);
  nand GNAME5392(G5392,G5094,G4568);
  nand GNAME5393(G5393,G5093,G13411);
  nand GNAME5394(G5394,G5092,G12614);
  nand GNAME5395(G5395,G5391,G4547);
  nand GNAME5396(G5396,G5392,G5393,G5394,G5395);
  nand GNAME5397(G5397,G6710,G36377);
  nand GNAME5398(G5398,G6713,G36345);
  nand GNAME5399(G5399,G6716,G36313);
  nand GNAME5400(G5400,G4569,G13357);
  nand GNAME5401(G5401,G5094,G4570);
  nand GNAME5402(G5402,G5401,G4971,G5400);
  nand GNAME5403(G5403,G4569,G13358);
  nand GNAME5404(G5404,G5094,G4571);
  nand GNAME5405(G5405,G5404,G4971,G5403);
  nand GNAME5406(G5406,G4573,G4962,G4545);
  nand GNAME5407(G5407,G5406,G4580);
  not GNAME5408(G5408,G4594);
  or GNAME5409(G5409,G4588,G4949,G4950);
  nor GNAME5410(G5410,G6728,G6722);
  or GNAME5411(G5411,G5410,G4557);
  nand GNAME5412(G5412,G4608,G4576);
  nand GNAME5413(G5413,G12609,G4577);
  nand GNAME5414(G5414,G13406,G4579);
  nand GNAME5415(G5415,G36440,G4581);
  nand GNAME5416(G5416,G4701,G4582);
  nand GNAME5417(G5417,G4575,G36346);
  or GNAME5418(G5418,G4961,G4587);
  nand GNAME5419(G5419,G4637,G4583);
  nand GNAME5420(G5420,G4610,G4576);
  nand GNAME5421(G5421,G13421,G4579);
  nand GNAME5422(G5422,G36450,G4581);
  nand GNAME5423(G5423,G4706,G4582);
  nand GNAME5424(G5424,G4608,G4583);
  nand GNAME5425(G5425,G4606,G4576);
  nand GNAME5426(G5426,G12558,G4577);
  nand GNAME5427(G5427,G13356,G4579);
  nand GNAME5428(G5428,G36435,G4581);
  nand GNAME5429(G5429,G4709,G4582);
  nand GNAME5430(G5430,G4575,G36348);
  nand GNAME5431(G5431,G4610,G4583);
  nand GNAME5432(G5432,G4609,G4576);
  nand GNAME5433(G5433,G12561,G4577);
  nand GNAME5434(G5434,G13359,G4579);
  nand GNAME5435(G5435,G13901,G4581);
  nand GNAME5436(G5436,G4712,G4582);
  nand GNAME5437(G5437,G4575,G36349);
  nand GNAME5438(G5438,G4606,G4583);
  nand GNAME5439(G5439,G4613,G4576);
  nand GNAME5440(G5440,G12613,G4577);
  nand GNAME5441(G5441,G13410,G4579);
  nand GNAME5442(G5442,G13945,G4581);
  nand GNAME5443(G5443,G4715,G4582);
  nand GNAME5444(G5444,G4575,G36350);
  nand GNAME5445(G5445,G4609,G4583);
  nand GNAME5446(G5446,G4611,G4576);
  nand GNAME5447(G5447,G12612,G4577);
  nand GNAME5448(G5448,G13409,G4579);
  nand GNAME5449(G5449,G13944,G4581);
  nand GNAME5450(G5450,G4718,G4582);
  nand GNAME5451(G5451,G4575,G36351);
  nand GNAME5452(G5452,G4613,G4583);
  nand GNAME5453(G5453,G4612,G4576);
  nand GNAME5454(G5454,G12562,G4577);
  nand GNAME5455(G5455,G13360,G4579);
  nand GNAME5456(G5456,G13943,G4581);
  nand GNAME5457(G5457,G4721,G4582);
  nand GNAME5458(G5458,G4575,G36352);
  nand GNAME5459(G5459,G4611,G4583);
  nand GNAME5460(G5460,G4607,G4576);
  nand GNAME5461(G5461,G12563,G4577);
  nand GNAME5462(G5462,G13361,G4579);
  nand GNAME5463(G5463,G13942,G4581);
  nand GNAME5464(G5464,G4724,G4582);
  nand GNAME5465(G5465,G4575,G36353);
  nand GNAME5466(G5466,G4612,G4583);
  nand GNAME5467(G5467,G4615,G4576);
  nand GNAME5468(G5468,G12611,G4577);
  nand GNAME5469(G5469,G13408,G4579);
  nand GNAME5470(G5470,G13941,G4581);
  nand GNAME5471(G5471,G4727,G4582);
  nand GNAME5472(G5472,G4575,G36354);
  nand GNAME5473(G5473,G4607,G4583);
  nand GNAME5474(G5474,G4614,G4576);
  nand GNAME5475(G5475,G12610,G4577);
  nand GNAME5476(G5476,G13407,G4579);
  nand GNAME5477(G5477,G13940,G4581);
  nand GNAME5478(G5478,G4730,G4582);
  nand GNAME5479(G5479,G4575,G36355);
  nand GNAME5480(G5480,G4615,G4583);
  nand GNAME5481(G5481,G4627,G4576);
  nand GNAME5482(G5482,G12555,G4577);
  nand GNAME5483(G5483,G13353,G4579);
  nand GNAME5484(G5484,G13964,G4581);
  nand GNAME5485(G5485,G4733,G4582);
  nand GNAME5486(G5486,G4575,G36356);
  nand GNAME5487(G5487,G4614,G4583);
  nand GNAME5488(G5488,G4631,G4576);
  nand GNAME5489(G5489,G12556,G4577);
  nand GNAME5490(G5490,G13354,G4579);
  nand GNAME5491(G5491,G13963,G4581);
  nand GNAME5492(G5492,G4736,G4582);
  nand GNAME5493(G5493,G4575,G36357);
  nand GNAME5494(G5494,G4627,G4583);
  nand GNAME5495(G5495,G4629,G4576);
  nand GNAME5496(G5496,G12631,G4577);
  nand GNAME5497(G5497,G13428,G4579);
  nand GNAME5498(G5498,G13962,G4581);
  nand GNAME5499(G5499,G4739,G4582);
  nand GNAME5500(G5500,G4575,G36358);
  nand GNAME5501(G5501,G4631,G4583);
  nand GNAME5502(G5502,G4628,G4576);
  nand GNAME5503(G5503,G12630,G4577);
  nand GNAME5504(G5504,G13427,G4579);
  nand GNAME5505(G5505,G13961,G4581);
  nand GNAME5506(G5506,G4742,G4582);
  nand GNAME5507(G5507,G4575,G36359);
  nand GNAME5508(G5508,G4629,G4583);
  nand GNAME5509(G5509,G4625,G4576);
  nand GNAME5510(G5510,G12557,G4577);
  nand GNAME5511(G5511,G13355,G4579);
  nand GNAME5512(G5512,G13960,G4581);
  nand GNAME5513(G5513,G4745,G4582);
  nand GNAME5514(G5514,G4575,G36360);
  nand GNAME5515(G5515,G4628,G4583);
  nand GNAME5516(G5516,G4630,G4576);
  nand GNAME5517(G5517,G12629,G4577);
  nand GNAME5518(G5518,G13426,G4579);
  nand GNAME5519(G5519,G13959,G4581);
  nand GNAME5520(G5520,G4748,G4582);
  nand GNAME5521(G5521,G4575,G36361);
  nand GNAME5522(G5522,G4625,G4583);
  nand GNAME5523(G5523,G4632,G4576);
  nand GNAME5524(G5524,G12628,G4577);
  nand GNAME5525(G5525,G13425,G4579);
  nand GNAME5526(G5526,G13958,G4581);
  nand GNAME5527(G5527,G4751,G4582);
  nand GNAME5528(G5528,G4575,G36362);
  nand GNAME5529(G5529,G4630,G4583);
  nand GNAME5530(G5530,G4634,G4576);
  nand GNAME5531(G5531,G12627,G4577);
  nand GNAME5532(G5532,G13424,G4579);
  nand GNAME5533(G5533,G13957,G4581);
  nand GNAME5534(G5534,G4754,G4582);
  nand GNAME5535(G5535,G4575,G36363);
  nand GNAME5536(G5536,G4632,G4583);
  nand GNAME5537(G5537,G4633,G4576);
  nand GNAME5538(G5538,G12626,G4577);
  nand GNAME5539(G5539,G13423,G4579);
  nand GNAME5540(G5540,G13956,G4581);
  nand GNAME5541(G5541,G4757,G4582);
  nand GNAME5542(G5542,G4575,G36364);
  nand GNAME5543(G5543,G4634,G4583);
  nand GNAME5544(G5544,G4621,G4576);
  nand GNAME5545(G5545,G12625,G4577);
  nand GNAME5546(G5546,G13422,G4579);
  nand GNAME5547(G5547,G13955,G4581);
  nand GNAME5548(G5548,G4759,G4582);
  nand GNAME5549(G5549,G4575,G36365);
  nand GNAME5550(G5550,G4633,G4583);
  nand GNAME5551(G5551,G4617,G4576);
  nand GNAME5552(G5552,G12623,G4577);
  nand GNAME5553(G5553,G13420,G4579);
  nand GNAME5554(G5554,G13954,G4581);
  nand GNAME5555(G5555,G4559,G4582);
  nand GNAME5556(G5556,G4575,G36366);
  nand GNAME5557(G5557,G4621,G4583);
  nand GNAME5558(G5558,G4622,G4576);
  nand GNAME5559(G5559,G12622,G4577);
  nand GNAME5560(G5560,G13419,G4579);
  nand GNAME5561(G5561,G13953,G4581);
  nand GNAME5562(G5562,G4560,G4582);
  nand GNAME5563(G5563,G4575,G36367);
  nand GNAME5564(G5564,G4617,G4583);
  nand GNAME5565(G5565,G4620,G4576);
  nand GNAME5566(G5566,G12621,G4577);
  nand GNAME5567(G5567,G13418,G4579);
  nand GNAME5568(G5568,G13952,G4581);
  nand GNAME5569(G5569,G4561,G4582);
  nand GNAME5570(G5570,G4575,G36368);
  nand GNAME5571(G5571,G4622,G4583);
  nand GNAME5572(G5572,G4616,G4576);
  nand GNAME5573(G5573,G12620,G4577);
  nand GNAME5574(G5574,G13417,G4579);
  nand GNAME5575(G5575,G13951,G4581);
  nand GNAME5576(G5576,G4562,G4582);
  nand GNAME5577(G5577,G4575,G36369);
  nand GNAME5578(G5578,G4620,G4583);
  nand GNAME5579(G5579,G4619,G4576);
  nand GNAME5580(G5580,G12619,G4577);
  nand GNAME5581(G5581,G13416,G4579);
  nand GNAME5582(G5582,G13950,G4581);
  nand GNAME5583(G5583,G4563,G4582);
  nand GNAME5584(G5584,G4575,G36370);
  nand GNAME5585(G5585,G4616,G4583);
  nand GNAME5586(G5586,G4626,G4576);
  nand GNAME5587(G5587,G12618,G4577);
  nand GNAME5588(G5588,G13415,G4579);
  nand GNAME5589(G5589,G13949,G4581);
  nand GNAME5590(G5590,G4564,G4582);
  nand GNAME5591(G5591,G4575,G36371);
  nand GNAME5592(G5592,G4619,G4583);
  nand GNAME5593(G5593,G4623,G4576);
  nand GNAME5594(G5594,G12617,G4577);
  nand GNAME5595(G5595,G13414,G4579);
  nand GNAME5596(G5596,G13948,G4581);
  nand GNAME5597(G5597,G4565,G4582);
  nand GNAME5598(G5598,G4575,G36372);
  nand GNAME5599(G5599,G4626,G4583);
  nand GNAME5600(G5600,G4624,G4576);
  nand GNAME5601(G5601,G12616,G4577);
  nand GNAME5602(G5602,G13413,G4579);
  nand GNAME5603(G5603,G13947,G4581);
  nand GNAME5604(G5604,G4566,G4582);
  nand GNAME5605(G5605,G4575,G36373);
  nand GNAME5606(G5606,G4623,G4583);
  nand GNAME5607(G5607,G4618,G4576);
  nand GNAME5608(G5608,G12615,G4577);
  nand GNAME5609(G5609,G13412,G4579);
  nand GNAME5610(G5610,G13946,G4581);
  nand GNAME5611(G5611,G4567,G4582);
  nand GNAME5612(G5612,G4575,G36374);
  nand GNAME5613(G5613,G12614,G4577);
  nand GNAME5614(G5614,G13411,G4579);
  nand GNAME5615(G5615,G13902,G4581);
  nand GNAME5616(G5616,G4568,G4582);
  nand GNAME5617(G5617,G13357,G4588);
  nand GNAME5618(G5618,G5617,G4971);
  nand GNAME5619(G5619,G4570,G4582);
  nand GNAME5620(G5620,G13358,G4588);
  nand GNAME5621(G5621,G5620,G4971);
  nand GNAME5622(G5622,G4571,G4582);
  or GNAME5623(G5623,G4597,G4598);
  or GNAME5624(G5624,G4601,G6736);
  nand GNAME5625(G5625,G12625,G4595);
  nand GNAME5626(G5626,G4596,G13143);
  nand GNAME5627(G5627,G4697,G4599);
  nand GNAME5628(G5628,G5627,G5625,G5626);
  nand GNAME5629(G5629,G4970,G4540);
  nand GNAME5630(G5630,G6700,G5629);
  nand GNAME5631(G5631,G4959,G5630);
  not GNAME5632(G5632,G4603);
  nand GNAME5633(G5633,G4691,G4601);
  nand GNAME5634(G5634,G5633,G4952);
  nand GNAME5635(G5635,G12625,G4592);
  nand GNAME5636(G5636,G6686,G4697);
  nand GNAME5637(G5637,G5628,G4600);
  nand GNAME5638(G5638,G13143,G4602);
  nand GNAME5639(G5639,G5632,G36378);
  nand GNAME5640(G5640,G12626,G4595);
  nand GNAME5641(G5641,G4596,G13186);
  nand GNAME5642(G5642,G4756,G4599);
  nand GNAME5643(G5643,G5642,G5640,G5641);
  nand GNAME5644(G5644,G12626,G4592);
  nand GNAME5645(G5645,G6686,G4756);
  nand GNAME5646(G5646,G5643,G4600);
  nand GNAME5647(G5647,G4602,G13186);
  nand GNAME5648(G5648,G5632,G36379);
  nand GNAME5649(G5649,G12627,G4595);
  nand GNAME5650(G5650,G4596,G13187);
  nand GNAME5651(G5651,G4753,G4599);
  nand GNAME5652(G5652,G5651,G5649,G5650);
  nand GNAME5653(G5653,G12627,G4592);
  nand GNAME5654(G5654,G6686,G4753);
  nand GNAME5655(G5655,G5652,G4600);
  nand GNAME5656(G5656,G4602,G13187);
  nand GNAME5657(G5657,G5632,G36380);
  nand GNAME5658(G5658,G12628,G4595);
  nand GNAME5659(G5659,G4596,G13188);
  nand GNAME5660(G5660,G4750,G4599);
  nand GNAME5661(G5661,G5660,G5658,G5659);
  nand GNAME5662(G5662,G12628,G4592);
  nand GNAME5663(G5663,G6686,G4750);
  nand GNAME5664(G5664,G5661,G4600);
  nand GNAME5665(G5665,G4602,G13188);
  nand GNAME5666(G5666,G5632,G36381);
  nand GNAME5667(G5667,G12629,G4595);
  nand GNAME5668(G5668,G4596,G13142);
  nand GNAME5669(G5669,G4747,G4599);
  nand GNAME5670(G5670,G5669,G5667,G5668);
  nand GNAME5671(G5671,G12629,G4592);
  nand GNAME5672(G5672,G6686,G4747);
  nand GNAME5673(G5673,G5670,G4600);
  nand GNAME5674(G5674,G4602,G13142);
  nand GNAME5675(G5675,G5632,G36382);
  nand GNAME5676(G5676,G12557,G4595);
  nand GNAME5677(G5677,G4596,G13141);
  nand GNAME5678(G5678,G4744,G4599);
  nand GNAME5679(G5679,G5678,G5676,G5677);
  nand GNAME5680(G5680,G12557,G4592);
  nand GNAME5681(G5681,G6686,G4744);
  nand GNAME5682(G5682,G5679,G4600);
  nand GNAME5683(G5683,G4602,G13141);
  nand GNAME5684(G5684,G5632,G36383);
  nand GNAME5685(G5685,G12630,G4595);
  nand GNAME5686(G5686,G4596,G13189);
  nand GNAME5687(G5687,G4741,G4599);
  nand GNAME5688(G5688,G5687,G5685,G5686);
  nand GNAME5689(G5689,G12630,G4592);
  nand GNAME5690(G5690,G6686,G4741);
  nand GNAME5691(G5691,G5688,G4600);
  nand GNAME5692(G5692,G4602,G13189);
  nand GNAME5693(G5693,G5632,G36384);
  nand GNAME5694(G5694,G12631,G4595);
  nand GNAME5695(G5695,G4596,G13190);
  nand GNAME5696(G5696,G4738,G4599);
  nand GNAME5697(G5697,G5696,G5694,G5695);
  nand GNAME5698(G5698,G12631,G4592);
  nand GNAME5699(G5699,G6686,G4738);
  nand GNAME5700(G5700,G5697,G4600);
  nand GNAME5701(G5701,G4602,G13190);
  nand GNAME5702(G5702,G5632,G36385);
  nand GNAME5703(G5703,G12556,G4595);
  nand GNAME5704(G5704,G4596,G13140);
  nand GNAME5705(G5705,G4735,G4599);
  nand GNAME5706(G5706,G5705,G5703,G5704);
  nand GNAME5707(G5707,G12556,G4592);
  nand GNAME5708(G5708,G6686,G4735);
  nand GNAME5709(G5709,G5706,G4600);
  nand GNAME5710(G5710,G4602,G13140);
  nand GNAME5711(G5711,G5632,G36386);
  nand GNAME5712(G5712,G12555,G4595);
  nand GNAME5713(G5713,G4596,G13139);
  nand GNAME5714(G5714,G4732,G4599);
  nand GNAME5715(G5715,G5714,G5712,G5713);
  nand GNAME5716(G5716,G12555,G4592);
  nand GNAME5717(G5717,G6686,G4732);
  nand GNAME5718(G5718,G5715,G4600);
  nand GNAME5719(G5719,G4602,G13139);
  nand GNAME5720(G5720,G5632,G36387);
  nand GNAME5721(G5721,G12610,G4595);
  nand GNAME5722(G5722,G4596,G13178);
  nand GNAME5723(G5723,G4729,G4599);
  nand GNAME5724(G5724,G5723,G5721,G5722);
  nand GNAME5725(G5725,G12610,G4592);
  nand GNAME5726(G5726,G6686,G4729);
  nand GNAME5727(G5727,G5724,G4600);
  nand GNAME5728(G5728,G4602,G13178);
  nand GNAME5729(G5729,G5632,G36388);
  nand GNAME5730(G5730,G12611,G4595);
  nand GNAME5731(G5731,G4596,G13179);
  nand GNAME5732(G5732,G4726,G4599);
  nand GNAME5733(G5733,G5732,G5730,G5731);
  nand GNAME5734(G5734,G12611,G4592);
  nand GNAME5735(G5735,G6686,G4726);
  nand GNAME5736(G5736,G5733,G4600);
  nand GNAME5737(G5737,G4602,G13179);
  nand GNAME5738(G5738,G5632,G36389);
  nand GNAME5739(G5739,G12563,G4595);
  nand GNAME5740(G5740,G4596,G13180);
  nand GNAME5741(G5741,G4723,G4599);
  nand GNAME5742(G5742,G5741,G5739,G5740);
  nand GNAME5743(G5743,G12563,G4592);
  nand GNAME5744(G5744,G6686,G4723);
  nand GNAME5745(G5745,G5742,G4600);
  nand GNAME5746(G5746,G4602,G13180);
  nand GNAME5747(G5747,G5632,G36390);
  nand GNAME5748(G5748,G12562,G4595);
  nand GNAME5749(G5749,G4596,G13181);
  nand GNAME5750(G5750,G4720,G4599);
  nand GNAME5751(G5751,G5750,G5748,G5749);
  nand GNAME5752(G5752,G12562,G4592);
  nand GNAME5753(G5753,G6686,G4720);
  nand GNAME5754(G5754,G5751,G4600);
  nand GNAME5755(G5755,G4602,G13181);
  nand GNAME5756(G5756,G5632,G36391);
  nand GNAME5757(G5757,G12612,G4595);
  nand GNAME5758(G5758,G4596,G13182);
  nand GNAME5759(G5759,G4717,G4599);
  nand GNAME5760(G5760,G5759,G5757,G5758);
  nand GNAME5761(G5761,G12612,G4592);
  nand GNAME5762(G5762,G6686,G4717);
  nand GNAME5763(G5763,G5760,G4600);
  nand GNAME5764(G5764,G4602,G13182);
  nand GNAME5765(G5765,G5632,G36392);
  nand GNAME5766(G5766,G12613,G4595);
  nand GNAME5767(G5767,G4596,G13183);
  nand GNAME5768(G5768,G4714,G4599);
  nand GNAME5769(G5769,G5768,G5766,G5767);
  nand GNAME5770(G5770,G12613,G4592);
  nand GNAME5771(G5771,G6686,G4714);
  nand GNAME5772(G5772,G5769,G4600);
  nand GNAME5773(G5773,G4602,G13183);
  nand GNAME5774(G5774,G5632,G36393);
  nand GNAME5775(G5775,G12561,G4595);
  nand GNAME5776(G5776,G4596,G13184);
  nand GNAME5777(G5777,G4711,G4599);
  nand GNAME5778(G5778,G5777,G5775,G5776);
  nand GNAME5779(G5779,G12561,G4592);
  nand GNAME5780(G5780,G6686,G4711);
  nand GNAME5781(G5781,G5778,G4600);
  nand GNAME5782(G5782,G4602,G13184);
  nand GNAME5783(G5783,G5632,G36394);
  nand GNAME5784(G5784,G12558,G4595);
  nand GNAME5785(G5785,G4596,G13185);
  nand GNAME5786(G5786,G4708,G4599);
  nand GNAME5787(G5787,G5786,G5784,G5785);
  nand GNAME5788(G5788,G12558,G4592);
  nand GNAME5789(G5789,G6686,G4708);
  nand GNAME5790(G5790,G5787,G4600);
  nand GNAME5791(G5791,G4602,G13185);
  nand GNAME5792(G5792,G5632,G36395);
  nand GNAME5793(G5793,G12624,G4595);
  nand GNAME5794(G5794,G4596,G13144);
  nand GNAME5795(G5795,G4705,G4599);
  nand GNAME5796(G5796,G5795,G5793,G5794);
  nand GNAME5797(G5797,G12624,G4592);
  nand GNAME5798(G5798,G6686,G4705);
  nand GNAME5799(G5799,G5796,G4600);
  nand GNAME5800(G5800,G4602,G13144);
  nand GNAME5801(G5801,G5632,G36396);
  nand GNAME5802(G5802,G12609,G4595);
  nand GNAME5803(G5803,G4596,G13177);
  nand GNAME5804(G5804,G4699,G4599);
  nand GNAME5805(G5805,G5804,G5802,G5803);
  nand GNAME5806(G5806,G12609,G4592);
  nand GNAME5807(G5807,G6686,G4699);
  nand GNAME5808(G5808,G5805,G4600);
  nand GNAME5809(G5809,G4602,G13177);
  nand GNAME5810(G5810,G5632,G36397);
  nand GNAME5811(G5811,G7118,G4638);
  nand GNAME5812(G5812,G6731,G4547);
  nand GNAME5813(G5813,G5812,G4958,G4984);
  nand GNAME5814(G5814,G6725,G4645);
  nand GNAME5815(G5815,G6728,G4554);
  nand GNAME5816(G5816,G5815,G4957,G5814);
  nand GNAME5817(G5817,G4639,G4638,G7118);
  nand GNAME5818(G5818,G4635,G7118,G4636,G4641);
  nand GNAME5819(G5819,G4963,G4642);
  nand GNAME5820(G5820,G5811,G4644);
  nand GNAME5821(G5821,G5820,G4939,G5819,G5817,G7120);
  nand GNAME5822(G5822,G7021,G7022,G36460,G4983);
  nand GNAME5823(G5823,G4605,G4938,G4543);
  nand GNAME5824(G5824,G5821,G4593);
  nand GNAME5825(G5825,G5822,G36430);
  nand GNAME5826(G5826,G4628,G4656);
  nand GNAME5827(G5827,G4630,G4657);
  nand GNAME5828(G5828,G4648,G13959);
  nand GNAME5829(G5829,G5828,G5826,G5827);
  nand GNAME5830(G5830,G4550,G4947);
  nand GNAME5831(G5831,G5830,G4695);
  or GNAME5832(G5832,G4650,G4651);
  nand GNAME5833(G5833,G4648,G5832);
  nand GNAME5834(G5834,G5833,G4962);
  and GNAME5835(G5835,G5834,G4543);
  nand GNAME5836(G5836,G6688,G4748);
  nand GNAME5837(G5837,G6687,G13959);
  nand GNAME5838(G5838,G13426,G4654);
  nand GNAME5839(G5839,G12629,G4655);
  nand GNAME5840(G5840,G5829,G4658);
  nand GNAME5841(G5841,G4389,G36431);
  nand GNAME5842(G5842,G4619,G4656);
  nand GNAME5843(G5843,G4623,G4657);
  nand GNAME5844(G5844,G4648,G13948);
  nand GNAME5845(G5845,G5844,G5842,G5843);
  nand GNAME5846(G5846,G4594,G4964);
  nand GNAME5847(G5847,G5846,G4580);
  nand GNAME5848(G5848,G4565,G4659);
  nand GNAME5849(G5849,G13414,G4654);
  nand GNAME5850(G5850,G12617,G4655);
  nand GNAME5851(G5851,G5845,G4658);
  nand GNAME5852(G5852,G6687,G13948);
  nand GNAME5853(G5853,G4389,G36432);
  nand GNAME5854(G5854,G4613,G4656);
  nand GNAME5855(G5855,G4612,G4657);
  nand GNAME5856(G5856,G4648,G13943);
  nand GNAME5857(G5857,G5856,G5854,G5855);
  nand GNAME5858(G5858,G6688,G4721);
  nand GNAME5859(G5859,G6687,G13943);
  nand GNAME5860(G5860,G13360,G4654);
  nand GNAME5861(G5861,G12562,G4655);
  nand GNAME5862(G5862,G5857,G4658);
  nand GNAME5863(G5863,G4389,G36433);
  nand GNAME5864(G5864,G4632,G4656);
  nand GNAME5865(G5865,G4633,G4657);
  nand GNAME5866(G5866,G4648,G13956);
  nand GNAME5867(G5867,G5866,G5864,G5865);
  nand GNAME5868(G5868,G6688,G4757);
  nand GNAME5869(G5869,G6687,G13956);
  nand GNAME5870(G5870,G13423,G4654);
  nand GNAME5871(G5871,G12626,G4655);
  nand GNAME5872(G5872,G5867,G4658);
  nand GNAME5873(G5873,G4389,G36434);
  nand GNAME5874(G5874,G4608,G4656);
  nand GNAME5875(G5875,G4606,G4657);
  nand GNAME5876(G5876,G4648,G36435);
  nand GNAME5877(G5877,G5876,G5874,G5875);
  nand GNAME5878(G5878,G6688,G4709);
  nand GNAME5879(G5879,G6687,G36435);
  nand GNAME5880(G5880,G13356,G4654);
  nand GNAME5881(G5881,G12558,G4655);
  nand GNAME5882(G5882,G5877,G4658);
  nand GNAME5883(G5883,G4389,G36435);
  nand GNAME5884(G5884,G4614,G4656);
  nand GNAME5885(G5885,G4631,G4657);
  nand GNAME5886(G5886,G4648,G13963);
  nand GNAME5887(G5887,G5886,G5884,G5885);
  nand GNAME5888(G5888,G6688,G4736);
  nand GNAME5889(G5889,G6687,G13963);
  nand GNAME5890(G5890,G13354,G4654);
  nand GNAME5891(G5891,G12556,G4655);
  nand GNAME5892(G5892,G5887,G4658);
  nand GNAME5893(G5893,G4389,G36436);
  nand GNAME5894(G5894,G4617,G4656);
  nand GNAME5895(G5895,G4620,G4657);
  nand GNAME5896(G5896,G4648,G13952);
  nand GNAME5897(G5897,G5896,G5894,G5895);
  nand GNAME5898(G5898,G4561,G4659);
  nand GNAME5899(G5899,G13418,G4654);
  nand GNAME5900(G5900,G12621,G4655);
  nand GNAME5901(G5901,G5897,G4658);
  nand GNAME5902(G5902,G6687,G13952);
  nand GNAME5903(G5903,G4389,G36437);
  nand GNAME5904(G5904,G4631,G4656);
  nand GNAME5905(G5905,G4628,G4657);
  nand GNAME5906(G5906,G4648,G13961);
  nand GNAME5907(G5907,G5906,G5904,G5905);
  nand GNAME5908(G5908,G6688,G4742);
  nand GNAME5909(G5909,G6687,G13961);
  nand GNAME5910(G5910,G13427,G4654);
  nand GNAME5911(G5911,G12630,G4655);
  nand GNAME5912(G5912,G5907,G4658);
  nand GNAME5913(G5913,G4389,G36438);
  nand GNAME5914(G5914,G4633,G4656);
  nand GNAME5915(G5915,G4617,G4657);
  nand GNAME5916(G5916,G4648,G13954);
  nand GNAME5917(G5917,G5916,G5914,G5915);
  nand GNAME5918(G5918,G4559,G4659);
  nand GNAME5919(G5919,G13420,G4654);
  nand GNAME5920(G5920,G12623,G4655);
  nand GNAME5921(G5921,G5917,G4658);
  nand GNAME5922(G5922,G6687,G13954);
  nand GNAME5923(G5923,G4389,G36439);
  or GNAME5924(G5924,G4647,G4658);
  nand GNAME5925(G5925,G4648,G5924);
  nand GNAME5926(G5926,G5925,G4652);
  nand GNAME5927(G5927,G4658,G4608,G4657);
  nand GNAME5928(G5928,G6688,G4701);
  nand GNAME5929(G5929,G5926,G36440);
  nand GNAME5930(G5930,G13406,G4654);
  nand GNAME5931(G5931,G12609,G4655);
  nand GNAME5932(G5932,G4389,G36440);
  nand GNAME5933(G5933,G4607,G4656);
  nand GNAME5934(G5934,G4614,G4657);
  nand GNAME5935(G5935,G4648,G13940);
  nand GNAME5936(G5936,G5935,G5933,G5934);
  nand GNAME5937(G5937,G6688,G4730);
  nand GNAME5938(G5938,G6687,G13940);
  nand GNAME5939(G5939,G13407,G4654);
  nand GNAME5940(G5940,G12610,G4655);
  nand GNAME5941(G5941,G5936,G4658);
  nand GNAME5942(G5942,G4389,G36441);
  nand GNAME5943(G5943,G4606,G4656);
  nand GNAME5944(G5944,G4613,G4657);
  nand GNAME5945(G5945,G4648,G13945);
  nand GNAME5946(G5946,G5945,G5943,G5944);
  nand GNAME5947(G5947,G6688,G4715);
  nand GNAME5948(G5948,G6687,G13945);
  nand GNAME5949(G5949,G13410,G4654);
  nand GNAME5950(G5950,G12613,G4655);
  nand GNAME5951(G5951,G5946,G4658);
  nand GNAME5952(G5952,G4389,G36442);
  nand GNAME5953(G5953,G4620,G4656);
  nand GNAME5954(G5954,G4619,G4657);
  nand GNAME5955(G5955,G4648,G13950);
  nand GNAME5956(G5956,G5955,G5953,G5954);
  nand GNAME5957(G5957,G4563,G4659);
  nand GNAME5958(G5958,G13416,G4654);
  nand GNAME5959(G5959,G12619,G4655);
  nand GNAME5960(G5960,G5956,G4658);
  nand GNAME5961(G5961,G6687,G13950);
  nand GNAME5962(G5962,G4389,G36443);
  nand GNAME5963(G5963,G4630,G4656);
  nand GNAME5964(G5964,G4634,G4657);
  nand GNAME5965(G5965,G4648,G13957);
  nand GNAME5966(G5966,G5965,G5963,G5964);
  nand GNAME5967(G5967,G6688,G4754);
  nand GNAME5968(G5968,G6687,G13957);
  nand GNAME5969(G5969,G13424,G4654);
  nand GNAME5970(G5970,G12627,G4655);
  nand GNAME5971(G5971,G5966,G4658);
  nand GNAME5972(G5972,G4389,G36444);
  nand GNAME5973(G5973,G4609,G4656);
  nand GNAME5974(G5974,G4611,G4657);
  nand GNAME5975(G5975,G4648,G13944);
  nand GNAME5976(G5976,G5975,G5973,G5974);
  nand GNAME5977(G5977,G6688,G4718);
  nand GNAME5978(G5978,G6687,G13944);
  nand GNAME5979(G5979,G13409,G4654);
  nand GNAME5980(G5980,G12612,G4655);
  nand GNAME5981(G5981,G5976,G4658);
  nand GNAME5982(G5982,G4389,G36445);
  nand GNAME5983(G5983,G4625,G4656);
  nand GNAME5984(G5984,G4632,G4657);
  nand GNAME5985(G5985,G4648,G13958);
  nand GNAME5986(G5986,G5985,G5983,G5984);
  nand GNAME5987(G5987,G6688,G4751);
  nand GNAME5988(G5988,G6687,G13958);
  nand GNAME5989(G5989,G13425,G4654);
  nand GNAME5990(G5990,G12628,G4655);
  nand GNAME5991(G5991,G5986,G4658);
  nand GNAME5992(G5992,G4389,G36446);
  nand GNAME5993(G5993,G4616,G4656);
  nand GNAME5994(G5994,G4626,G4657);
  nand GNAME5995(G5995,G4648,G13949);
  nand GNAME5996(G5996,G5995,G5993,G5994);
  nand GNAME5997(G5997,G4564,G4659);
  nand GNAME5998(G5998,G13415,G4654);
  nand GNAME5999(G5999,G12618,G4655);
  nand GNAME6000(G6000,G5996,G4658);
  nand GNAME6001(G6001,G6687,G13949);
  nand GNAME6002(G6002,G4389,G36447);
  nand GNAME6003(G6003,G4627,G4656);
  nand GNAME6004(G6004,G4629,G4657);
  nand GNAME6005(G6005,G4648,G13962);
  nand GNAME6006(G6006,G6005,G6003,G6004);
  nand GNAME6007(G6007,G6688,G4739);
  nand GNAME6008(G6008,G6687,G13962);
  nand GNAME6009(G6009,G13428,G4654);
  nand GNAME6010(G6010,G12631,G4655);
  nand GNAME6011(G6011,G6006,G4658);
  nand GNAME6012(G6012,G4389,G36448);
  nand GNAME6013(G6013,G4621,G4656);
  nand GNAME6014(G6014,G4622,G4657);
  nand GNAME6015(G6015,G4648,G13953);
  nand GNAME6016(G6016,G6015,G6013,G6014);
  nand GNAME6017(G6017,G4560,G4659);
  nand GNAME6018(G6018,G13419,G4654);
  nand GNAME6019(G6019,G12622,G4655);
  nand GNAME6020(G6020,G6016,G4658);
  nand GNAME6021(G6021,G6687,G13953);
  nand GNAME6022(G6022,G4389,G36449);
  nand GNAME6023(G6023,G4637,G4656);
  nand GNAME6024(G6024,G4610,G4657);
  nand GNAME6025(G6025,G4648,G36450);
  nand GNAME6026(G6026,G6025,G6023,G6024);
  nand GNAME6027(G6027,G6688,G4706);
  nand GNAME6028(G6028,G6687,G36450);
  nand GNAME6029(G6029,G13421,G4654);
  nand GNAME6030(G6030,G12624,G4655);
  nand GNAME6031(G6031,G6026,G4658);
  nand GNAME6032(G6032,G4389,G36450);
  nand GNAME6033(G6033,G4612,G4656);
  nand GNAME6034(G6034,G4615,G4657);
  nand GNAME6035(G6035,G4648,G13941);
  nand GNAME6036(G6036,G6035,G6033,G6034);
  nand GNAME6037(G6037,G6688,G4727);
  nand GNAME6038(G6038,G6687,G13941);
  nand GNAME6039(G6039,G13408,G4654);
  nand GNAME6040(G6040,G12611,G4655);
  nand GNAME6041(G6041,G6036,G4658);
  nand GNAME6042(G6042,G4389,G36451);
  nand GNAME6043(G6043,G4623,G4656);
  nand GNAME6044(G6044,G4618,G4657);
  nand GNAME6045(G6045,G4648,G13946);
  nand GNAME6046(G6046,G6045,G6043,G6044);
  nand GNAME6047(G6047,G4567,G4659);
  nand GNAME6048(G6048,G13412,G4654);
  nand GNAME6049(G6049,G12615,G4655);
  nand GNAME6050(G6050,G6046,G4658);
  nand GNAME6051(G6051,G6687,G13946);
  nand GNAME6052(G6052,G4389,G36452);
  nand GNAME6053(G6053,G4634,G4656);
  nand GNAME6054(G6054,G4621,G4657);
  nand GNAME6055(G6055,G4648,G13955);
  nand GNAME6056(G6056,G6055,G6053,G6054);
  nand GNAME6057(G6057,G6688,G4759);
  nand GNAME6058(G6058,G6687,G13955);
  nand GNAME6059(G6059,G13422,G4654);
  nand GNAME6060(G6060,G12625,G4655);
  nand GNAME6061(G6061,G6056,G4658);
  nand GNAME6062(G6062,G4389,G36453);
  nand GNAME6063(G6063,G4610,G4656);
  nand GNAME6064(G6064,G4609,G4657);
  nand GNAME6065(G6065,G4648,G13901);
  nand GNAME6066(G6066,G6065,G6063,G6064);
  nand GNAME6067(G6067,G6688,G4712);
  nand GNAME6068(G6068,G6687,G13901);
  nand GNAME6069(G6069,G13359,G4654);
  nand GNAME6070(G6070,G12561,G4655);
  nand GNAME6071(G6071,G6066,G4658);
  nand GNAME6072(G6072,G4389,G36454);
  nand GNAME6073(G6073,G4615,G4656);
  nand GNAME6074(G6074,G4627,G4657);
  nand GNAME6075(G6075,G4648,G13964);
  nand GNAME6076(G6076,G6075,G6073,G6074);
  nand GNAME6077(G6077,G6688,G4733);
  nand GNAME6078(G6078,G6687,G13964);
  nand GNAME6079(G6079,G13353,G4654);
  nand GNAME6080(G6080,G12555,G4655);
  nand GNAME6081(G6081,G6076,G4658);
  nand GNAME6082(G6082,G4389,G36455);
  nand GNAME6083(G6083,G4622,G4656);
  nand GNAME6084(G6084,G4616,G4657);
  nand GNAME6085(G6085,G4648,G13951);
  nand GNAME6086(G6086,G6085,G6083,G6084);
  nand GNAME6087(G6087,G4562,G4659);
  nand GNAME6088(G6088,G13417,G4654);
  nand GNAME6089(G6089,G12620,G4655);
  nand GNAME6090(G6090,G6086,G4658);
  nand GNAME6091(G6091,G6687,G13951);
  nand GNAME6092(G6092,G4389,G36456);
  nand GNAME6093(G6093,G4629,G4656);
  nand GNAME6094(G6094,G4625,G4657);
  nand GNAME6095(G6095,G4648,G13960);
  nand GNAME6096(G6096,G6095,G6093,G6094);
  nand GNAME6097(G6097,G6688,G4745);
  nand GNAME6098(G6098,G6687,G13960);
  nand GNAME6099(G6099,G13355,G4654);
  nand GNAME6100(G6100,G12557,G4655);
  nand GNAME6101(G6101,G6096,G4658);
  nand GNAME6102(G6102,G4389,G36457);
  nand GNAME6103(G6103,G4626,G4656);
  nand GNAME6104(G6104,G4624,G4657);
  nand GNAME6105(G6105,G4648,G13947);
  nand GNAME6106(G6106,G6105,G6103,G6104);
  nand GNAME6107(G6107,G4566,G4659);
  nand GNAME6108(G6108,G13413,G4654);
  nand GNAME6109(G6109,G12616,G4655);
  nand GNAME6110(G6110,G6106,G4658);
  nand GNAME6111(G6111,G6687,G13947);
  nand GNAME6112(G6112,G4389,G36458);
  nand GNAME6113(G6113,G4611,G4656);
  nand GNAME6114(G6114,G4607,G4657);
  nand GNAME6115(G6115,G4648,G13942);
  nand GNAME6116(G6116,G6115,G6113,G6114);
  nand GNAME6117(G6117,G6688,G4724);
  nand GNAME6118(G6118,G6687,G13942);
  nand GNAME6119(G6119,G13361,G4654);
  nand GNAME6120(G6120,G12563,G4655);
  nand GNAME6121(G6121,G6116,G4658);
  nand GNAME6122(G6122,G4389,G36459);
  or GNAME6123(G6123,G4685,G4686);
  nand GNAME6124(G6124,G4942,G4944,G4975,G4976);
  nand GNAME6125(G6125,G4684,G4730);
  nand GNAME6126(G6126,G4615,G6124);
  nand GNAME6127(G6127,G6123,G4729);
  nand GNAME6128(G6128,G36323,G4673);
  nand GNAME6129(G6129,G36355,G4674);
  nand GNAME6130(G6130,G4684,G4727);
  nand GNAME6131(G6131,G4607,G6124);
  nand GNAME6132(G6132,G6123,G4726);
  nand GNAME6133(G6133,G36322,G4673);
  nand GNAME6134(G6134,G36354,G4674);
  nand GNAME6135(G6135,G4684,G4724);
  nand GNAME6136(G6136,G4612,G6124);
  nand GNAME6137(G6137,G6123,G4723);
  nand GNAME6138(G6138,G36321,G4673);
  nand GNAME6139(G6139,G36353,G4674);
  nand GNAME6140(G6140,G4684,G4721);
  nand GNAME6141(G6141,G4611,G6124);
  nand GNAME6142(G6142,G6123,G4720);
  nand GNAME6143(G6143,G36320,G4673);
  nand GNAME6144(G6144,G36352,G4674);
  nand GNAME6145(G6145,G4684,G4718);
  nand GNAME6146(G6146,G4613,G6124);
  nand GNAME6147(G6147,G6123,G4717);
  nand GNAME6148(G6148,G36319,G4673);
  nand GNAME6149(G6149,G36351,G4674);
  nand GNAME6150(G6150,G4684,G4715);
  nand GNAME6151(G6151,G4609,G6124);
  nand GNAME6152(G6152,G6123,G4714);
  nand GNAME6153(G6153,G36318,G4673);
  nand GNAME6154(G6154,G36350,G4674);
  nand GNAME6155(G6155,G4976,G4975);
  nand GNAME6156(G6156,G4944,G4942);
  nand GNAME6157(G6157,G4624,G6156);
  nand GNAME6158(G6158,G4666,G4567);
  nand GNAME6159(G6159,G4618,G6155);
  nand GNAME6160(G6160,G4667,G4568);
  nand GNAME6161(G6161,G4684,G4712);
  nand GNAME6162(G6162,G4606,G6124);
  nand GNAME6163(G6163,G6123,G4711);
  nand GNAME6164(G6164,G36317,G4673);
  nand GNAME6165(G6165,G36349,G4674);
  nand GNAME6166(G6166,G4624,G6124);
  nand GNAME6167(G6167,G4684,G4567);
  nand GNAME6168(G6168,G4623,G6124);
  nand GNAME6169(G6169,G4684,G4566);
  nand GNAME6170(G6170,G4626,G6124);
  nand GNAME6171(G6171,G4684,G4565);
  nand GNAME6172(G6172,G4619,G6124);
  nand GNAME6173(G6173,G4684,G4564);
  nand GNAME6174(G6174,G4616,G6124);
  nand GNAME6175(G6175,G4684,G4563);
  nand GNAME6176(G6176,G4620,G6124);
  nand GNAME6177(G6177,G4684,G4562);
  nand GNAME6178(G6178,G4622,G6124);
  nand GNAME6179(G6179,G4684,G4561);
  nand GNAME6180(G6180,G4617,G6124);
  nand GNAME6181(G6181,G4684,G4560);
  nand GNAME6182(G6182,G4621,G6124);
  nand GNAME6183(G6183,G4684,G4559);
  nand GNAME6184(G6184,G4684,G4709);
  nand GNAME6185(G6185,G4610,G6124);
  nand GNAME6186(G6186,G6123,G4708);
  nand GNAME6187(G6187,G36316,G4673);
  nand GNAME6188(G6188,G36348,G4674);
  nand GNAME6189(G6189,G4684,G4759);
  nand GNAME6190(G6190,G4633,G6124);
  nand GNAME6191(G6191,G36333,G4673);
  nand GNAME6192(G6192,G36365,G4674);
  nand GNAME6193(G6193,G4684,G4757);
  nand GNAME6194(G6194,G4634,G6124);
  nand GNAME6195(G6195,G6123,G4756);
  nand GNAME6196(G6196,G36332,G4673);
  nand GNAME6197(G6197,G36364,G4674);
  nand GNAME6198(G6198,G4684,G4754);
  nand GNAME6199(G6199,G4632,G6124);
  nand GNAME6200(G6200,G6123,G4753);
  nand GNAME6201(G6201,G36331,G4673);
  nand GNAME6202(G6202,G36363,G4674);
  nand GNAME6203(G6203,G4684,G4751);
  nand GNAME6204(G6204,G4630,G6124);
  nand GNAME6205(G6205,G6123,G4750);
  nand GNAME6206(G6206,G36330,G4673);
  nand GNAME6207(G6207,G36362,G4674);
  nand GNAME6208(G6208,G4684,G4748);
  nand GNAME6209(G6209,G4625,G6124);
  nand GNAME6210(G6210,G6123,G4747);
  nand GNAME6211(G6211,G36329,G4673);
  nand GNAME6212(G6212,G36361,G4674);
  nand GNAME6213(G6213,G4684,G4745);
  nand GNAME6214(G6214,G4628,G6124);
  nand GNAME6215(G6215,G6123,G4744);
  nand GNAME6216(G6216,G36328,G4673);
  nand GNAME6217(G6217,G36360,G4674);
  nand GNAME6218(G6218,G4684,G4742);
  nand GNAME6219(G6219,G4629,G6124);
  nand GNAME6220(G6220,G6123,G4741);
  nand GNAME6221(G6221,G36327,G4673);
  nand GNAME6222(G6222,G36359,G4674);
  nand GNAME6223(G6223,G4684,G4739);
  nand GNAME6224(G6224,G4631,G6124);
  nand GNAME6225(G6225,G6123,G4738);
  nand GNAME6226(G6226,G36326,G4673);
  nand GNAME6227(G6227,G36358,G4674);
  nand GNAME6228(G6228,G4684,G4736);
  nand GNAME6229(G6229,G4627,G6124);
  nand GNAME6230(G6230,G6123,G4735);
  nand GNAME6231(G6231,G36325,G4673);
  nand GNAME6232(G6232,G36357,G4674);
  nand GNAME6233(G6233,G4684,G4733);
  nand GNAME6234(G6234,G4614,G6124);
  nand GNAME6235(G6235,G6123,G4732);
  nand GNAME6236(G6236,G36324,G4673);
  nand GNAME6237(G6237,G36356,G4674);
  nand GNAME6238(G6238,G4684,G4706);
  nand GNAME6239(G6239,G4608,G6124);
  nand GNAME6240(G6240,G6123,G4705);
  nand GNAME6241(G6241,G36315,G4673);
  nand GNAME6242(G6242,G36347,G4674);
  nand GNAME6243(G6243,G4684,G4701);
  nand GNAME6244(G6244,G4637,G6124);
  nand GNAME6245(G6245,G6123,G4699);
  nand GNAME6246(G6246,G36314,G4673);
  nand GNAME6247(G6247,G36346,G4674);
  nor GNAME6248(G6248,G5082,G4643);
  nand GNAME6249(G6249,G4954,G4671,G4981,G4675);
  nand GNAME6250(G6250,G4676,G4567);
  nand GNAME6251(G6251,G4677,G4568);
  or GNAME6252(G6252,G4676,G4677);
  or GNAME6253(G6253,G4679,G4678);
  nand GNAME6254(G6254,G6253,G4730);
  nand GNAME6255(G6255,G4615,G6252);
  nand GNAME6256(G6256,G6253,G4727);
  nand GNAME6257(G6257,G4607,G6252);
  nand GNAME6258(G6258,G6253,G4724);
  nand GNAME6259(G6259,G4612,G6252);
  nand GNAME6260(G6260,G6253,G4721);
  nand GNAME6261(G6261,G4611,G6252);
  nand GNAME6262(G6262,G6253,G4718);
  nand GNAME6263(G6263,G4613,G6252);
  nand GNAME6264(G6264,G6253,G4715);
  nand GNAME6265(G6265,G4609,G6252);
  nand GNAME6266(G6266,G4624,G4676);
  nand GNAME6267(G6267,G4618,G4677);
  nand GNAME6268(G6268,G4567,G4678);
  nand GNAME6269(G6269,G4571,G4679);
  nand GNAME6270(G6270,G4570,G4679);
  nand GNAME6271(G6271,G6253,G4712);
  nand GNAME6272(G6272,G4606,G6252);
  nand GNAME6273(G6273,G4568,G4679);
  nand GNAME6274(G6274,G6253,G4567);
  nand GNAME6275(G6275,G4624,G6252);
  nand GNAME6276(G6276,G6253,G4566);
  nand GNAME6277(G6277,G4623,G6252);
  nand GNAME6278(G6278,G6253,G4565);
  nand GNAME6279(G6279,G4626,G6252);
  nand GNAME6280(G6280,G6253,G4564);
  nand GNAME6281(G6281,G4619,G6252);
  nand GNAME6282(G6282,G6253,G4563);
  nand GNAME6283(G6283,G4616,G6252);
  nand GNAME6284(G6284,G6253,G4562);
  nand GNAME6285(G6285,G4620,G6252);
  nand GNAME6286(G6286,G6253,G4561);
  nand GNAME6287(G6287,G4622,G6252);
  nand GNAME6288(G6288,G6253,G4560);
  nand GNAME6289(G6289,G4617,G6252);
  nand GNAME6290(G6290,G6253,G4559);
  nand GNAME6291(G6291,G4621,G6252);
  nand GNAME6292(G6292,G6253,G4709);
  nand GNAME6293(G6293,G4610,G6252);
  nand GNAME6294(G6294,G6253,G4759);
  nand GNAME6295(G6295,G4633,G6252);
  nand GNAME6296(G6296,G6253,G4757);
  nand GNAME6297(G6297,G4634,G6252);
  nand GNAME6298(G6298,G6253,G4754);
  nand GNAME6299(G6299,G4632,G6252);
  nand GNAME6300(G6300,G6253,G4751);
  nand GNAME6301(G6301,G4630,G6252);
  nand GNAME6302(G6302,G6253,G4748);
  nand GNAME6303(G6303,G4625,G6252);
  nand GNAME6304(G6304,G6253,G4745);
  nand GNAME6305(G6305,G4628,G6252);
  nand GNAME6306(G6306,G6253,G4742);
  nand GNAME6307(G6307,G4629,G6252);
  nand GNAME6308(G6308,G6253,G4739);
  nand GNAME6309(G6309,G4631,G6252);
  nand GNAME6310(G6310,G6253,G4736);
  nand GNAME6311(G6311,G4627,G6252);
  nand GNAME6312(G6312,G6253,G4733);
  nand GNAME6313(G6313,G4614,G6252);
  nand GNAME6314(G6314,G6253,G4706);
  nand GNAME6315(G6315,G4608,G6252);
  nand GNAME6316(G6316,G6253,G4701);
  nand GNAME6317(G6317,G4637,G6252);
  nand GNAME6318(G6318,G4672,G4952);
  nand GNAME6319(G6319,G6318,G36323);
  nand GNAME6320(G6320,G4700,G36355);
  nand GNAME6321(G6321,G6318,G36322);
  nand GNAME6322(G6322,G4700,G36354);
  nand GNAME6323(G6323,G6318,G36321);
  nand GNAME6324(G6324,G4700,G36353);
  nand GNAME6325(G6325,G6318,G36320);
  nand GNAME6326(G6326,G4700,G36352);
  nand GNAME6327(G6327,G6318,G36319);
  nand GNAME6328(G6328,G4700,G36351);
  nand GNAME6329(G6329,G6318,G36318);
  nand GNAME6330(G6330,G4700,G36350);
  nand GNAME6331(G6331,G6318,G36317);
  nand GNAME6332(G6332,G4700,G36349);
  nand GNAME6333(G6333,G6318,G36316);
  nand GNAME6334(G6334,G4700,G36348);
  nand GNAME6335(G6335,G6318,G36333);
  nand GNAME6336(G6336,G4700,G36365);
  nand GNAME6337(G6337,G6318,G36332);
  nand GNAME6338(G6338,G4700,G36364);
  nand GNAME6339(G6339,G6318,G36331);
  nand GNAME6340(G6340,G4700,G36363);
  nand GNAME6341(G6341,G6318,G36330);
  nand GNAME6342(G6342,G4700,G36362);
  nand GNAME6343(G6343,G6318,G36329);
  nand GNAME6344(G6344,G4700,G36361);
  nand GNAME6345(G6345,G6318,G36328);
  nand GNAME6346(G6346,G4700,G36360);
  nand GNAME6347(G6347,G6318,G36327);
  nand GNAME6348(G6348,G4700,G36359);
  nand GNAME6349(G6349,G6318,G36326);
  nand GNAME6350(G6350,G4700,G36358);
  nand GNAME6351(G6351,G6318,G36325);
  nand GNAME6352(G6352,G4700,G36357);
  nand GNAME6353(G6353,G6318,G36324);
  nand GNAME6354(G6354,G4700,G36356);
  nand GNAME6355(G6355,G6318,G36315);
  nand GNAME6356(G6356,G4700,G36347);
  nand GNAME6357(G6357,G6318,G36314);
  nand GNAME6358(G6358,G4700,G36346);
  nand GNAME6359(G6359,G4691,G4604);
  nand GNAME6360(G6360,G6359,G4951);
  or GNAME6361(G6361,G6725,G4649);
  nand GNAME6362(G6362,G4681,G7123);
  nand GNAME6363(G6363,G6362,G4730);
  nand GNAME6364(G6364,G4615,G6360);
  nand GNAME6365(G6365,G6700,G4607);
  nand GNAME6366(G6366,G6362,G4727);
  nand GNAME6367(G6367,G4607,G6360);
  nand GNAME6368(G6368,G6700,G4612);
  nand GNAME6369(G6369,G6362,G4724);
  nand GNAME6370(G6370,G4612,G6360);
  nand GNAME6371(G6371,G6700,G4611);
  nand GNAME6372(G6372,G6362,G4721);
  nand GNAME6373(G6373,G4611,G6360);
  nand GNAME6374(G6374,G6700,G4613);
  nand GNAME6375(G6375,G6362,G4718);
  nand GNAME6376(G6376,G4613,G6360);
  nand GNAME6377(G6377,G6700,G4609);
  nand GNAME6378(G6378,G6362,G4715);
  nand GNAME6379(G6379,G4609,G6360);
  nand GNAME6380(G6380,G6700,G4606);
  nand GNAME6381(G6381,G6362,G4571);
  nand GNAME6382(G6382,G4207,G6360);
  nand GNAME6383(G6383,G6362,G4570);
  nand GNAME6384(G6384,G4209,G6360);
  nand GNAME6385(G6385,G6362,G4712);
  nand GNAME6386(G6386,G4606,G6360);
  nand GNAME6387(G6387,G6700,G4610);
  nand GNAME6388(G6388,G6362,G4568);
  nand GNAME6389(G6389,G4618,G6360);
  nand GNAME6390(G6390,G6700,G4624);
  nand GNAME6391(G6391,G6362,G4567);
  nand GNAME6392(G6392,G4624,G6360);
  nand GNAME6393(G6393,G6700,G4623);
  nand GNAME6394(G6394,G6362,G4566);
  nand GNAME6395(G6395,G4623,G6360);
  nand GNAME6396(G6396,G6700,G4626);
  nand GNAME6397(G6397,G6362,G4565);
  nand GNAME6398(G6398,G4626,G6360);
  nand GNAME6399(G6399,G6700,G4619);
  nand GNAME6400(G6400,G6362,G4564);
  nand GNAME6401(G6401,G4619,G6360);
  nand GNAME6402(G6402,G6700,G4616);
  nand GNAME6403(G6403,G6362,G4563);
  nand GNAME6404(G6404,G4616,G6360);
  nand GNAME6405(G6405,G6700,G4620);
  nand GNAME6406(G6406,G6362,G4562);
  nand GNAME6407(G6407,G4620,G6360);
  nand GNAME6408(G6408,G6700,G4622);
  nand GNAME6409(G6409,G6362,G4561);
  nand GNAME6410(G6410,G4622,G6360);
  nand GNAME6411(G6411,G6700,G4617);
  nand GNAME6412(G6412,G6362,G4560);
  nand GNAME6413(G6413,G4617,G6360);
  nand GNAME6414(G6414,G6700,G4621);
  nand GNAME6415(G6415,G6362,G4559);
  nand GNAME6416(G6416,G4621,G6360);
  nand GNAME6417(G6417,G6700,G4633);
  nand GNAME6418(G6418,G6362,G4709);
  nand GNAME6419(G6419,G4610,G6360);
  nand GNAME6420(G6420,G6700,G4608);
  nand GNAME6421(G6421,G6362,G4759);
  nand GNAME6422(G6422,G4633,G6360);
  nand GNAME6423(G6423,G6700,G4634);
  nand GNAME6424(G6424,G6362,G4757);
  nand GNAME6425(G6425,G4634,G6360);
  nand GNAME6426(G6426,G6700,G4632);
  nand GNAME6427(G6427,G6362,G4754);
  nand GNAME6428(G6428,G4632,G6360);
  nand GNAME6429(G6429,G6700,G4630);
  nand GNAME6430(G6430,G6362,G4751);
  nand GNAME6431(G6431,G4630,G6360);
  nand GNAME6432(G6432,G6700,G4625);
  nand GNAME6433(G6433,G6362,G4748);
  nand GNAME6434(G6434,G4625,G6360);
  nand GNAME6435(G6435,G6700,G4628);
  nand GNAME6436(G6436,G6362,G4745);
  nand GNAME6437(G6437,G4628,G6360);
  nand GNAME6438(G6438,G6700,G4629);
  nand GNAME6439(G6439,G6362,G4742);
  nand GNAME6440(G6440,G4629,G6360);
  nand GNAME6441(G6441,G6700,G4631);
  nand GNAME6442(G6442,G6362,G4739);
  nand GNAME6443(G6443,G4631,G6360);
  nand GNAME6444(G6444,G6700,G4627);
  nand GNAME6445(G6445,G6362,G4736);
  nand GNAME6446(G6446,G4627,G6360);
  nand GNAME6447(G6447,G6700,G4614);
  nand GNAME6448(G6448,G6362,G4733);
  nand GNAME6449(G6449,G4614,G6360);
  nand GNAME6450(G6450,G6700,G4615);
  nand GNAME6451(G6451,G6362,G4706);
  nand GNAME6452(G6452,G4608,G6360);
  nand GNAME6453(G6453,G6700,G4637);
  nand GNAME6454(G6454,G6362,G4701);
  nand GNAME6455(G6455,G4637,G6360);
  or GNAME6456(G6456,G13899,G7123);
  nand GNAME6457(G6457,G6456,G4681);
  nand GNAME6458(G6458,G12610,G4683);
  nand GNAME6459(G6459,G4615,G6457);
  nand GNAME6460(G6460,G6360,G4730);
  nand GNAME6461(G6461,G12611,G4683);
  nand GNAME6462(G6462,G4607,G6457);
  nand GNAME6463(G6463,G6360,G4727);
  nand GNAME6464(G6464,G12563,G4683);
  nand GNAME6465(G6465,G4612,G6457);
  nand GNAME6466(G6466,G6360,G4724);
  nand GNAME6467(G6467,G12562,G4683);
  nand GNAME6468(G6468,G4611,G6457);
  nand GNAME6469(G6469,G6360,G4721);
  nand GNAME6470(G6470,G12612,G4683);
  nand GNAME6471(G6471,G4613,G6457);
  nand GNAME6472(G6472,G6360,G4718);
  nand GNAME6473(G6473,G12613,G4683);
  nand GNAME6474(G6474,G4609,G6457);
  nand GNAME6475(G6475,G6360,G4715);
  nand GNAME6476(G6476,G4683,G12560);
  nand GNAME6477(G6477,G4207,G6457);
  nand GNAME6478(G6478,G6360,G4571);
  nand GNAME6479(G6479,G4683,G12559);
  nand GNAME6480(G6480,G4209,G6457);
  nand GNAME6481(G6481,G6360,G4570);
  nand GNAME6482(G6482,G12561,G4683);
  nand GNAME6483(G6483,G4606,G6457);
  nand GNAME6484(G6484,G6360,G4712);
  nand GNAME6485(G6485,G12614,G4683);
  nand GNAME6486(G6486,G4618,G6457);
  nand GNAME6487(G6487,G6360,G4568);
  nand GNAME6488(G6488,G12615,G4683);
  nand GNAME6489(G6489,G4624,G6457);
  nand GNAME6490(G6490,G6360,G4567);
  nand GNAME6491(G6491,G12616,G4683);
  nand GNAME6492(G6492,G4623,G6457);
  nand GNAME6493(G6493,G6360,G4566);
  nand GNAME6494(G6494,G12617,G4683);
  nand GNAME6495(G6495,G4626,G6457);
  nand GNAME6496(G6496,G6360,G4565);
  nand GNAME6497(G6497,G12618,G4683);
  nand GNAME6498(G6498,G4619,G6457);
  nand GNAME6499(G6499,G6360,G4564);
  nand GNAME6500(G6500,G12619,G4683);
  nand GNAME6501(G6501,G4616,G6457);
  nand GNAME6502(G6502,G6360,G4563);
  nand GNAME6503(G6503,G12620,G4683);
  nand GNAME6504(G6504,G4620,G6457);
  nand GNAME6505(G6505,G6360,G4562);
  nand GNAME6506(G6506,G12621,G4683);
  nand GNAME6507(G6507,G4622,G6457);
  nand GNAME6508(G6508,G6360,G4561);
  nand GNAME6509(G6509,G12622,G4683);
  nand GNAME6510(G6510,G4617,G6457);
  nand GNAME6511(G6511,G6360,G4560);
  nand GNAME6512(G6512,G12623,G4683);
  nand GNAME6513(G6513,G4621,G6457);
  nand GNAME6514(G6514,G6360,G4559);
  nand GNAME6515(G6515,G12558,G4683);
  nand GNAME6516(G6516,G4610,G6457);
  nand GNAME6517(G6517,G6360,G4709);
  nand GNAME6518(G6518,G12625,G4683);
  nand GNAME6519(G6519,G4633,G6457);
  nand GNAME6520(G6520,G6360,G4759);
  nand GNAME6521(G6521,G12626,G4683);
  nand GNAME6522(G6522,G4634,G6457);
  nand GNAME6523(G6523,G6360,G4757);
  nand GNAME6524(G6524,G12627,G4683);
  nand GNAME6525(G6525,G4632,G6457);
  nand GNAME6526(G6526,G6360,G4754);
  nand GNAME6527(G6527,G12628,G4683);
  nand GNAME6528(G6528,G4630,G6457);
  nand GNAME6529(G6529,G6360,G4751);
  nand GNAME6530(G6530,G12629,G4683);
  nand GNAME6531(G6531,G4625,G6457);
  nand GNAME6532(G6532,G6360,G4748);
  nand GNAME6533(G6533,G12557,G4683);
  nand GNAME6534(G6534,G4628,G6457);
  nand GNAME6535(G6535,G6360,G4745);
  nand GNAME6536(G6536,G12630,G4683);
  nand GNAME6537(G6537,G4629,G6457);
  nand GNAME6538(G6538,G6360,G4742);
  nand GNAME6539(G6539,G12631,G4683);
  nand GNAME6540(G6540,G4631,G6457);
  nand GNAME6541(G6541,G6360,G4739);
  nand GNAME6542(G6542,G12556,G4683);
  nand GNAME6543(G6543,G4627,G6457);
  nand GNAME6544(G6544,G6360,G4736);
  nand GNAME6545(G6545,G12555,G4683);
  nand GNAME6546(G6546,G4614,G6457);
  nand GNAME6547(G6547,G6360,G4733);
  nand GNAME6548(G6548,G12624,G4683);
  nand GNAME6549(G6549,G4608,G6457);
  nand GNAME6550(G6550,G6360,G4706);
  nand GNAME6551(G6551,G12609,G4683);
  nand GNAME6552(G6552,G4637,G6457);
  nand GNAME6553(G6553,G6360,G4701);
  or GNAME6554(G6554,G4673,G4674);
  or GNAME6555(G6555,G4691,G4684);
  nand GNAME6556(G6556,G4615,G6555);
  nand GNAME6557(G6557,G6554,G4729);
  nand GNAME6558(G6558,G6124,G4730);
  nand GNAME6559(G6559,G36323,G4685);
  nand GNAME6560(G6560,G36355,G4686);
  nand GNAME6561(G6561,G4607,G6555);
  nand GNAME6562(G6562,G6554,G4726);
  nand GNAME6563(G6563,G6124,G4727);
  nand GNAME6564(G6564,G36322,G4685);
  nand GNAME6565(G6565,G36354,G4686);
  nand GNAME6566(G6566,G4612,G6555);
  nand GNAME6567(G6567,G6554,G4723);
  nand GNAME6568(G6568,G6124,G4724);
  nand GNAME6569(G6569,G36321,G4685);
  nand GNAME6570(G6570,G36353,G4686);
  nand GNAME6571(G6571,G4611,G6555);
  nand GNAME6572(G6572,G6554,G4720);
  nand GNAME6573(G6573,G6124,G4721);
  nand GNAME6574(G6574,G36320,G4685);
  nand GNAME6575(G6575,G36352,G4686);
  nand GNAME6576(G6576,G4613,G6555);
  nand GNAME6577(G6577,G6554,G4717);
  nand GNAME6578(G6578,G6124,G4718);
  nand GNAME6579(G6579,G36319,G4685);
  nand GNAME6580(G6580,G36351,G4686);
  nand GNAME6581(G6581,G4609,G6555);
  nand GNAME6582(G6582,G6554,G4714);
  nand GNAME6583(G6583,G6124,G4715);
  nand GNAME6584(G6584,G36318,G4685);
  nand GNAME6585(G6585,G36350,G4686);
  nand GNAME6586(G6586,G36333,G4685);
  nand GNAME6587(G6587,G36365,G4686);
  nand GNAME6588(G6588,G6156,G4567);
  nand GNAME6589(G6589,G4624,G4666);
  nand GNAME6590(G6590,G6155,G4568);
  nand GNAME6591(G6591,G4618,G4667);
  nand GNAME6592(G6592,G4207,G4691);
  nand GNAME6593(G6593,G4209,G4691);
  nand GNAME6594(G6594,G4606,G6555);
  nand GNAME6595(G6595,G6554,G4711);
  nand GNAME6596(G6596,G6124,G4712);
  nand GNAME6597(G6597,G36317,G4685);
  nand GNAME6598(G6598,G36349,G4686);
  nand GNAME6599(G6599,G4618,G4691);
  nand GNAME6600(G6600,G4624,G6555);
  nand GNAME6601(G6601,G6124,G4567);
  nand GNAME6602(G6602,G4623,G6555);
  nand GNAME6603(G6603,G6124,G4566);
  nand GNAME6604(G6604,G4626,G6555);
  nand GNAME6605(G6605,G6124,G4565);
  nand GNAME6606(G6606,G4619,G6555);
  nand GNAME6607(G6607,G6124,G4564);
  nand GNAME6608(G6608,G4616,G6555);
  nand GNAME6609(G6609,G6124,G4563);
  nand GNAME6610(G6610,G4620,G6555);
  nand GNAME6611(G6611,G6124,G4562);
  nand GNAME6612(G6612,G4622,G6555);
  nand GNAME6613(G6613,G6124,G4561);
  nand GNAME6614(G6614,G4617,G6555);
  nand GNAME6615(G6615,G6124,G4560);
  nand GNAME6616(G6616,G4621,G6555);
  nand GNAME6617(G6617,G6124,G4559);
  nand GNAME6618(G6618,G4610,G6555);
  nand GNAME6619(G6619,G6554,G4708);
  nand GNAME6620(G6620,G6124,G4709);
  nand GNAME6621(G6621,G36316,G4685);
  nand GNAME6622(G6622,G36348,G4686);
  nand GNAME6623(G6623,G4633,G6555);
  nand GNAME6624(G6624,G6554,G4697);
  nand GNAME6625(G6625,G6124,G4759);
  nand GNAME6626(G6626,G4634,G6555);
  nand GNAME6627(G6627,G6554,G4756);
  nand GNAME6628(G6628,G6124,G4757);
  nand GNAME6629(G6629,G36332,G4685);
  nand GNAME6630(G6630,G36364,G4686);
  nand GNAME6631(G6631,G4632,G6555);
  nand GNAME6632(G6632,G6554,G4753);
  nand GNAME6633(G6633,G6124,G4754);
  nand GNAME6634(G6634,G36331,G4685);
  nand GNAME6635(G6635,G36363,G4686);
  nand GNAME6636(G6636,G4630,G6555);
  nand GNAME6637(G6637,G6554,G4750);
  nand GNAME6638(G6638,G6124,G4751);
  nand GNAME6639(G6639,G36330,G4685);
  nand GNAME6640(G6640,G36362,G4686);
  nand GNAME6641(G6641,G4625,G6555);
  nand GNAME6642(G6642,G6554,G4747);
  nand GNAME6643(G6643,G6124,G4748);
  nand GNAME6644(G6644,G36329,G4685);
  nand GNAME6645(G6645,G36361,G4686);
  nand GNAME6646(G6646,G4628,G6555);
  nand GNAME6647(G6647,G6554,G4744);
  nand GNAME6648(G6648,G6124,G4745);
  nand GNAME6649(G6649,G36328,G4685);
  nand GNAME6650(G6650,G36360,G4686);
  nand GNAME6651(G6651,G4629,G6555);
  nand GNAME6652(G6652,G6554,G4741);
  nand GNAME6653(G6653,G6124,G4742);
  nand GNAME6654(G6654,G36327,G4685);
  nand GNAME6655(G6655,G36359,G4686);
  nand GNAME6656(G6656,G4631,G6555);
  nand GNAME6657(G6657,G6554,G4738);
  nand GNAME6658(G6658,G6124,G4739);
  nand GNAME6659(G6659,G36326,G4685);
  nand GNAME6660(G6660,G36358,G4686);
  nand GNAME6661(G6661,G4627,G6555);
  nand GNAME6662(G6662,G6554,G4735);
  nand GNAME6663(G6663,G6124,G4736);
  nand GNAME6664(G6664,G36325,G4685);
  nand GNAME6665(G6665,G36357,G4686);
  nand GNAME6666(G6666,G4614,G6555);
  nand GNAME6667(G6667,G6554,G4732);
  nand GNAME6668(G6668,G6124,G4733);
  nand GNAME6669(G6669,G36324,G4685);
  nand GNAME6670(G6670,G36356,G4686);
  nand GNAME6671(G6671,G4608,G6555);
  nand GNAME6672(G6672,G6554,G4705);
  nand GNAME6673(G6673,G6124,G4706);
  nand GNAME6674(G6674,G36315,G4685);
  nand GNAME6675(G6675,G36347,G4686);
  nand GNAME6676(G6676,G4637,G6555);
  nand GNAME6677(G6677,G6554,G4699);
  nand GNAME6678(G6678,G6124,G4701);
  nand GNAME6679(G6679,G36314,G4685);
  nand GNAME6680(G6680,G36346,G4686);
  nand GNAME6681(G6681,G4648,G4647);
  nand GNAME6682(G6682,G6719,G4591);
  nand GNAME6683(G6683,G4647,G4964);
  or GNAME6684(G6684,G4546,G4573,G4572);
  or GNAME6685(G6685,G4960,G4930,G4641,G4639,G4642);
  nand GNAME6686(G6686,G4972,G6682);
  nand GNAME6687(G6687,G6681,G4652);
  nand GNAME6688(G6688,G4973,G6683);
  nand GNAME6689(G6689,G4932,G36243);
  nand GNAME6690(G6690,G13842,G36249);
  nand GNAME6691(G6691,G4932,G36244);
  nand GNAME6692(G6692,G13811,G36249);
  nand GNAME6693(G6693,G6691,G6692);
  nand GNAME6694(G6694,G4932,G36242);
  nand GNAME6695(G6695,G13843,G36249);
  nand GNAME6696(G6696,G4542,G4689,G7124);
  or GNAME6697(G6697,G4542,G4690,G4541);
  nand GNAME6698(G6698,G4932,G36241);
  nand GNAME6699(G6699,G13810,G36249);
  not GNAME6700(G6700,G4691);
  nand GNAME6701(G6701,G4933,G36250);
  nand GNAME6702(G6702,G5083,G4966);
  nand GNAME6703(G6703,G4933,G36251);
  nand GNAME6704(G6704,G5084,G4966);
  nand GNAME6705(G6705,G4932,G36247,G36248);
  nand GNAME6706(G6706,G36249,G13813,G13840);
  nand GNAME6707(G6707,G6705,G6706);
  nand GNAME6708(G6708,G4932,G4537,G36248);
  nand GNAME6709(G6709,G36249,G4536,G13840);
  nand GNAME6710(G6710,G6708,G6709);
  nand GNAME6711(G6711,G4932,G4538,G36247);
  or GNAME6712(G6712,G4932,G13840,G4536);
  nand GNAME6713(G6713,G6711,G6712);
  or GNAME6714(G6714,G36249,G36248,G36247);
  or GNAME6715(G6715,G4932,G13813,G13840);
  nand GNAME6716(G6716,G6714,G6715);
  nand GNAME6717(G6717,G4932,G36246);
  nand GNAME6718(G6718,G13841,G36249);
  not GNAME6719(G6719,G4694);
  nand GNAME6720(G6720,G4932,G36239);
  nand GNAME6721(G6721,G13844,G36249);
  not GNAME6722(G6722,G4695);
  nand GNAME6723(G6723,G4932,G36240);
  nand GNAME6724(G6724,G13809,G36249);
  not GNAME6725(G6725,G4696);
  nand GNAME6726(G6726,G4932,G36237);
  nand GNAME6727(G6727,G13808,G36249);
  not GNAME6728(G6728,G4697);
  nand GNAME6729(G6729,G4932,G36238);
  nand GNAME6730(G6730,G13845,G36249);
  not GNAME6731(G6731,G4698);
  nand GNAME6732(G6732,G4932,G36218);
  nand GNAME6733(G6733,G36218,G36249);
  nand GNAME6734(G6734,G4932,G36245);
  nand GNAME6735(G6735,G13812,G36249);
  not GNAME6736(G6736,G4700);
  nand GNAME6737(G6737,G4959,G857);
  nand GNAME6738(G6738,G4699,G4934);
  nand GNAME6739(G6739,G6722,G4696);
  or GNAME6740(G6740,G4554,G4696);
  nand GNAME6741(G6741,G5081,G36250);
  nand GNAME6742(G6742,G4544,G5083);
  not GNAME6743(G6743,G4702);
  nand GNAME6744(G6744,G5081,G36251);
  nand GNAME6745(G6745,G4544,G5084);
  not GNAME6746(G6746,G4703);
  nand GNAME6747(G6747,G4935,G36282);
  nand GNAME6748(G6748,G5099,G4967);
  nand GNAME6749(G6749,G4932,G36219);
  nand GNAME6750(G6750,G13833,G36249);
  nand GNAME6751(G6751,G4959,G846);
  nand GNAME6752(G6752,G4934,G4705);
  nand GNAME6753(G6753,G4935,G36283);
  nand GNAME6754(G6754,G5113,G4967);
  nand GNAME6755(G6755,G4932,G36220);
  nand GNAME6756(G6756,G13814,G36249);
  nand GNAME6757(G6757,G4959,G835);
  nand GNAME6758(G6758,G4934,G4708);
  nand GNAME6759(G6759,G4935,G36284);
  nand GNAME6760(G6760,G5123,G4967);
  nand GNAME6761(G6761,G4932,G36221);
  nand GNAME6762(G6762,G13815,G36249);
  nand GNAME6763(G6763,G4959,G832);
  nand GNAME6764(G6764,G4934,G4711);
  nand GNAME6765(G6765,G4935,G36285);
  nand GNAME6766(G6766,G5133,G4967);
  nand GNAME6767(G6767,G4932,G36222);
  nand GNAME6768(G6768,G13838,G36249);
  nand GNAME6769(G6769,G4959,G831);
  nand GNAME6770(G6770,G4934,G4714);
  nand GNAME6771(G6771,G4935,G36286);
  nand GNAME6772(G6772,G5143,G4967);
  nand GNAME6773(G6773,G4932,G36223);
  nand GNAME6774(G6774,G13837,G36249);
  nand GNAME6775(G6775,G4959,G830);
  nand GNAME6776(G6776,G4934,G4717);
  nand GNAME6777(G6777,G4935,G36287);
  nand GNAME6778(G6778,G5153,G4967);
  nand GNAME6779(G6779,G4932,G36224);
  nand GNAME6780(G6780,G13816,G36249);
  nand GNAME6781(G6781,G4959,G829);
  nand GNAME6782(G6782,G4934,G4720);
  nand GNAME6783(G6783,G4935,G36288);
  nand GNAME6784(G6784,G5163,G4967);
  nand GNAME6785(G6785,G4932,G36225);
  nand GNAME6786(G6786,G13817,G36249);
  nand GNAME6787(G6787,G4959,G828);
  nand GNAME6788(G6788,G4934,G4723);
  nand GNAME6789(G6789,G4935,G36289);
  nand GNAME6790(G6790,G5173,G4967);
  nand GNAME6791(G6791,G4932,G36226);
  nand GNAME6792(G6792,G13836,G36249);
  nand GNAME6793(G6793,G4959,G827);
  nand GNAME6794(G6794,G4934,G4726);
  nand GNAME6795(G6795,G4935,G36290);
  nand GNAME6796(G6796,G5183,G4967);
  nand GNAME6797(G6797,G4932,G36227);
  nand GNAME6798(G6798,G13835,G36249);
  nand GNAME6799(G6799,G4959,G826);
  nand GNAME6800(G6800,G4934,G4729);
  nand GNAME6801(G6801,G4935,G36291);
  nand GNAME6802(G6802,G5193,G4967);
  nand GNAME6803(G6803,G4932,G36228);
  nand GNAME6804(G6804,G13803,G36249);
  nand GNAME6805(G6805,G4959,G856);
  nand GNAME6806(G6806,G4934,G4732);
  nand GNAME6807(G6807,G4935,G36292);
  nand GNAME6808(G6808,G5203,G4967);
  nand GNAME6809(G6809,G4932,G36229);
  nand GNAME6810(G6810,G13804,G36249);
  nand GNAME6811(G6811,G4959,G855);
  nand GNAME6812(G6812,G4934,G4735);
  nand GNAME6813(G6813,G4935,G36293);
  nand GNAME6814(G6814,G5213,G4967);
  nand GNAME6815(G6815,G4932,G36230);
  nand GNAME6816(G6816,G13850,G36249);
  nand GNAME6817(G6817,G4959,G854);
  nand GNAME6818(G6818,G4934,G4738);
  nand GNAME6819(G6819,G4935,G36294);
  nand GNAME6820(G6820,G5223,G4967);
  nand GNAME6821(G6821,G4932,G36231);
  nand GNAME6822(G6822,G13849,G36249);
  nand GNAME6823(G6823,G4959,G853);
  nand GNAME6824(G6824,G4934,G4741);
  nand GNAME6825(G6825,G4935,G36295);
  nand GNAME6826(G6826,G5233,G4967);
  nand GNAME6827(G6827,G4932,G36232);
  nand GNAME6828(G6828,G13805,G36249);
  nand GNAME6829(G6829,G4959,G852);
  nand GNAME6830(G6830,G4934,G4744);
  nand GNAME6831(G6831,G4935,G36296);
  nand GNAME6832(G6832,G5243,G4967);
  nand GNAME6833(G6833,G4932,G36233);
  nand GNAME6834(G6834,G13806,G36249);
  nand GNAME6835(G6835,G4959,G851);
  nand GNAME6836(G6836,G4934,G4747);
  nand GNAME6837(G6837,G4935,G36297);
  nand GNAME6838(G6838,G5253,G4967);
  nand GNAME6839(G6839,G4932,G36234);
  nand GNAME6840(G6840,G13848,G36249);
  nand GNAME6841(G6841,G4959,G850);
  nand GNAME6842(G6842,G4934,G4750);
  nand GNAME6843(G6843,G4935,G36298);
  nand GNAME6844(G6844,G5263,G4967);
  nand GNAME6845(G6845,G4932,G36235);
  nand GNAME6846(G6846,G13847,G36249);
  nand GNAME6847(G6847,G4959,G849);
  nand GNAME6848(G6848,G4934,G4753);
  nand GNAME6849(G6849,G4935,G36299);
  nand GNAME6850(G6850,G5273,G4967);
  nand GNAME6851(G6851,G4932,G36236);
  nand GNAME6852(G6852,G13807,G36249);
  nand GNAME6853(G6853,G4959,G848);
  nand GNAME6854(G6854,G4934,G4756);
  nand GNAME6855(G6855,G4935,G36300);
  nand GNAME6856(G6856,G5283,G4967);
  nand GNAME6857(G6857,G4959,G847);
  nand GNAME6858(G6858,G4697,G4934);
  nand GNAME6859(G6859,G4935,G36301);
  nand GNAME6860(G6860,G5293,G4967);
  nand GNAME6861(G6861,G4935,G36302);
  nand GNAME6862(G6862,G5303,G4967);
  nand GNAME6863(G6863,G4935,G36303);
  nand GNAME6864(G6864,G5313,G4967);
  nand GNAME6865(G6865,G4935,G36304);
  nand GNAME6866(G6866,G5323,G4967);
  nand GNAME6867(G6867,G4935,G36305);
  nand GNAME6868(G6868,G5333,G4967);
  nand GNAME6869(G6869,G4935,G36306);
  nand GNAME6870(G6870,G5343,G4967);
  nand GNAME6871(G6871,G4935,G36307);
  nand GNAME6872(G6872,G5353,G4967);
  nand GNAME6873(G6873,G4935,G36308);
  nand GNAME6874(G6874,G5363,G4967);
  nand GNAME6875(G6875,G4935,G36309);
  nand GNAME6876(G6876,G5373,G4967);
  nand GNAME6877(G6877,G4935,G36310);
  nand GNAME6878(G6878,G5383,G4967);
  nand GNAME6879(G6879,G4935,G36311);
  nand GNAME6880(G6880,G5396,G4967);
  nand GNAME6881(G6881,G4935,G36312);
  nand GNAME6882(G6882,G5402,G4967);
  nand GNAME6883(G6883,G4935,G36313);
  nand GNAME6884(G6884,G5405,G4967);
  nand GNAME6885(G6885,G4936,G36314);
  nand GNAME6886(G6886,G5099,G4968);
  nand GNAME6887(G6887,G4936,G36315);
  nand GNAME6888(G6888,G5113,G4968);
  nand GNAME6889(G6889,G4936,G36316);
  nand GNAME6890(G6890,G5123,G4968);
  nand GNAME6891(G6891,G4936,G36317);
  nand GNAME6892(G6892,G5133,G4968);
  nand GNAME6893(G6893,G4936,G36318);
  nand GNAME6894(G6894,G5143,G4968);
  nand GNAME6895(G6895,G4936,G36319);
  nand GNAME6896(G6896,G5153,G4968);
  nand GNAME6897(G6897,G4936,G36320);
  nand GNAME6898(G6898,G5163,G4968);
  nand GNAME6899(G6899,G4936,G36321);
  nand GNAME6900(G6900,G5173,G4968);
  nand GNAME6901(G6901,G4936,G36322);
  nand GNAME6902(G6902,G5183,G4968);
  nand GNAME6903(G6903,G4936,G36323);
  nand GNAME6904(G6904,G5193,G4968);
  nand GNAME6905(G6905,G4936,G36324);
  nand GNAME6906(G6906,G5203,G4968);
  nand GNAME6907(G6907,G4936,G36325);
  nand GNAME6908(G6908,G5213,G4968);
  nand GNAME6909(G6909,G4936,G36326);
  nand GNAME6910(G6910,G5223,G4968);
  nand GNAME6911(G6911,G4936,G36327);
  nand GNAME6912(G6912,G5233,G4968);
  nand GNAME6913(G6913,G4936,G36328);
  nand GNAME6914(G6914,G5243,G4968);
  nand GNAME6915(G6915,G4936,G36329);
  nand GNAME6916(G6916,G5253,G4968);
  nand GNAME6917(G6917,G4936,G36330);
  nand GNAME6918(G6918,G5263,G4968);
  nand GNAME6919(G6919,G4936,G36331);
  nand GNAME6920(G6920,G5273,G4968);
  nand GNAME6921(G6921,G4936,G36332);
  nand GNAME6922(G6922,G5283,G4968);
  nand GNAME6923(G6923,G4936,G36333);
  nand GNAME6924(G6924,G5293,G4968);
  nand GNAME6925(G6925,G4936,G36334);
  nand GNAME6926(G6926,G5303,G4968);
  nand GNAME6927(G6927,G4936,G36335);
  nand GNAME6928(G6928,G5313,G4968);
  nand GNAME6929(G6929,G4936,G36336);
  nand GNAME6930(G6930,G5323,G4968);
  nand GNAME6931(G6931,G4936,G36337);
  nand GNAME6932(G6932,G5333,G4968);
  nand GNAME6933(G6933,G4936,G36338);
  nand GNAME6934(G6934,G5343,G4968);
  nand GNAME6935(G6935,G4936,G36339);
  nand GNAME6936(G6936,G5353,G4968);
  nand GNAME6937(G6937,G4936,G36340);
  nand GNAME6938(G6938,G5363,G4968);
  nand GNAME6939(G6939,G4936,G36341);
  nand GNAME6940(G6940,G5373,G4968);
  nand GNAME6941(G6941,G4936,G36342);
  nand GNAME6942(G6942,G5383,G4968);
  nand GNAME6943(G6943,G4936,G36343);
  nand GNAME6944(G6944,G5396,G4968);
  nand GNAME6945(G6945,G4936,G36344);
  nand GNAME6946(G6946,G5402,G4968);
  nand GNAME6947(G6947,G4936,G36345);
  nand GNAME6948(G6948,G5405,G4968);
  nand GNAME6949(G6949,G4575,G36347);
  nand GNAME6950(G6950,G4969,G5418,G12624);
  nand GNAME6951(G6951,G4575,G36375);
  nand GNAME6952(G6952,G4969,G5391,G4547);
  nand GNAME6953(G6953,G4575,G36376);
  nand GNAME6954(G6954,G5618,G4969);
  nand GNAME6955(G6955,G4575,G36377);
  nand GNAME6956(G6956,G5621,G4969);
  nand GNAME6957(G6957,G4965,G36398);
  nand GNAME6958(G6958,G4637,G4591);
  nand GNAME6959(G6959,G4965,G36399);
  nand GNAME6960(G6960,G4608,G4591);
  nand GNAME6961(G6961,G4965,G36400);
  nand GNAME6962(G6962,G4610,G4591);
  nand GNAME6963(G6963,G4965,G36401);
  nand GNAME6964(G6964,G4606,G4591);
  nand GNAME6965(G6965,G4965,G36402);
  nand GNAME6966(G6966,G4609,G4591);
  nand GNAME6967(G6967,G4965,G36403);
  nand GNAME6968(G6968,G4613,G4591);
  nand GNAME6969(G6969,G4965,G36404);
  nand GNAME6970(G6970,G4611,G4591);
  nand GNAME6971(G6971,G4965,G36405);
  nand GNAME6972(G6972,G4612,G4591);
  nand GNAME6973(G6973,G4965,G36406);
  nand GNAME6974(G6974,G4607,G4591);
  nand GNAME6975(G6975,G4965,G36407);
  nand GNAME6976(G6976,G4615,G4591);
  nand GNAME6977(G6977,G4965,G36408);
  nand GNAME6978(G6978,G4614,G4591);
  nand GNAME6979(G6979,G4965,G36409);
  nand GNAME6980(G6980,G4627,G4591);
  nand GNAME6981(G6981,G4965,G36410);
  nand GNAME6982(G6982,G4631,G4591);
  nand GNAME6983(G6983,G4965,G36411);
  nand GNAME6984(G6984,G4629,G4591);
  nand GNAME6985(G6985,G4965,G36412);
  nand GNAME6986(G6986,G4628,G4591);
  nand GNAME6987(G6987,G4965,G36413);
  nand GNAME6988(G6988,G4625,G4591);
  nand GNAME6989(G6989,G4965,G36414);
  nand GNAME6990(G6990,G4630,G4591);
  nand GNAME6991(G6991,G4965,G36415);
  nand GNAME6992(G6992,G4632,G4591);
  nand GNAME6993(G6993,G4965,G36416);
  nand GNAME6994(G6994,G4634,G4591);
  nand GNAME6995(G6995,G4965,G36417);
  nand GNAME6996(G6996,G4633,G4591);
  nand GNAME6997(G6997,G4965,G36418);
  nand GNAME6998(G6998,G4621,G4591);
  nand GNAME6999(G6999,G4965,G36419);
  nand GNAME7000(G7000,G4617,G4591);
  nand GNAME7001(G7001,G4965,G36420);
  nand GNAME7002(G7002,G4622,G4591);
  nand GNAME7003(G7003,G4965,G36421);
  nand GNAME7004(G7004,G4620,G4591);
  nand GNAME7005(G7005,G4965,G36422);
  nand GNAME7006(G7006,G4616,G4591);
  nand GNAME7007(G7007,G4965,G36423);
  nand GNAME7008(G7008,G4619,G4591);
  nand GNAME7009(G7009,G4965,G36424);
  nand GNAME7010(G7010,G4626,G4591);
  nand GNAME7011(G7011,G4965,G36425);
  nand GNAME7012(G7012,G4623,G4591);
  nand GNAME7013(G7013,G4965,G36426);
  nand GNAME7014(G7014,G4624,G4591);
  nand GNAME7015(G7015,G4965,G36427);
  nand GNAME7016(G7016,G4618,G4591);
  nand GNAME7017(G7017,G4965,G36428);
  nand GNAME7018(G7018,G4209,G4591);
  nand GNAME7019(G7019,G4965,G36429);
  nand GNAME7020(G7020,G4207,G4591);
  nand GNAME7021(G7021,G4691,G4696);
  or GNAME7022(G7022,G4605,G4691);
  or GNAME7023(G7023,G4608,G4706);
  nand GNAME7024(G7024,G4608,G4706);
  nand GNAME7025(G7025,G7023,G7024);
  or GNAME7026(G7026,G4606,G4712);
  nand GNAME7027(G7027,G4606,G4712);
  nand GNAME7028(G7028,G7026,G7027);
  or GNAME7029(G7029,G4607,G4727);
  nand GNAME7030(G7030,G4607,G4727);
  nand GNAME7031(G7031,G7029,G7030);
  or GNAME7032(G7032,G4609,G4715);
  nand GNAME7033(G7033,G4609,G4715);
  nand GNAME7034(G7034,G7032,G7033);
  or GNAME7035(G7035,G4610,G4709);
  nand GNAME7036(G7036,G4610,G4709);
  nand GNAME7037(G7037,G7035,G7036);
  or GNAME7038(G7038,G4613,G4718);
  nand GNAME7039(G7039,G4613,G4718);
  nand GNAME7040(G7040,G7038,G7039);
  or GNAME7041(G7041,G4611,G4721);
  nand GNAME7042(G7042,G4611,G4721);
  nand GNAME7043(G7043,G7041,G7042);
  or GNAME7044(G7044,G4612,G4724);
  nand GNAME7045(G7045,G4612,G4724);
  nand GNAME7046(G7046,G7044,G7045);
  or GNAME7047(G7047,G4614,G4733);
  nand GNAME7048(G7048,G4614,G4733);
  nand GNAME7049(G7049,G7047,G7048);
  or GNAME7050(G7050,G4615,G4730);
  nand GNAME7051(G7051,G4615,G4730);
  nand GNAME7052(G7052,G7050,G7051);
  nand GNAME7053(G7053,G4617,G4560);
  or GNAME7054(G7054,G4560,G4617);
  nand GNAME7055(G7055,G7053,G7054);
  nand GNAME7056(G7056,G4616,G4563);
  or GNAME7057(G7057,G4563,G4616);
  nand GNAME7058(G7058,G7056,G7057);
  nand GNAME7059(G7059,G4209,G4570);
  or GNAME7060(G7060,G4209,G4570);
  nand GNAME7061(G7061,G7059,G7060);
  nand GNAME7062(G7062,G4620,G4562);
  or GNAME7063(G7063,G4562,G4620);
  nand GNAME7064(G7064,G7062,G7063);
  nand GNAME7065(G7065,G4618,G4568);
  or GNAME7066(G7066,G4568,G4618);
  nand GNAME7067(G7067,G7065,G7066);
  nand GNAME7068(G7068,G4619,G4564);
  or GNAME7069(G7069,G4564,G4619);
  nand GNAME7070(G7070,G7068,G7069);
  nand GNAME7071(G7071,G4623,G4566);
  or GNAME7072(G7072,G4566,G4623);
  nand GNAME7073(G7073,G7071,G7072);
  nand GNAME7074(G7074,G4621,G4559);
  or GNAME7075(G7075,G4559,G4621);
  nand GNAME7076(G7076,G7074,G7075);
  nand GNAME7077(G7077,G4622,G4561);
  or GNAME7078(G7078,G4561,G4622);
  nand GNAME7079(G7079,G7077,G7078);
  nand GNAME7080(G7080,G4207,G4571);
  or GNAME7081(G7081,G4207,G4571);
  nand GNAME7082(G7082,G7080,G7081);
  nand GNAME7083(G7083,G4624,G4567);
  or GNAME7084(G7084,G4567,G4624);
  nand GNAME7085(G7085,G7083,G7084);
  or GNAME7086(G7086,G4627,G4736);
  nand GNAME7087(G7087,G4627,G4736);
  nand GNAME7088(G7088,G7086,G7087);
  nand GNAME7089(G7089,G4626,G4565);
  or GNAME7090(G7090,G4565,G4626);
  nand GNAME7091(G7091,G7089,G7090);
  or GNAME7092(G7092,G4625,G4748);
  nand GNAME7093(G7093,G4625,G4748);
  nand GNAME7094(G7094,G7092,G7093);
  or GNAME7095(G7095,G4628,G4745);
  nand GNAME7096(G7096,G4628,G4745);
  nand GNAME7097(G7097,G7095,G7096);
  or GNAME7098(G7098,G4629,G4742);
  nand GNAME7099(G7099,G4629,G4742);
  nand GNAME7100(G7100,G7098,G7099);
  or GNAME7101(G7101,G4632,G4754);
  nand GNAME7102(G7102,G4632,G4754);
  nand GNAME7103(G7103,G7101,G7102);
  or GNAME7104(G7104,G4630,G4751);
  nand GNAME7105(G7105,G4630,G4751);
  nand GNAME7106(G7106,G7104,G7105);
  or GNAME7107(G7107,G4631,G4739);
  nand GNAME7108(G7108,G4631,G4739);
  nand GNAME7109(G7109,G7107,G7108);
  or GNAME7110(G7110,G4633,G4759);
  nand GNAME7111(G7111,G4633,G4759);
  nand GNAME7112(G7112,G7110,G7111);
  or GNAME7113(G7113,G4634,G4757);
  nand GNAME7114(G7114,G4634,G4757);
  nand GNAME7115(G7115,G7113,G7114);
  or GNAME7116(G7116,G4637,G4701);
  nand GNAME7117(G7117,G4637,G4701);
  nand GNAME7118(G7118,G7116,G7117);
  nand GNAME7119(G7119,G5813,G13005);
  nand GNAME7120(G7120,G4938,G5816);
  not GNAME7121(G7121,G4961);
  not GNAME7122(G7122,G4950);
  not GNAME7123(G7123,G4682);
  not GNAME7124(G7124,G4539);
  not GNAME7125(G7125,G4639);
  nand GNAME7126(G7126,G15015,G7568);
  or GNAME7127(G7127,G7758,G15014);
  nand GNAME7128(G7128,G7129,G7131,G7130);
  nand GNAME7129(G7129,G15014,G7758);
  or GNAME7130(G7130,G7566,G15013);
  nand GNAME7131(G7131,G7132,G7134,G7133);
  nand GNAME7132(G7132,G15013,G7566);
  or GNAME7133(G7133,G7761,G15012);
  nand GNAME7134(G7134,G9923,G9925,G9924);
  nand GNAME7135(G7135,G9108,G9109);
  nand GNAME7136(G7136,G9110,G9111);
  nand GNAME7137(G7137,G9112,G9113);
  nand GNAME7138(G7138,G9114,G9115);
  nand GNAME7139(G7139,G9116,G9117);
  nand GNAME7140(G7140,G9118,G9119);
  nand GNAME7141(G7141,G9120,G9121);
  nand GNAME7142(G7142,G9122,G9123);
  nand GNAME7143(G7143,G9124,G9125);
  nand GNAME7144(G7144,G9126,G9127);
  nand GNAME7145(G7145,G9092,G9093);
  nand GNAME7146(G7146,G9094,G9095);
  nand GNAME7147(G7147,G9096,G9097);
  nand GNAME7148(G7148,G9098,G9099);
  nand GNAME7149(G7149,G9100,G9101);
  nand GNAME7150(G7150,G9102,G9103);
  nand GNAME7151(G7151,G9104,G9105);
  nand GNAME7152(G7152,G9106,G9107);
  nand GNAME7153(G7153,G9128,G9129);
  nand GNAME7154(G7154,G9130,G9131);
  nand GNAME7155(G7155,G9537,G7611);
  nand GNAME7156(G7156,G9443,G9441,G9442);
  nand GNAME7157(G7157,G7876,G8337,G8338,G8339);
  nand GNAME7158(G7158,G9446,G9444,G9445);
  nand GNAME7159(G7159,G7876,G8329,G8330,G8331);
  nand GNAME7160(G7160,G9450,G9451,G9452,G7656);
  nand GNAME7161(G7161,G7876,G8321,G8322,G8323);
  nand GNAME7162(G7162,G9453,G9454,G9455,G7656);
  nand GNAME7163(G7163,G8312,G8313,G8314,G8315);
  nand GNAME7164(G7164,G9456,G9457,G9458,G7656);
  nand GNAME7165(G7165,G8303,G8304,G8305,G8306);
  nand GNAME7166(G7166,G9459,G9460,G9461,G7656);
  nand GNAME7167(G7167,G8294,G8295,G8296,G8297);
  nand GNAME7168(G7168,G9462,G9463,G9464,G7656);
  nand GNAME7169(G7169,G8285,G8286,G8287,G8288);
  nand GNAME7170(G7170,G9465,G9466,G9467,G7656);
  nand GNAME7171(G7171,G8276,G8277,G8278,G8279);
  nand GNAME7172(G7172,G9468,G9469,G9470,G7656);
  nand GNAME7173(G7173,G8267,G8268,G8269,G8270);
  nand GNAME7174(G7174,G9471,G9472,G9473,G7656);
  nand GNAME7175(G7175,G8258,G8259,G8260,G8261);
  nand GNAME7176(G7176,G9474,G9475,G9476,G7656);
  nand GNAME7177(G7177,G8249,G8250,G8251,G8252);
  nand GNAME7178(G7178,G9477,G9478,G9479,G7656);
  nand GNAME7179(G7179,G8238,G8239,G8240,G8241);
  nand GNAME7180(G7180,G9483,G9484,G9485,G7656);
  nand GNAME7181(G7181,G8226,G8227,G8228,G8229);
  nand GNAME7182(G7182,G9486,G9487,G9488,G7656);
  nand GNAME7183(G7183,G8214,G8215,G8216,G8217);
  nand GNAME7184(G7184,G9489,G9490,G9491,G7656);
  nand GNAME7185(G7185,G8202,G8203,G8204,G8205);
  nand GNAME7186(G7186,G9492,G9493,G9494,G7656);
  nand GNAME7187(G7187,G8190,G8191,G8192,G8193);
  nand GNAME7188(G7188,G9495,G9496,G9497,G7656);
  nand GNAME7189(G7189,G8178,G8179,G8180,G8181);
  nand GNAME7190(G7190,G9498,G9499,G9500,G7656);
  nand GNAME7191(G7191,G8166,G8167,G8168,G8169);
  nand GNAME7192(G7192,G9501,G9502,G9503,G7656);
  nand GNAME7193(G7193,G8154,G8155,G8156,G8157);
  nand GNAME7194(G7194,G9504,G9505,G9506,G7656);
  nand GNAME7195(G7195,G8142,G8143,G8144,G8145);
  nand GNAME7196(G7196,G9507,G9508,G9509,G7656);
  nand GNAME7197(G7197,G8130,G8131,G8132,G8133);
  nand GNAME7198(G7198,G9510,G9511,G9512,G7656);
  nand GNAME7199(G7199,G8118,G8119,G8120,G8121);
  nand GNAME7200(G7200,G9423,G9424,G9425,G7656);
  nand GNAME7201(G7201,G8106,G8107,G8108,G8109);
  nand GNAME7202(G7202,G9426,G9427,G9428,G7656);
  nand GNAME7203(G7203,G8094,G8095,G8096,G8097);
  nand GNAME7204(G7204,G9429,G9430,G9431,G7656);
  nand GNAME7205(G7205,G8082,G8083,G8084,G8085);
  nand GNAME7206(G7206,G9432,G9433,G9434,G7656);
  nand GNAME7207(G7207,G8070,G8071,G8072,G8073);
  nand GNAME7208(G7208,G9435,G9436,G9437,G7656);
  nand GNAME7209(G7209,G8058,G8059,G8060,G8061);
  nand GNAME7210(G7210,G9438,G9439,G9440,G7656);
  nand GNAME7211(G7211,G8046,G8047,G8048,G8049);
  nand GNAME7212(G7212,G9447,G9448,G9449,G7656);
  nand GNAME7213(G7213,G8034,G8035,G8036,G8037);
  nand GNAME7214(G7214,G9480,G9481,G9482,G7656);
  nand GNAME7215(G7215,G8016,G8017,G8018,G8019);
  nand GNAME7216(G7216,G9513,G9514,G9515,G7656);
  nand GNAME7217(G7217,G7984,G7985,G7986,G7987);
  nand GNAME7218(G7218,G9516,G9517,G9518,G7656);
  nand GNAME7219(G7219,G8021,G8022,G8023,G8024);
  nand GNAME7220(G7220,G9346,G9347);
  nand GNAME7221(G7221,G9348,G9349);
  nand GNAME7222(G7222,G9355,G9353,G9354);
  nand GNAME7223(G7223,G9358,G9356,G9357);
  nand GNAME7224(G7224,G9361,G9359,G9360);
  nand GNAME7225(G7225,G9364,G9362,G9363);
  nand GNAME7226(G7226,G9367,G9365,G9366);
  nand GNAME7227(G7227,G9370,G9368,G9369);
  nand GNAME7228(G7228,G9373,G9371,G9372);
  nand GNAME7229(G7229,G9376,G9374,G9375);
  nand GNAME7230(G7230,G9379,G9377,G9378);
  nand GNAME7231(G7231,G9382,G9380,G9381);
  nand GNAME7232(G7232,G9388,G9386,G9387);
  nand GNAME7233(G7233,G9391,G9389,G9390);
  nand GNAME7234(G7234,G9394,G9392,G9393);
  nand GNAME7235(G7235,G9397,G9395,G9396);
  nand GNAME7236(G7236,G9400,G9398,G9399);
  nand GNAME7237(G7237,G9403,G9401,G9402);
  nand GNAME7238(G7238,G9406,G9404,G9405);
  nand GNAME7239(G7239,G9409,G9407,G9408);
  nand GNAME7240(G7240,G9412,G9410,G9411);
  nand GNAME7241(G7241,G9415,G9413,G9414);
  nand GNAME7242(G7242,G9330,G9328,G9329);
  nand GNAME7243(G7243,G9333,G9331,G9332);
  nand GNAME7244(G7244,G9336,G9334,G9335);
  nand GNAME7245(G7245,G9339,G9337,G9338);
  nand GNAME7246(G7246,G9342,G9340,G9341);
  nand GNAME7247(G7247,G9345,G9343,G9344);
  nand GNAME7248(G7248,G9352,G9350,G9351);
  nand GNAME7249(G7249,G9385,G9383,G9384);
  nand GNAME7250(G7250,G9418,G9416,G9417);
  nand GNAME7251(G7251,G9419,G9420);
  or GNAME7252(G7252,G7535,G7642,G9323);
  or GNAME7253(G7253,G7254,G7659);
  nand GNAME7254(G7254,G9262,G9263,G9261,G7873,G9260);
  nand GNAME7255(G7255,G9268,G7873,G9267);
  nand GNAME7256(G7256,G9270,G7873,G9269);
  nand GNAME7257(G7257,G9272,G7873,G9271);
  nand GNAME7258(G7258,G9274,G7873,G9273);
  nand GNAME7259(G7259,G9276,G7873,G9275);
  nand GNAME7260(G7260,G9278,G7873,G9277);
  nand GNAME7261(G7261,G9280,G7873,G9279);
  nand GNAME7262(G7262,G9282,G7873,G9281);
  nand GNAME7263(G7263,G9284,G7873,G9283);
  nand GNAME7264(G7264,G9289,G7873,G9288);
  nand GNAME7265(G7265,G9292,G9290,G9291);
  nand GNAME7266(G7266,G9295,G9293,G9294);
  nand GNAME7267(G7267,G9298,G9296,G9297);
  nand GNAME7268(G7268,G9301,G9299,G9300);
  nand GNAME7269(G7269,G9304,G9302,G9303);
  nand GNAME7270(G7270,G9307,G9305,G9306);
  nand GNAME7271(G7271,G9310,G9308,G9309);
  nand GNAME7272(G7272,G9313,G9311,G9312);
  nand GNAME7273(G7273,G9316,G9314,G9315);
  nand GNAME7274(G7274,G9244,G9242,G9243);
  nand GNAME7275(G7275,G9247,G9245,G9246);
  nand GNAME7276(G7276,G9250,G9248,G9249);
  nand GNAME7277(G7277,G9253,G9251,G9252);
  nand GNAME7278(G7278,G9256,G9254,G9255);
  nand GNAME7279(G7279,G9259,G9257,G9258);
  nand GNAME7280(G7280,G9266,G9264,G9265);
  nand GNAME7281(G7281,G9287,G9285,G9286);
  nand GNAME7282(G7282,G9319,G9317,G9318);
  nand GNAME7283(G7283,G9322,G9320,G9321);
  nand GNAME7284(G7284,G9164,G7651);
  nand GNAME7285(G7285,G9165,G7651);
  nand GNAME7286(G7286,G9170,G7651);
  nand GNAME7287(G7287,G7650,G9172,G9173);
  nand GNAME7288(G7288,G7650,G9174,G9175);
  nand GNAME7289(G7289,G7650,G9176,G9177);
  nand GNAME7290(G7290,G7650,G9178,G9179);
  nand GNAME7291(G7291,G7650,G9180,G9181);
  nand GNAME7292(G7292,G7650,G9182,G9183);
  nand GNAME7293(G7293,G7650,G9184,G9185);
  nand GNAME7294(G7294,G7650,G9186,G9187);
  nand GNAME7295(G7295,G7650,G9188,G9189);
  nand GNAME7296(G7296,G7650,G9194,G9195);
  nand GNAME7297(G7297,G9196,G9197,G9198,G9199);
  nand GNAME7298(G7298,G9200,G9201,G9202,G9203);
  nand GNAME7299(G7299,G9204,G9205,G9206,G9207);
  nand GNAME7300(G7300,G9208,G9209,G9210,G9211);
  nand GNAME7301(G7301,G9212,G9213,G9214,G9215);
  nand GNAME7302(G7302,G9216,G9217,G9218,G9219);
  nand GNAME7303(G7303,G9220,G9221,G9222,G9223);
  nand GNAME7304(G7304,G9224,G9225,G9226,G9227);
  nand GNAME7305(G7305,G9228,G9229,G9230,G9231);
  nand GNAME7306(G7306,G9134,G9135,G9136,G9137);
  nand GNAME7307(G7307,G9138,G9139,G9140,G9141);
  nand GNAME7308(G7308,G9142,G9143,G9144,G9145);
  nand GNAME7309(G7309,G9146,G9147,G9148,G9149);
  nand GNAME7310(G7310,G9150,G9151,G9152,G9153);
  nand GNAME7311(G7311,G9154,G9155,G9156,G9157);
  nand GNAME7312(G7312,G9166,G9167,G9168,G9169);
  nand GNAME7313(G7313,G9190,G9191,G9192,G9193);
  nand GNAME7314(G7314,G9232,G9233,G9234,G9235);
  nand GNAME7315(G7315,G9236,G9237,G9238,G9239);
  nand GNAME7316(G7316,G36705,G8691);
  not GNAME7317(G7317,G36705);
  nand GNAME7318(G7318,G7887,G7885,G7886);
  nand GNAME7319(G7319,G7890,G7888,G7889);
  nand GNAME7320(G7320,G7893,G7891,G7892);
  nand GNAME7321(G7321,G7896,G7894,G7895);
  nand GNAME7322(G7322,G7899,G7897,G7898);
  nand GNAME7323(G7323,G7902,G7900,G7901);
  nand GNAME7324(G7324,G7905,G7903,G7904);
  nand GNAME7325(G7325,G7908,G7906,G7907);
  nand GNAME7326(G7326,G7911,G7909,G7910);
  nand GNAME7327(G7327,G7914,G7912,G7913);
  nand GNAME7328(G7328,G7917,G7915,G7916);
  nand GNAME7329(G7329,G7920,G7918,G7919);
  nand GNAME7330(G7330,G7923,G7921,G7922);
  nand GNAME7331(G7331,G7926,G7924,G7925);
  nand GNAME7332(G7332,G7929,G7927,G7928);
  nand GNAME7333(G7333,G7932,G7930,G7931);
  nand GNAME7334(G7334,G7935,G7933,G7934);
  nand GNAME7335(G7335,G7938,G7936,G7937);
  nand GNAME7336(G7336,G7941,G7939,G7940);
  nand GNAME7337(G7337,G7944,G7942,G7943);
  nand GNAME7338(G7338,G7947,G7945,G7946);
  nand GNAME7339(G7339,G7950,G7948,G7949);
  nand GNAME7340(G7340,G7953,G7951,G7952);
  nand GNAME7341(G7341,G7956,G7954,G7955);
  nand GNAME7342(G7342,G7959,G7957,G7958);
  nand GNAME7343(G7343,G7962,G7960,G7961);
  nand GNAME7344(G7344,G7965,G7963,G7964);
  nand GNAME7345(G7345,G7968,G7966,G7967);
  nand GNAME7346(G7346,G7971,G7969,G7970);
  nand GNAME7347(G7347,G7974,G7972,G7973);
  nand GNAME7348(G7348,G7977,G7975,G7976);
  nand GNAME7349(G7349,G7980,G7978,G7979);
  and GNAME7350(G7350,G7868,G36497);
  and GNAME7351(G7351,G7868,G36498);
  and GNAME7352(G7352,G7868,G36499);
  and GNAME7353(G7353,G7868,G36500);
  and GNAME7354(G7354,G7868,G36501);
  and GNAME7355(G7355,G7868,G36502);
  and GNAME7356(G7356,G7868,G36503);
  and GNAME7357(G7357,G7868,G36504);
  and GNAME7358(G7358,G7868,G36505);
  and GNAME7359(G7359,G7868,G36506);
  and GNAME7360(G7360,G7868,G36507);
  and GNAME7361(G7361,G7868,G36508);
  and GNAME7362(G7362,G7868,G36509);
  and GNAME7363(G7363,G7868,G36510);
  and GNAME7364(G7364,G7868,G36511);
  and GNAME7365(G7365,G7868,G36512);
  and GNAME7366(G7366,G7868,G36513);
  and GNAME7367(G7367,G7868,G36514);
  and GNAME7368(G7368,G7868,G36515);
  and GNAME7369(G7369,G7868,G36516);
  and GNAME7370(G7370,G7868,G36517);
  and GNAME7371(G7371,G7868,G36518);
  and GNAME7372(G7372,G7868,G36519);
  and GNAME7373(G7373,G7868,G36520);
  and GNAME7374(G7374,G7868,G36521);
  and GNAME7375(G7375,G7868,G36522);
  and GNAME7376(G7376,G7868,G36523);
  and GNAME7377(G7377,G7868,G36524);
  and GNAME7378(G7378,G7868,G36525);
  and GNAME7379(G7379,G7868,G36526);
  nand GNAME7380(G7380,G8012,G8013,G8014,G8015);
  nand GNAME7381(G7381,G8032,G8033,G8031,G8029,G8030);
  nand GNAME7382(G7382,G8044,G8045,G8043,G8041,G8042);
  nand GNAME7383(G7383,G8056,G8057,G8055,G8053,G8054);
  nand GNAME7384(G7384,G8068,G8069,G8067,G8065,G8066);
  nand GNAME7385(G7385,G8080,G8081,G8079,G8077,G8078);
  nand GNAME7386(G7386,G8092,G8093,G8091,G8089,G8090);
  nand GNAME7387(G7387,G8104,G8105,G8103,G8101,G8102);
  nand GNAME7388(G7388,G8116,G8117,G8115,G8113,G8114);
  nand GNAME7389(G7389,G8128,G8129,G8127,G8125,G8126);
  nand GNAME7390(G7390,G8140,G8141,G8139,G8137,G8138);
  nand GNAME7391(G7391,G8152,G8153,G8151,G8149,G8150);
  nand GNAME7392(G7392,G8164,G8165,G8163,G8161,G8162);
  nand GNAME7393(G7393,G8176,G8177,G8175,G8173,G8174);
  nand GNAME7394(G7394,G8188,G8189,G8187,G8185,G8186);
  nand GNAME7395(G7395,G8200,G8201,G8199,G8197,G8198);
  nand GNAME7396(G7396,G8212,G8213,G8211,G8209,G8210);
  nand GNAME7397(G7397,G8224,G8225,G8223,G8221,G8222);
  nand GNAME7398(G7398,G8236,G8237,G8235,G8233,G8234);
  nand GNAME7399(G7399,G8247,G8248,G8246,G8244,G8245);
  nand GNAME7400(G7400,G8256,G8257,G8255,G8253,G8254);
  nand GNAME7401(G7401,G8265,G8266,G8264,G8262,G8263);
  nand GNAME7402(G7402,G8274,G8275,G8273,G8271,G8272);
  nand GNAME7403(G7403,G8283,G8284,G8282,G8280,G8281);
  nand GNAME7404(G7404,G8292,G8293,G8291,G8289,G8290);
  nand GNAME7405(G7405,G8301,G8302,G8300,G8298,G8299);
  nand GNAME7406(G7406,G8310,G8311,G8309,G8307,G8308);
  nand GNAME7407(G7407,G8319,G8320,G8318,G8316,G8317);
  nand GNAME7408(G7408,G8327,G8328,G8326,G8324,G8325);
  nand GNAME7409(G7409,G8334,G8335,G8336,G9620,G9621);
  nand GNAME7410(G7410,G8341,G7874,G8340);
  nand GNAME7411(G7411,G8343,G7874,G8342);
  nand GNAME7412(G7412,G8349,G8350,G8351,G8352);
  nand GNAME7413(G7413,G8356,G8357,G8355,G8353,G8354);
  nand GNAME7414(G7414,G8361,G8362,G8360,G8358,G8359);
  nand GNAME7415(G7415,G8366,G8367,G8365,G8363,G8364);
  nand GNAME7416(G7416,G8371,G8372,G8370,G8368,G8369);
  nand GNAME7417(G7417,G8376,G8377,G8375,G8373,G8374);
  nand GNAME7418(G7418,G8381,G8382,G8380,G8378,G8379);
  nand GNAME7419(G7419,G8386,G8387,G8385,G8383,G8384);
  nand GNAME7420(G7420,G8391,G8392,G8390,G8388,G8389);
  nand GNAME7421(G7421,G8396,G8397,G8395,G8393,G8394);
  nand GNAME7422(G7422,G8401,G8402,G8400,G8398,G8399);
  nand GNAME7423(G7423,G8406,G8407,G8405,G8403,G8404);
  nand GNAME7424(G7424,G8411,G8412,G8410,G8408,G8409);
  nand GNAME7425(G7425,G8416,G8417,G8415,G8413,G8414);
  nand GNAME7426(G7426,G8421,G8422,G8420,G8418,G8419);
  nand GNAME7427(G7427,G8426,G8427,G8425,G8423,G8424);
  nand GNAME7428(G7428,G8431,G8432,G8430,G8428,G8429);
  nand GNAME7429(G7429,G8436,G8437,G8435,G8433,G8434);
  nand GNAME7430(G7430,G8441,G8442,G8440,G8438,G8439);
  nand GNAME7431(G7431,G8446,G8447,G8445,G8443,G8444);
  nand GNAME7432(G7432,G8451,G8452,G8450,G8448,G8449);
  nand GNAME7433(G7433,G8456,G8457,G8455,G8453,G8454);
  nand GNAME7434(G7434,G8461,G8462,G8460,G8458,G8459);
  nand GNAME7435(G7435,G8466,G8467,G8465,G8463,G8464);
  nand GNAME7436(G7436,G8471,G8472,G8470,G8468,G8469);
  nand GNAME7437(G7437,G8476,G8477,G8475,G8473,G8474);
  nand GNAME7438(G7438,G8481,G8482,G8480,G8478,G8479);
  nand GNAME7439(G7439,G8486,G8487,G8485,G8483,G8484);
  nand GNAME7440(G7440,G8491,G8492,G8490,G8488,G8489);
  nand GNAME7441(G7441,G8493,G8494,G8495,G9624,G9625);
  nand GNAME7442(G7442,G8497,G7875,G8496);
  nand GNAME7443(G7443,G8499,G7875,G8498);
  nand GNAME7444(G7444,G8511,G8512,G8510,G8508,G8509);
  nand GNAME7445(G7445,G8517,G7837,G8516,G8514,G8515);
  nand GNAME7446(G7446,G7781,G8523,G8521,G8522);
  nand GNAME7447(G7447,G7782,G8529,G8527,G8528);
  nand GNAME7448(G7448,G7783,G8532,G8533,G8534);
  nand GNAME7449(G7449,G7784,G8538,G8539,G8540);
  nand GNAME7450(G7450,G7785,G8544,G8545,G8546);
  nand GNAME7451(G7451,G7786,G8550,G8551,G8552);
  nand GNAME7452(G7452,G7787,G8556,G8557,G8558);
  nand GNAME7453(G7453,G7788,G8562,G8563,G8564);
  nand GNAME7454(G7454,G7789,G8568,G8569,G8570);
  nand GNAME7455(G7455,G7790,G8574,G8575,G8576);
  nand GNAME7456(G7456,G7791,G8580,G8581,G8582);
  nand GNAME7457(G7457,G7792,G8586,G8587,G8588);
  nand GNAME7458(G7458,G7793,G8592,G8593,G8594);
  nand GNAME7459(G7459,G7794,G8598,G8599,G8600);
  nand GNAME7460(G7460,G7795,G8604,G8605,G8606);
  nand GNAME7461(G7461,G7796,G8610,G8611,G8612);
  nand GNAME7462(G7462,G7797,G8616,G8617,G8618);
  nand GNAME7463(G7463,G7798,G8622,G8623,G8624);
  nand GNAME7464(G7464,G7799,G8628,G8629,G8630);
  nand GNAME7465(G7465,G7800,G8634,G8635,G8636);
  nand GNAME7466(G7466,G7801,G8640,G8641,G8642);
  nand GNAME7467(G7467,G7802,G8646,G8647,G8648);
  nand GNAME7468(G7468,G7803,G8652,G8653,G8654);
  nand GNAME7469(G7469,G7804,G8658,G8659,G8660);
  nand GNAME7470(G7470,G7805,G8664,G8665,G8666);
  nand GNAME7471(G7471,G7806,G8670,G8671,G8672);
  nand GNAME7472(G7472,G7807,G8676,G8677,G8678);
  nand GNAME7473(G7473,G8682,G7838,G8684,G8680,G8681);
  nand GNAME7474(G7474,G7602,G8685,G8686);
  nand GNAME7475(G7475,G7602,G8687,G8688);
  nand GNAME7476(G7476,G9028,G8696,G8695,G8693,G8694);
  nand GNAME7477(G7477,G8846,G8700,G8699,G8697,G8698);
  nand GNAME7478(G7478,G8941,G8704,G8703,G8701,G8702);
  nand GNAME7479(G7479,G8961,G8708,G8707,G8705,G8706);
  nand GNAME7480(G7480,G8815,G8712,G8711,G8709,G8710);
  nand GNAME7481(G7481,G9067,G8716,G8715,G8713,G8714);
  nand GNAME7482(G7482,G8885,G8720,G8719,G8717,G8718);
  nand GNAME7483(G7483,G8980,G8724,G8723,G8721,G8722);
  nand GNAME7484(G7484,G8866,G8728,G8727,G8725,G8726);
  nand GNAME7485(G7485,G9048,G8732,G8731,G8729,G8730);
  nand GNAME7486(G7486,G8912,G8736,G8735,G8733,G8734);
  nand GNAME7487(G7487,G9009,G8740,G8739,G8737,G8738);
  nand GNAME7488(G7488,G9086,G8744,G8743,G8741,G8742);
  nand GNAME7489(G7489,G8836,G8748,G8747,G8745,G8746);
  nand GNAME7490(G7490,G8951,G8752,G8751,G8749,G8750);
  nand GNAME7491(G7491,G8922,G8756,G8755,G8753,G8754);
  nand GNAME7492(G7492,G9038,G8760,G8759,G8757,G8758);
  nand GNAME7493(G7493,G8856,G8764,G8763,G8761,G8762);
  nand GNAME7494(G7494,G8999,G8768,G8767,G8765,G8766);
  nand GNAME7495(G7495,G8902,G8772,G8771,G8769,G8770);
  nand GNAME7496(G7496,G8791,G8789,G8790);
  nand GNAME7497(G7497,G7815,G8812,G8810,G8811);
  nand GNAME7498(G7498,G8825,G8826,G8824,G8822,G8823);
  nand GNAME7499(G7499,G7816,G8834,G8831,G8832);
  nand GNAME7500(G7500,G7817,G8843,G8841,G8844);
  nand GNAME7501(G7501,G7818,G8855,G8854,G8852);
  nand GNAME7502(G7502,G7819,G8864,G8861,G8862);
  nand GNAME7503(G7503,G8874,G8875,G8873,G8871,G8872);
  nand GNAME7504(G7504,G7820,G8883,G8880,G8881);
  nand GNAME7505(G7505,G8893,G8894,G8892,G8890,G8891);
  nand GNAME7506(G7506,G7821,G8899,G8897,G8898);
  nand GNAME7507(G7507,G7822,G8910,G8907,G8908);
  nand GNAME7508(G7508,G7823,G8920,G8917,G8918);
  nand GNAME7509(G7509,G8930,G8931,G8929,G8927,G8928);
  nand GNAME7510(G7510,G7824,G8938,G8936,G8939);
  nand GNAME7511(G7511,G7825,G8949,G8946,G8947);
  nand GNAME7512(G7512,G7826,G8958,G8956,G8959);
  nand GNAME7513(G7513,G8969,G8970,G8968,G8966,G8967);
  nand GNAME7514(G7514,G7827,G8978,G8975,G8976);
  nand GNAME7515(G7515,G8988,G8989,G8987,G8985,G8986);
  nand GNAME7516(G7516,G7828,G8998,G8997,G8995);
  nand GNAME7517(G7517,G7829,G9007,G9004,G9005);
  nand GNAME7518(G7518,G9017,G9018,G9016,G9014,G9015);
  nand GNAME7519(G7519,G7830,G9025,G9023,G9026);
  nand GNAME7520(G7520,G7831,G9037,G9036,G9034);
  nand GNAME7521(G7521,G7832,G9046,G9043,G9044);
  nand GNAME7522(G7522,G9056,G9057,G9055,G9053,G9054);
  nand GNAME7523(G7523,G7833,G9065,G9062,G9063);
  nand GNAME7524(G7524,G9075,G9076,G9074,G9072,G9073);
  nand GNAME7525(G7525,G7834,G9084,G9081,G9082);
  nor GNAME7526(G7526,G7317,G7527);
  and GNAME7527(G7527,G36705,G7533);
  not GNAME7528(G7528,G14405);
  not GNAME7529(G7529,G36491);
  not GNAME7530(G7530,G14377);
  not GNAME7531(G7531,G36492);
  not GNAME7532(G7532,G36493);
  not GNAME7533(G7533,G36494);
  nand GNAME7534(G7534,G9530,G7658);
  or GNAME7535(G7535,G7603,G7659);
  nand GNAME7536(G7536,G7657,G9530);
  not GNAME7537(G7537,G36675);
  nor GNAME7538(G7538,G7317,G7535);
  nand GNAME7539(G7539,G9530,G9533,G9534);
  and GNAME7540(G7540,G7840,G7990);
  and GNAME7541(G7541,G7667,G7668);
  nand GNAME7542(G7542,G9565,G7663,G9568);
  nor GNAME7543(G7543,G9562,G7663);
  nand GNAME7544(G7544,G7665,G7543);
  nand GNAME7545(G7545,G7540,G7541);
  and GNAME7546(G7546,G9574,G9571);
  nand GNAME7547(G7547,G7540,G7546);
  and GNAME7548(G7548,G14376,G36494);
  and GNAME7549(G7549,G7533,G36490);
  nand GNAME7550(G7550,G8008,G8009);
  and GNAME7551(G7551,G7663,G7664);
  and GNAME7552(G7552,G8011,G7551);
  nand GNAME7553(G7553,G7999,G7538);
  and GNAME7554(G7554,G7552,G7869);
  and GNAME7555(G7555,G7849,G7843);
  nand GNAME7556(G7556,G8006,G7555);
  and GNAME7557(G7557,G8007,G7869);
  nor GNAME7558(G7558,G7664,G9568);
  and GNAME7559(G7559,G9568,G7666);
  and GNAME7560(G7560,G9562,G7559);
  and GNAME7561(G7561,G9565,G9559);
  or GNAME7562(G7562,G7548,G7549);
  and GNAME7563(G7563,G8002,G7869);
  and GNAME7564(G7564,G8028,G7551);
  and GNAME7565(G7565,G7869,G7564);
  and GNAME7566(G7566,G7866,G813);
  and GNAME7567(G7567,G7866,G812);
  and GNAME7568(G7568,G7866,G811);
  and GNAME7569(G7569,G7866,G810);
  and GNAME7570(G7570,G7866,G809);
  and GNAME7571(G7571,G7866,G808);
  and GNAME7572(G7572,G7866,G807);
  and GNAME7573(G7573,G7866,G806);
  and GNAME7574(G7574,G7866,G805);
  and GNAME7575(G7575,G7866,G804);
  and GNAME7576(G7576,G8333,G7551);
  and GNAME7577(G7577,G7157,G7576);
  and GNAME7578(G7578,G7866,G802);
  and GNAME7579(G7579,G7866,G801);
  and GNAME7580(G7580,G7668,G9571);
  and GNAME7581(G7581,G7667,G9574);
  and GNAME7582(G7582,G7664,G7559);
  and GNAME7583(G7583,G7540,G7581);
  nand GNAME7584(G7584,G8348,G7538);
  and GNAME7585(G7585,G7552,G7870);
  and GNAME7586(G7586,G8007,G7870);
  and GNAME7587(G7587,G8002,G7870);
  and GNAME7588(G7588,G7564,G7870);
  nand GNAME7589(G7589,G9559,G7558);
  nand GNAME7590(G7590,G8504,G7538);
  and GNAME7591(G7591,G7552,G7871);
  and GNAME7592(G7592,G8507,G7871);
  or GNAME7593(G7593,G7666,G7589);
  nor GNAME7594(G7594,G7590,G7593);
  and GNAME7595(G7595,G9562,G9559);
  nand GNAME7596(G7596,G7666,G7558);
  nor GNAME7597(G7597,G8505,G7590);
  and GNAME7598(G7598,G7564,G7871);
  nor GNAME7599(G7599,G9568,G9565);
  and GNAME7600(G7600,G7665,G9565);
  and GNAME7601(G7601,G7619,G7851,G7850,G7847,G7620);
  and GNAME7602(G7602,G8683,G8684);
  nor GNAME7603(G7603,G7657,G7534);
  and GNAME7604(G7604,G9537,G7603);
  and GNAME7605(G7605,G36705,G7604);
  nor GNAME7606(G7606,G7670,G7867);
  and GNAME7607(G7607,G7542,G9562,G7593,G7601);
  nand GNAME7608(G7608,G7848,G7861);
  nor GNAME7609(G7609,G7610,G9922);
  nor GNAME7610(G7610,G7316,G7604);
  nor GNAME7611(G7611,G9562,G7542);
  and GNAME7612(G7612,G7611,G7670,G8003);
  not GNAME7613(G7613,G14239);
  and GNAME7614(G7614,G7659,G7664);
  and GNAME7615(G7615,G7811,G7812,G7810,G7808,G7809);
  and GNAME7616(G7616,G7813,G7814);
  and GNAME7617(G7617,G7615,G7616);
  and GNAME7618(G7618,G9559,G7842);
  nand GNAME7619(G7619,G7663,G7599);
  nand GNAME7620(G7620,G7663,G7600);
  and GNAME7621(G7621,G7608,G7538);
  and GNAME7622(G7622,G7865,G7621);
  nor GNAME7623(G7623,G9565,G7544);
  nor GNAME7624(G7624,G9922,G7593);
  and GNAME7625(G7625,G8802,G7538);
  and GNAME7626(G7626,G8028,G7864);
  and GNAME7627(G7627,G8011,G7864);
  nor GNAME7628(G7628,G7603,G7155,G7317);
  and GNAME7629(G7629,G8821,G7538);
  nand GNAME7630(G7630,G7867,G8808,G8809,G9519);
  nor GNAME7631(G7631,G8003,G7659);
  nor GNAME7632(G7632,G7659,G7562);
  nor GNAME7633(G7633,G7535,G9559,G9565);
  and GNAME7634(G7634,G7665,G7633);
  nor GNAME7635(G7635,G7603,G7663);
  and GNAME7636(G7636,G7600,G7635);
  and GNAME7637(G7637,G9568,G7633);
  and GNAME7638(G7638,G7599,G7635);
  nand GNAME7639(G7639,G7852,G7857,G7858,G7859);
  nand GNAME7640(G7640,G7877,G7878,G7879,G7880);
  nor GNAME7641(G7641,G7603,G7542);
  and GNAME7642(G7642,G9568,G7635);
  and GNAME7643(G7643,G7666,G7642);
  nor GNAME7644(G7644,G7603,G7620);
  and GNAME7645(G7645,G9565,G7642);
  nand GNAME7646(G7646,G7853,G7854,G7855,G7856);
  nand GNAME7647(G7647,G7881,G7882,G7883,G7884);
  and GNAME7648(G7648,G7603,G7631);
  and GNAME7649(G7649,G7603,G7632);
  and GNAME7650(G7650,G9158,G9159);
  and GNAME7651(G7651,G9163,G7650,G9162,G9160,G9161);
  and GNAME7652(G7652,G7847,G7596,G7846);
  nand GNAME7653(G7653,G7620,G7843,G9325);
  and GNAME7654(G7654,G7544,G7848,G7849,G7589);
  and GNAME7655(G7655,G7582,G791);
  and GNAME7656(G7656,G7659,G7652);
  and GNAME7657(G7657,G9526,G9527);
  nand GNAME7658(G7658,G9531,G9532);
  nand GNAME7659(G7659,G9535,G9536);
  nand GNAME7660(G7660,G9538,G9539);
  nand GNAME7661(G7661,G9540,G9541);
  nand GNAME7662(G7662,G9554,G9555);
  nand GNAME7663(G7663,G9557,G9558);
  nand GNAME7664(G7664,G9560,G9561);
  nand GNAME7665(G7665,G9566,G9567);
  nand GNAME7666(G7666,G9563,G9564);
  nand GNAME7667(G7667,G9569,G9570);
  nand GNAME7668(G7668,G9572,G9573);
  nand GNAME7669(G7669,G9575,G9576);
  nand GNAME7670(G7670,G9577,G9578);
  nand GNAME7671(G7671,G9584,G9585);
  nand GNAME7672(G7672,G9586,G9587);
  nand GNAME7673(G7673,G9588,G9589);
  nand GNAME7674(G7674,G9590,G9591);
  nand GNAME7675(G7675,G9592,G9593);
  nand GNAME7676(G7676,G9594,G9595);
  nand GNAME7677(G7677,G9596,G9597);
  nand GNAME7678(G7678,G9598,G9599);
  nand GNAME7679(G7679,G9600,G9601);
  nand GNAME7680(G7680,G9602,G9603);
  nand GNAME7681(G7681,G9604,G9605);
  nand GNAME7682(G7682,G9606,G9607);
  nand GNAME7683(G7683,G9608,G9609);
  nand GNAME7684(G7684,G9610,G9611);
  nand GNAME7685(G7685,G9612,G9613);
  nand GNAME7686(G7686,G9614,G9615);
  nand GNAME7687(G7687,G9616,G9617);
  nand GNAME7688(G7688,G9618,G9619);
  nand GNAME7689(G7689,G9632,G9633);
  nand GNAME7690(G7690,G9634,G9635);
  nand GNAME7691(G7691,G9636,G9637);
  nand GNAME7692(G7692,G9638,G9639);
  nand GNAME7693(G7693,G9640,G9641);
  nand GNAME7694(G7694,G9642,G9643);
  nand GNAME7695(G7695,G9644,G9645);
  nand GNAME7696(G7696,G9646,G9647);
  nand GNAME7697(G7697,G9648,G9649);
  nand GNAME7698(G7698,G9650,G9651);
  nand GNAME7699(G7699,G9652,G9653);
  nand GNAME7700(G7700,G9654,G9655);
  nand GNAME7701(G7701,G9656,G9657);
  nand GNAME7702(G7702,G9658,G9659);
  nand GNAME7703(G7703,G9660,G9661);
  nand GNAME7704(G7704,G9662,G9663);
  nand GNAME7705(G7705,G9664,G9665);
  nand GNAME7706(G7706,G9666,G9667);
  nand GNAME7707(G7707,G9668,G9669);
  nand GNAME7708(G7708,G9670,G9671);
  nand GNAME7709(G7709,G9672,G9673);
  nand GNAME7710(G7710,G9674,G9675);
  nand GNAME7711(G7711,G9676,G9677);
  nand GNAME7712(G7712,G9678,G9679);
  nand GNAME7713(G7713,G9680,G9681);
  nand GNAME7714(G7714,G9682,G9683);
  nand GNAME7715(G7715,G9684,G9685);
  nand GNAME7716(G7716,G9686,G9687);
  nand GNAME7717(G7717,G9688,G9689);
  nand GNAME7718(G7718,G9690,G9691);
  nand GNAME7719(G7719,G9692,G9693);
  nand GNAME7720(G7720,G9694,G9695);
  nand GNAME7721(G7721,G9848,G9849);
  nand GNAME7722(G7722,G9800,G9801);
  nand GNAME7723(G7723,G9791,G9792);
  nand GNAME7724(G7724,G9806,G9807);
  nand GNAME7725(G7725,G9812,G9813);
  nand GNAME7726(G7726,G9824,G9825);
  nand GNAME7727(G7727,G9830,G9831);
  nand GNAME7728(G7728,G9818,G9819);
  nand GNAME7729(G7729,G9836,G9837);
  nand GNAME7730(G7730,G9842,G9843);
  nand GNAME7731(G7731,G9704,G9705);
  nand GNAME7732(G7732,G9710,G9711);
  nand GNAME7733(G7733,G9698,G9699);
  nand GNAME7734(G7734,G9716,G9717);
  nand GNAME7735(G7735,G9722,G9723);
  nand GNAME7736(G7736,G9734,G9735);
  nand GNAME7737(G7737,G9740,G9741);
  nand GNAME7738(G7738,G9728,G9729);
  nand GNAME7739(G7739,G9746,G9747);
  nand GNAME7740(G7740,G9752,G9753);
  nand GNAME7741(G7741,G9858,G9859);
  nand GNAME7742(G7742,G9860,G9861);
  nand GNAME7743(G7743,G9862,G9863);
  nand GNAME7744(G7744,G9864,G9865);
  nand GNAME7745(G7745,G9866,G9867);
  nand GNAME7746(G7746,G9868,G9869);
  nand GNAME7747(G7747,G9870,G9871);
  nand GNAME7748(G7748,G9872,G9873);
  nand GNAME7749(G7749,G9874,G9875);
  nand GNAME7750(G7750,G9876,G9877);
  nand GNAME7751(G7751,G9878,G9879);
  nand GNAME7752(G7752,G9880,G9881);
  nand GNAME7753(G7753,G9882,G9883);
  nand GNAME7754(G7754,G9884,G9885);
  nand GNAME7755(G7755,G9886,G9887);
  nand GNAME7756(G7756,G9888,G9889);
  nand GNAME7757(G7757,G9890,G9891);
  nand GNAME7758(G7758,G9892,G9893);
  nand GNAME7759(G7759,G9894,G9895);
  nand GNAME7760(G7760,G9896,G9897);
  nand GNAME7761(G7761,G9898,G9899);
  nand GNAME7762(G7762,G9900,G9901);
  nand GNAME7763(G7763,G9902,G9903);
  nand GNAME7764(G7764,G9904,G9905);
  nand GNAME7765(G7765,G9906,G9907);
  nand GNAME7766(G7766,G9908,G9909);
  nand GNAME7767(G7767,G9910,G9911);
  nand GNAME7768(G7768,G9912,G9913);
  nand GNAME7769(G7769,G9914,G9915);
  nand GNAME7770(G7770,G9916,G9917);
  nand GNAME7771(G7771,G9918,G9919);
  nand GNAME7772(G7772,G9920,G9921);
  or GNAME7773(G7773,G36523,G36524,G36525,G36526);
  nor GNAME7774(G7774,G7773,G36522,G36521,G36520,G36519);
  or GNAME7775(G7775,G36515,G36516,G36517,G36518);
  nor GNAME7776(G7776,G7775,G36512,G36514,G36513);
  or GNAME7777(G7777,G36508,G36509,G36510,G36511);
  nor GNAME7778(G7778,G7777,G36505,G36507,G36506);
  or GNAME7779(G7779,G36501,G36502,G36503,G36504);
  nor GNAME7780(G7780,G7779,G36498,G36500,G36499);
  and GNAME7781(G7781,G8520,G8518,G8519);
  and GNAME7782(G7782,G8526,G8524,G8525);
  and GNAME7783(G7783,G8535,G8530,G8531);
  and GNAME7784(G7784,G8541,G8536,G8537);
  and GNAME7785(G7785,G8547,G8542,G8543);
  and GNAME7786(G7786,G8553,G8548,G8549);
  and GNAME7787(G7787,G8559,G8554,G8555);
  and GNAME7788(G7788,G8565,G8560,G8561);
  and GNAME7789(G7789,G8571,G8566,G8567);
  and GNAME7790(G7790,G8577,G8572,G8573);
  and GNAME7791(G7791,G8583,G8578,G8579);
  and GNAME7792(G7792,G8589,G8584,G8585);
  and GNAME7793(G7793,G8595,G8590,G8591);
  and GNAME7794(G7794,G8601,G8596,G8597);
  and GNAME7795(G7795,G8607,G8602,G8603);
  and GNAME7796(G7796,G8613,G8608,G8609);
  and GNAME7797(G7797,G8619,G8614,G8615);
  and GNAME7798(G7798,G8625,G8620,G8621);
  and GNAME7799(G7799,G8631,G8626,G8627);
  and GNAME7800(G7800,G8637,G8632,G8633);
  and GNAME7801(G7801,G8643,G8638,G8639);
  and GNAME7802(G7802,G8649,G8644,G8645);
  and GNAME7803(G7803,G8655,G8650,G8651);
  and GNAME7804(G7804,G8661,G8656,G8657);
  and GNAME7805(G7805,G8667,G8662,G8663);
  and GNAME7806(G7806,G8673,G8668,G8669);
  and GNAME7807(G7807,G8679,G8674,G8675);
  and GNAME7808(G7808,G9760,G9763,G9766);
  and GNAME7809(G7809,G9769,G9772,G9775);
  and GNAME7810(G7810,G9787,G9790,G9778,G9781,G9784);
  and GNAME7811(G7811,G9811,G9817,G9796,G9799,G9805);
  and GNAME7812(G7812,G9841,G9847,G9823,G9829,G9835);
  and GNAME7813(G7813,G9721,G9727,G9703,G9709,G9715);
  and GNAME7814(G7814,G9751,G9757,G9733,G9739,G9745);
  and GNAME7815(G7815,G8815,G8813,G8814);
  and GNAME7816(G7816,G8836,G8833,G8835);
  and GNAME7817(G7817,G8846,G8842,G8845);
  and GNAME7818(G7818,G8856,G8851,G8853);
  and GNAME7819(G7819,G8866,G8863,G8865);
  and GNAME7820(G7820,G8885,G8882,G8884);
  and GNAME7821(G7821,G8902,G8900,G8901);
  and GNAME7822(G7822,G8912,G8909,G8911);
  and GNAME7823(G7823,G8922,G8919,G8921);
  and GNAME7824(G7824,G8941,G8937,G8940);
  and GNAME7825(G7825,G8951,G8948,G8950);
  and GNAME7826(G7826,G8961,G8957,G8960);
  and GNAME7827(G7827,G8980,G8977,G8979);
  and GNAME7828(G7828,G8999,G8994,G8996);
  and GNAME7829(G7829,G9009,G9006,G9008);
  and GNAME7830(G7830,G9028,G9024,G9027);
  and GNAME7831(G7831,G9038,G9033,G9035);
  and GNAME7832(G7832,G9048,G9045,G9047);
  and GNAME7833(G7833,G9067,G9064,G9066);
  and GNAME7834(G7834,G9086,G9083,G9085);
  and GNAME7835(G7835,G7539,G7538);
  and GNAME7836(G7836,G7159,G7576);
  and GNAME7837(G7837,G9626,G9627);
  and GNAME7838(G7838,G9628,G9629);
  and GNAME7839(G7839,G9579,G8003);
  nand GNAME7840(G7840,G7989,G7981);
  nand GNAME7841(G7841,G7659,G8003);
  not GNAME7842(G7842,G7596);
  or GNAME7843(G7843,G7664,G7542);
  not GNAME7844(G7844,G7582);
  or GNAME7845(G7845,G7664,G7620);
  not GNAME7846(G7846,G7560);
  nand GNAME7847(G7847,G7664,G7599);
  nand GNAME7848(G7848,G9568,G7595);
  nand GNAME7849(G7849,G9568,G7543);
  nand GNAME7850(G7850,G7663,G7559);
  nand GNAME7851(G7851,G7664,G7600);
  nand GNAME7852(G7852,G7541,G7636);
  nand GNAME7853(G7853,G7541,G7645);
  nand GNAME7854(G7854,G7541,G7644);
  nand GNAME7855(G7855,G7541,G7641);
  nand GNAME7856(G7856,G7541,G7643);
  nand GNAME7857(G7857,G7541,G7634);
  nand GNAME7858(G7858,G7546,G7638);
  nand GNAME7859(G7859,G7541,G7637);
  nand GNAME7860(G7860,G9559,G7560);
  not GNAME7861(G7861,G7618);
  and GNAME7862(G7862,G9559,G7582);
  nand GNAME7863(G7863,G7616,G7615,G9853);
  not GNAME7864(G7864,G7547);
  not GNAME7865(G7865,G7545);
  not GNAME7866(G7866,G7839);
  not GNAME7867(G7867,G7605);
  not GNAME7868(G7868,G7835);
  not GNAME7869(G7869,G7553);
  not GNAME7870(G7870,G7584);
  not GNAME7871(G7871,G7590);
  nand GNAME7872(G7872,G7670,G36705,G7659);
  nand GNAME7873(G7873,G9240,G7665);
  nand GNAME7874(G7874,G7869,G7577);
  nand GNAME7875(G7875,G7577,G7870);
  nand GNAME7876(G7876,G9544,G14967);
  nand GNAME7877(G7877,G9521,G7634);
  nand GNAME7878(G7878,G9521,G7636);
  nand GNAME7879(G7879,G9521,G7637);
  nand GNAME7880(G7880,G9133,G7638);
  nand GNAME7881(G7881,G9521,G7641);
  nand GNAME7882(G7882,G9521,G7643);
  nand GNAME7883(G7883,G9521,G7644);
  nand GNAME7884(G7884,G9521,G7645);
  nand GNAME7885(G7885,G7317,G825);
  nand GNAME7886(G7886,G7526,G36463);
  nand GNAME7887(G7887,G7527,G36463);
  nand GNAME7888(G7888,G7317,G814);
  nand GNAME7889(G7889,G7526,G14397);
  nand GNAME7890(G7890,G7527,G36464);
  nand GNAME7891(G7891,G7317,G803);
  nand GNAME7892(G7892,G7526,G14378);
  nand GNAME7893(G7893,G7527,G36465);
  nand GNAME7894(G7894,G7317,G800);
  nand GNAME7895(G7895,G7526,G14379);
  nand GNAME7896(G7896,G7527,G36466);
  nand GNAME7897(G7897,G7317,G799);
  nand GNAME7898(G7898,G7526,G14402);
  nand GNAME7899(G7899,G7527,G36467);
  nand GNAME7900(G7900,G7317,G798);
  nand GNAME7901(G7901,G7526,G14401);
  nand GNAME7902(G7902,G7527,G36468);
  nand GNAME7903(G7903,G7317,G797);
  nand GNAME7904(G7904,G7526,G14380);
  nand GNAME7905(G7905,G7527,G36469);
  nand GNAME7906(G7906,G7317,G796);
  nand GNAME7907(G7907,G7526,G14381);
  nand GNAME7908(G7908,G7527,G36470);
  nand GNAME7909(G7909,G7317,G795);
  nand GNAME7910(G7910,G7526,G14400);
  nand GNAME7911(G7911,G7527,G36471);
  nand GNAME7912(G7912,G7317,G794);
  nand GNAME7913(G7913,G7526,G14399);
  nand GNAME7914(G7914,G7527,G36472);
  nand GNAME7915(G7915,G7317,G824);
  nand GNAME7916(G7916,G7526,G14367);
  nand GNAME7917(G7917,G7527,G36473);
  nand GNAME7918(G7918,G7317,G823);
  nand GNAME7919(G7919,G7526,G14368);
  nand GNAME7920(G7920,G7527,G36474);
  nand GNAME7921(G7921,G7317,G822);
  nand GNAME7922(G7922,G7526,G14414);
  nand GNAME7923(G7923,G7527,G36475);
  nand GNAME7924(G7924,G7317,G821);
  nand GNAME7925(G7925,G7526,G14413);
  nand GNAME7926(G7926,G7527,G36476);
  nand GNAME7927(G7927,G7317,G820);
  nand GNAME7928(G7928,G7526,G14369);
  nand GNAME7929(G7929,G7527,G36477);
  nand GNAME7930(G7930,G7317,G819);
  nand GNAME7931(G7931,G7526,G14370);
  nand GNAME7932(G7932,G7527,G36478);
  nand GNAME7933(G7933,G7317,G818);
  nand GNAME7934(G7934,G7526,G14412);
  nand GNAME7935(G7935,G7527,G36479);
  nand GNAME7936(G7936,G7317,G817);
  nand GNAME7937(G7937,G7526,G14411);
  nand GNAME7938(G7938,G7527,G36480);
  nand GNAME7939(G7939,G7317,G816);
  nand GNAME7940(G7940,G7526,G14371);
  nand GNAME7941(G7941,G7527,G36481);
  nand GNAME7942(G7942,G7317,G815);
  nand GNAME7943(G7943,G7526,G14372);
  nand GNAME7944(G7944,G7527,G36482);
  nand GNAME7945(G7945,G7317,G813);
  nand GNAME7946(G7946,G7526,G14409);
  nand GNAME7947(G7947,G7527,G36483);
  nand GNAME7948(G7948,G7317,G812);
  nand GNAME7949(G7949,G7526,G14408);
  nand GNAME7950(G7950,G7527,G36484);
  nand GNAME7951(G7951,G7317,G811);
  nand GNAME7952(G7952,G7526,G14373);
  nand GNAME7953(G7953,G7527,G36485);
  nand GNAME7954(G7954,G7317,G810);
  nand GNAME7955(G7955,G7526,G14374);
  nand GNAME7956(G7956,G7527,G36486);
  nand GNAME7957(G7957,G7317,G809);
  nand GNAME7958(G7958,G7526,G14407);
  nand GNAME7959(G7959,G7527,G36487);
  nand GNAME7960(G7960,G7317,G808);
  nand GNAME7961(G7961,G7526,G14406);
  nand GNAME7962(G7962,G7527,G36488);
  nand GNAME7963(G7963,G7317,G807);
  nand GNAME7964(G7964,G7526,G14375);
  nand GNAME7965(G7965,G7527,G36489);
  nand GNAME7966(G7966,G7317,G806);
  nand GNAME7967(G7967,G7526,G14376);
  nand GNAME7968(G7968,G7527,G36490);
  nand GNAME7969(G7969,G7317,G805);
  nand GNAME7970(G7970,G7526,G14405);
  nand GNAME7971(G7971,G7527,G36491);
  nand GNAME7972(G7972,G7317,G804);
  nand GNAME7973(G7973,G7526,G14377);
  nand GNAME7974(G7974,G7527,G36492);
  nand GNAME7975(G7975,G7317,G802);
  nand GNAME7976(G7976,G7526,G14404);
  nand GNAME7977(G7977,G7527,G36493);
  nand GNAME7978(G7978,G7317,G801);
  nand GNAME7979(G7979,G7526,G14398);
  nand GNAME7980(G7980,G7527,G36494);
  not GNAME7981(G7981,G7539);
  nand GNAME7982(G7982,G7536,G9531,G9532);
  nand GNAME7983(G7983,G7657,G7536);
  nand GNAME7984(G7984,G9544,G36695);
  nand GNAME7985(G7985,G9547,G36592);
  nand GNAME7986(G7986,G9550,G36560);
  nand GNAME7987(G7987,G9553,G36528);
  not GNAME7988(G7988,G7217);
  nand GNAME7989(G7989,G7774,G7776,G7778,G7780);
  nand GNAME7990(G7990,G36497,G7981);
  not GNAME7991(G7991,G7561);
  nand GNAME7992(G7992,G7664,G9565);
  nand GNAME7993(G7993,G7992,G7665);
  nand GNAME7994(G7994,G7993,G9559);
  nand GNAME7995(G7995,G7994,G9622);
  or GNAME7996(G7996,G7611,G7623);
  nand GNAME7997(G7997,G7996,G7865);
  nand GNAME7998(G7998,G7995,G7864);
  nand GNAME7999(G7999,G7997,G7998);
  not GNAME8000(G8000,G7559);
  nand GNAME8001(G8001,G9562,G7561);
  nand GNAME8002(G8002,G8001,G7589,G7860);
  not GNAME8003(G8003,G7562);
  nand GNAME8004(G8004,G7662,G7669);
  nand GNAME8005(G8005,G8004,G9848);
  or GNAME8006(G8006,G7595,G9565);
  or GNAME8007(G8007,G7600,G7556);
  nand GNAME8008(G8008,G14405,G7548);
  nand GNAME8009(G8009,G36491,G7549);
  not GNAME8010(G8010,G7550);
  nand GNAME8011(G8011,G9556,G8010);
  nand GNAME8012(G8012,G7217,G7554);
  nand GNAME8013(G8013,G7557,G14517);
  nand GNAME8014(G8014,G8005,G7563);
  nand GNAME8015(G8015,G7553,G36527);
  nand GNAME8016(G8016,G9553,G36529);
  nand GNAME8017(G8017,G9544,G36680);
  nand GNAME8018(G8018,G9547,G36593);
  nand GNAME8019(G8019,G9550,G36561);
  not GNAME8020(G8020,G7215);
  nand GNAME8021(G8021,G9544,G36685);
  nand GNAME8022(G8022,G9547,G36591);
  nand GNAME8023(G8023,G9550,G36559);
  nand GNAME8024(G8024,G9553,G36527);
  not GNAME8025(G8025,G7219);
  nand GNAME8026(G8026,G7662,G7671);
  nand GNAME8027(G8027,G8026,G9698);
  nand GNAME8028(G8028,G9580,G9581,G9582,G9583);
  nand GNAME8029(G8029,G7215,G7554);
  nand GNAME8030(G8030,G7219,G7565);
  nand GNAME8031(G8031,G7557,G14532);
  nand GNAME8032(G8032,G8027,G7563);
  nand GNAME8033(G8033,G7553,G36528);
  nand GNAME8034(G8034,G9553,G36530);
  nand GNAME8035(G8035,G9544,G14937);
  nand GNAME8036(G8036,G9547,G36594);
  nand GNAME8037(G8037,G9550,G36562);
  not GNAME8038(G8038,G7213);
  nand GNAME8039(G8039,G7662,G7672);
  nand GNAME8040(G8040,G8039,G9722);
  nand GNAME8041(G8041,G7213,G7554);
  nand GNAME8042(G8042,G7217,G7565);
  nand GNAME8043(G8043,G7557,G14466);
  nand GNAME8044(G8044,G8040,G7563);
  nand GNAME8045(G8045,G7553,G36529);
  nand GNAME8046(G8046,G9553,G36531);
  nand GNAME8047(G8047,G9544,G14941);
  nand GNAME8048(G8048,G9547,G36595);
  nand GNAME8049(G8049,G9550,G36563);
  not GNAME8050(G8050,G7211);
  nand GNAME8051(G8051,G7662,G7673);
  nand GNAME8052(G8052,G8051,G9704);
  nand GNAME8053(G8053,G7211,G7554);
  nand GNAME8054(G8054,G7215,G7565);
  nand GNAME8055(G8055,G7557,G14469);
  nand GNAME8056(G8056,G8052,G7563);
  nand GNAME8057(G8057,G7553,G36530);
  nand GNAME8058(G8058,G9553,G36532);
  nand GNAME8059(G8059,G9544,G14933);
  nand GNAME8060(G8060,G9547,G36596);
  nand GNAME8061(G8061,G9550,G36564);
  not GNAME8062(G8062,G7209);
  nand GNAME8063(G8063,G7662,G7674);
  nand GNAME8064(G8064,G8063,G9716);
  nand GNAME8065(G8065,G7209,G7554);
  nand GNAME8066(G8066,G7213,G7565);
  nand GNAME8067(G8067,G7557,G14521);
  nand GNAME8068(G8068,G8064,G7563);
  nand GNAME8069(G8069,G7553,G36531);
  nand GNAME8070(G8070,G9553,G36533);
  nand GNAME8071(G8071,G9544,G14919);
  nand GNAME8072(G8072,G9547,G36597);
  nand GNAME8073(G8073,G9550,G36565);
  not GNAME8074(G8074,G7207);
  nand GNAME8075(G8075,G7662,G7675);
  nand GNAME8076(G8076,G8075,G9728);
  nand GNAME8077(G8077,G7207,G7554);
  nand GNAME8078(G8078,G7211,G7565);
  nand GNAME8079(G8079,G7557,G14520);
  nand GNAME8080(G8080,G8076,G7563);
  nand GNAME8081(G8081,G7553,G36532);
  nand GNAME8082(G8082,G9553,G36534);
  nand GNAME8083(G8083,G9544,G14929);
  nand GNAME8084(G8084,G9547,G36598);
  nand GNAME8085(G8085,G9550,G36566);
  not GNAME8086(G8086,G7205);
  nand GNAME8087(G8087,G7662,G7676);
  nand GNAME8088(G8088,G8087,G9734);
  nand GNAME8089(G8089,G7205,G7554);
  nand GNAME8090(G8090,G7209,G7565);
  nand GNAME8091(G8091,G7557,G14470);
  nand GNAME8092(G8092,G8088,G7563);
  nand GNAME8093(G8093,G7553,G36533);
  nand GNAME8094(G8094,G9553,G36535);
  nand GNAME8095(G8095,G9544,G14923);
  nand GNAME8096(G8096,G9547,G36599);
  nand GNAME8097(G8097,G9550,G36567);
  not GNAME8098(G8098,G7203);
  nand GNAME8099(G8099,G7662,G7677);
  nand GNAME8100(G8100,G8099,G9740);
  nand GNAME8101(G8101,G7203,G7554);
  nand GNAME8102(G8102,G7207,G7565);
  nand GNAME8103(G8103,G7557,G14471);
  nand GNAME8104(G8104,G8100,G7563);
  nand GNAME8105(G8105,G7553,G36534);
  nand GNAME8106(G8106,G9553,G36536);
  nand GNAME8107(G8107,G9544,G14925);
  nand GNAME8108(G8108,G9547,G36600);
  nand GNAME8109(G8109,G9550,G36568);
  not GNAME8110(G8110,G7201);
  nand GNAME8111(G8111,G7662,G7678);
  nand GNAME8112(G8112,G8111,G9710);
  nand GNAME8113(G8113,G7201,G7554);
  nand GNAME8114(G8114,G7205,G7565);
  nand GNAME8115(G8115,G7557,G14519);
  nand GNAME8116(G8116,G8112,G7563);
  nand GNAME8117(G8117,G7553,G36535);
  nand GNAME8118(G8118,G9553,G36537);
  nand GNAME8119(G8119,G9544,G14924);
  nand GNAME8120(G8120,G9547,G36601);
  nand GNAME8121(G8121,G9550,G36569);
  not GNAME8122(G8122,G7199);
  nand GNAME8123(G8123,G7662,G7679);
  nand GNAME8124(G8124,G8123,G9752);
  nand GNAME8125(G8125,G7199,G7554);
  nand GNAME8126(G8126,G7203,G7565);
  nand GNAME8127(G8127,G7557,G14518);
  nand GNAME8128(G8128,G8124,G7563);
  nand GNAME8129(G8129,G7553,G36536);
  nand GNAME8130(G8130,G9553,G36538);
  nand GNAME8131(G8131,G9544,G14920);
  nand GNAME8132(G8132,G9547,G36602);
  nand GNAME8133(G8133,G9550,G36570);
  not GNAME8134(G8134,G7197);
  nand GNAME8135(G8135,G7662,G7680);
  nand GNAME8136(G8136,G8135,G9746);
  nand GNAME8137(G8137,G7197,G7554);
  nand GNAME8138(G8138,G7201,G7565);
  nand GNAME8139(G8139,G7557,G14463);
  nand GNAME8140(G8140,G8136,G7563);
  nand GNAME8141(G8141,G7553,G36537);
  nand GNAME8142(G8142,G9553,G36539);
  nand GNAME8143(G8143,G9544,G14935);
  nand GNAME8144(G8144,G9547,G36603);
  nand GNAME8145(G8145,G9550,G36571);
  not GNAME8146(G8146,G7195);
  nand GNAME8147(G8147,G7662,G7681);
  nand GNAME8148(G8148,G8147,G9791);
  nand GNAME8149(G8149,G7195,G7554);
  nand GNAME8150(G8150,G7199,G7565);
  nand GNAME8151(G8151,G7557,G14464);
  nand GNAME8152(G8152,G8148,G7563);
  nand GNAME8153(G8153,G7553,G36538);
  nand GNAME8154(G8154,G9553,G36540);
  nand GNAME8155(G8155,G9544,G14936);
  nand GNAME8156(G8156,G9547,G36604);
  nand GNAME8157(G8157,G9550,G36572);
  not GNAME8158(G8158,G7193);
  nand GNAME8159(G8159,G7662,G7682);
  nand GNAME8160(G8160,G8159,G9830);
  nand GNAME8161(G8161,G7193,G7554);
  nand GNAME8162(G8162,G7197,G7565);
  nand GNAME8163(G8163,G7557,G14539);
  nand GNAME8164(G8164,G8160,G7563);
  nand GNAME8165(G8165,G7553,G36539);
  nand GNAME8166(G8166,G9553,G36541);
  nand GNAME8167(G8167,G9544,G14942);
  nand GNAME8168(G8168,G9547,G36605);
  nand GNAME8169(G8169,G9550,G36573);
  not GNAME8170(G8170,G7191);
  nand GNAME8171(G8171,G7662,G7683);
  nand GNAME8172(G8172,G8171,G9812);
  nand GNAME8173(G8173,G7191,G7554);
  nand GNAME8174(G8174,G7195,G7565);
  nand GNAME8175(G8175,G7557,G14538);
  nand GNAME8176(G8176,G8172,G7563);
  nand GNAME8177(G8177,G7553,G36540);
  nand GNAME8178(G8178,G9553,G36542);
  nand GNAME8179(G8179,G9544,G14932);
  nand GNAME8180(G8180,G9547,G36606);
  nand GNAME8181(G8181,G9550,G36574);
  not GNAME8182(G8182,G7189);
  nand GNAME8183(G8183,G7662,G7684);
  nand GNAME8184(G8184,G8183,G9806);
  nand GNAME8185(G8185,G7189,G7554);
  nand GNAME8186(G8186,G7193,G7565);
  nand GNAME8187(G8187,G7557,G14465);
  nand GNAME8188(G8188,G8184,G7563);
  nand GNAME8189(G8189,G7553,G36541);
  nand GNAME8190(G8190,G9553,G36543);
  nand GNAME8191(G8191,G9544,G14918);
  nand GNAME8192(G8192,G9547,G36607);
  nand GNAME8193(G8193,G9550,G36575);
  not GNAME8194(G8194,G7187);
  nand GNAME8195(G8195,G7662,G7685);
  nand GNAME8196(G8196,G8195,G9800);
  nand GNAME8197(G8197,G7187,G7554);
  nand GNAME8198(G8198,G7191,G7565);
  nand GNAME8199(G8199,G7557,G14537);
  nand GNAME8200(G8200,G8196,G7563);
  nand GNAME8201(G8201,G7553,G36542);
  nand GNAME8202(G8202,G9553,G36544);
  nand GNAME8203(G8203,G9544,G14930);
  nand GNAME8204(G8204,G9547,G36608);
  nand GNAME8205(G8205,G9550,G36576);
  not GNAME8206(G8206,G7185);
  nand GNAME8207(G8207,G7662,G7686);
  nand GNAME8208(G8208,G8207,G9824);
  nand GNAME8209(G8209,G7185,G7554);
  nand GNAME8210(G8210,G7189,G7565);
  nand GNAME8211(G8211,G7557,G14536);
  nand GNAME8212(G8212,G8208,G7563);
  nand GNAME8213(G8213,G7553,G36543);
  nand GNAME8214(G8214,G9553,G36545);
  nand GNAME8215(G8215,G9544,G14922);
  nand GNAME8216(G8216,G9547,G36609);
  nand GNAME8217(G8217,G9550,G36577);
  not GNAME8218(G8218,G7183);
  nand GNAME8219(G8219,G7662,G7687);
  nand GNAME8220(G8220,G8219,G9818);
  nand GNAME8221(G8221,G7183,G7554);
  nand GNAME8222(G8222,G7187,G7565);
  nand GNAME8223(G8223,G7557,G14535);
  nand GNAME8224(G8224,G8220,G7563);
  nand GNAME8225(G8225,G7553,G36544);
  nand GNAME8226(G8226,G9553,G36546);
  nand GNAME8227(G8227,G9544,G14926);
  nand GNAME8228(G8228,G9547,G36610);
  nand GNAME8229(G8229,G9550,G36578);
  not GNAME8230(G8230,G7181);
  nand GNAME8231(G8231,G7662,G7688);
  nand GNAME8232(G8232,G8231,G9842);
  nand GNAME8233(G8233,G7181,G7554);
  nand GNAME8234(G8234,G7185,G7565);
  nand GNAME8235(G8235,G7557,G14534);
  nand GNAME8236(G8236,G8232,G7563);
  nand GNAME8237(G8237,G7553,G36545);
  nand GNAME8238(G8238,G9547,G36611);
  nand GNAME8239(G8239,G9550,G36579);
  nand GNAME8240(G8240,G9553,G36547);
  nand GNAME8241(G8241,G9544,G14931);
  nand GNAME8242(G8242,G7665,G7662);
  nand GNAME8243(G8243,G8242,G9836);
  nand GNAME8244(G8244,G7179,G7554);
  nand GNAME8245(G8245,G7183,G7565);
  nand GNAME8246(G8246,G7557,G14533);
  nand GNAME8247(G8247,G8243,G7563);
  nand GNAME8248(G8248,G7553,G36546);
  nand GNAME8249(G8249,G9547,G36612);
  nand GNAME8250(G8250,G9550,G36580);
  nand GNAME8251(G8251,G9553,G36548);
  nand GNAME8252(G8252,G9544,G14939);
  nand GNAME8253(G8253,G7177,G7554);
  nand GNAME8254(G8254,G7181,G7565);
  nand GNAME8255(G8255,G7557,G14531);
  nand GNAME8256(G8256,G7563,G7566);
  nand GNAME8257(G8257,G7553,G36547);
  nand GNAME8258(G8258,G9547,G36613);
  nand GNAME8259(G8259,G9550,G36581);
  nand GNAME8260(G8260,G9553,G36549);
  nand GNAME8261(G8261,G9544,G14928);
  nand GNAME8262(G8262,G7175,G7554);
  nand GNAME8263(G8263,G7179,G7565);
  nand GNAME8264(G8264,G7557,G14530);
  nand GNAME8265(G8265,G7563,G7567);
  nand GNAME8266(G8266,G7553,G36548);
  nand GNAME8267(G8267,G9547,G36614);
  nand GNAME8268(G8268,G9550,G36582);
  nand GNAME8269(G8269,G9553,G36550);
  nand GNAME8270(G8270,G9544,G14917);
  nand GNAME8271(G8271,G7173,G7554);
  nand GNAME8272(G8272,G7177,G7565);
  nand GNAME8273(G8273,G7557,G14529);
  nand GNAME8274(G8274,G7563,G7568);
  nand GNAME8275(G8275,G7553,G36549);
  nand GNAME8276(G8276,G9547,G36615);
  nand GNAME8277(G8277,G9550,G36583);
  nand GNAME8278(G8278,G9553,G36551);
  nand GNAME8279(G8279,G9544,G14921);
  nand GNAME8280(G8280,G7171,G7554);
  nand GNAME8281(G8281,G7175,G7565);
  nand GNAME8282(G8282,G7557,G14528);
  nand GNAME8283(G8283,G7563,G7569);
  nand GNAME8284(G8284,G7553,G36550);
  nand GNAME8285(G8285,G9547,G36616);
  nand GNAME8286(G8286,G9550,G36584);
  nand GNAME8287(G8287,G9553,G36552);
  nand GNAME8288(G8288,G9544,G14927);
  nand GNAME8289(G8289,G7169,G7554);
  nand GNAME8290(G8290,G7173,G7565);
  nand GNAME8291(G8291,G7557,G14527);
  nand GNAME8292(G8292,G7563,G7570);
  nand GNAME8293(G8293,G7553,G36551);
  nand GNAME8294(G8294,G9547,G36617);
  nand GNAME8295(G8295,G9550,G36585);
  nand GNAME8296(G8296,G9553,G36553);
  nand GNAME8297(G8297,G9544,G14938);
  nand GNAME8298(G8298,G7167,G7554);
  nand GNAME8299(G8299,G7171,G7565);
  nand GNAME8300(G8300,G7557,G14526);
  nand GNAME8301(G8301,G7563,G7571);
  nand GNAME8302(G8302,G7553,G36552);
  nand GNAME8303(G8303,G9547,G36618);
  nand GNAME8304(G8304,G9550,G36586);
  nand GNAME8305(G8305,G9553,G36554);
  nand GNAME8306(G8306,G9544,G14934);
  nand GNAME8307(G8307,G7165,G7554);
  nand GNAME8308(G8308,G7169,G7565);
  nand GNAME8309(G8309,G7557,G14525);
  nand GNAME8310(G8310,G7563,G7572);
  nand GNAME8311(G8311,G7553,G36553);
  nand GNAME8312(G8312,G9547,G36619);
  nand GNAME8313(G8313,G9550,G36587);
  nand GNAME8314(G8314,G9553,G36555);
  nand GNAME8315(G8315,G9544,G14940);
  nand GNAME8316(G8316,G7163,G7554);
  nand GNAME8317(G8317,G7167,G7565);
  nand GNAME8318(G8318,G7557,G14524);
  nand GNAME8319(G8319,G7563,G7573);
  nand GNAME8320(G8320,G7553,G36554);
  nand GNAME8321(G8321,G9547,G36620);
  nand GNAME8322(G8322,G9550,G36588);
  nand GNAME8323(G8323,G9553,G36556);
  nand GNAME8324(G8324,G7161,G7554);
  nand GNAME8325(G8325,G7165,G7565);
  nand GNAME8326(G8326,G7557,G14523);
  nand GNAME8327(G8327,G7563,G7574);
  nand GNAME8328(G8328,G7553,G36555);
  nand GNAME8329(G8329,G9547,G36621);
  nand GNAME8330(G8330,G9550,G36589);
  nand GNAME8331(G8331,G9553,G36557);
  nand GNAME8332(G8332,G7537,G7550);
  nand GNAME8333(G8333,G8332,G9556);
  nand GNAME8334(G8334,G7163,G7565);
  nand GNAME8335(G8335,G7557,G14522);
  nand GNAME8336(G8336,G7563,G7575);
  nand GNAME8337(G8337,G9547,G36622);
  nand GNAME8338(G8338,G9550,G36590);
  nand GNAME8339(G8339,G9553,G36558);
  nand GNAME8340(G8340,G7563,G7578);
  nand GNAME8341(G8341,G7553,G36557);
  nand GNAME8342(G8342,G7563,G7579);
  nand GNAME8343(G8343,G7553,G36558);
  nand GNAME8344(G8344,G7544,G9622,G9623);
  or GNAME8345(G8345,G7611,G7862);
  nand GNAME8346(G8346,G7580,G8344,G7540);
  nand GNAME8347(G8347,G8345,G7583);
  nand GNAME8348(G8348,G8346,G8347);
  nand GNAME8349(G8349,G7217,G7585);
  nand GNAME8350(G8350,G14517,G7586);
  nand GNAME8351(G8351,G8005,G7587);
  nand GNAME8352(G8352,G7584,G36559);
  nand GNAME8353(G8353,G7215,G7585);
  nand GNAME8354(G8354,G7219,G7588);
  nand GNAME8355(G8355,G14532,G7586);
  nand GNAME8356(G8356,G8027,G7587);
  nand GNAME8357(G8357,G7584,G36560);
  nand GNAME8358(G8358,G7213,G7585);
  nand GNAME8359(G8359,G7217,G7588);
  nand GNAME8360(G8360,G14466,G7586);
  nand GNAME8361(G8361,G8040,G7587);
  nand GNAME8362(G8362,G7584,G36561);
  nand GNAME8363(G8363,G7211,G7585);
  nand GNAME8364(G8364,G7215,G7588);
  nand GNAME8365(G8365,G14469,G7586);
  nand GNAME8366(G8366,G8052,G7587);
  nand GNAME8367(G8367,G7584,G36562);
  nand GNAME8368(G8368,G7209,G7585);
  nand GNAME8369(G8369,G7213,G7588);
  nand GNAME8370(G8370,G14521,G7586);
  nand GNAME8371(G8371,G8064,G7587);
  nand GNAME8372(G8372,G7584,G36563);
  nand GNAME8373(G8373,G7207,G7585);
  nand GNAME8374(G8374,G7211,G7588);
  nand GNAME8375(G8375,G14520,G7586);
  nand GNAME8376(G8376,G8076,G7587);
  nand GNAME8377(G8377,G7584,G36564);
  nand GNAME8378(G8378,G7205,G7585);
  nand GNAME8379(G8379,G7209,G7588);
  nand GNAME8380(G8380,G14470,G7586);
  nand GNAME8381(G8381,G8088,G7587);
  nand GNAME8382(G8382,G7584,G36565);
  nand GNAME8383(G8383,G7203,G7585);
  nand GNAME8384(G8384,G7207,G7588);
  nand GNAME8385(G8385,G14471,G7586);
  nand GNAME8386(G8386,G8100,G7587);
  nand GNAME8387(G8387,G7584,G36566);
  nand GNAME8388(G8388,G7201,G7585);
  nand GNAME8389(G8389,G7205,G7588);
  nand GNAME8390(G8390,G14519,G7586);
  nand GNAME8391(G8391,G8112,G7587);
  nand GNAME8392(G8392,G7584,G36567);
  nand GNAME8393(G8393,G7199,G7585);
  nand GNAME8394(G8394,G7203,G7588);
  nand GNAME8395(G8395,G14518,G7586);
  nand GNAME8396(G8396,G8124,G7587);
  nand GNAME8397(G8397,G7584,G36568);
  nand GNAME8398(G8398,G7197,G7585);
  nand GNAME8399(G8399,G7201,G7588);
  nand GNAME8400(G8400,G14463,G7586);
  nand GNAME8401(G8401,G8136,G7587);
  nand GNAME8402(G8402,G7584,G36569);
  nand GNAME8403(G8403,G7195,G7585);
  nand GNAME8404(G8404,G7199,G7588);
  nand GNAME8405(G8405,G14464,G7586);
  nand GNAME8406(G8406,G8148,G7587);
  nand GNAME8407(G8407,G7584,G36570);
  nand GNAME8408(G8408,G7193,G7585);
  nand GNAME8409(G8409,G7197,G7588);
  nand GNAME8410(G8410,G14539,G7586);
  nand GNAME8411(G8411,G8160,G7587);
  nand GNAME8412(G8412,G7584,G36571);
  nand GNAME8413(G8413,G7191,G7585);
  nand GNAME8414(G8414,G7195,G7588);
  nand GNAME8415(G8415,G14538,G7586);
  nand GNAME8416(G8416,G8172,G7587);
  nand GNAME8417(G8417,G7584,G36572);
  nand GNAME8418(G8418,G7189,G7585);
  nand GNAME8419(G8419,G7193,G7588);
  nand GNAME8420(G8420,G14465,G7586);
  nand GNAME8421(G8421,G8184,G7587);
  nand GNAME8422(G8422,G7584,G36573);
  nand GNAME8423(G8423,G7187,G7585);
  nand GNAME8424(G8424,G7191,G7588);
  nand GNAME8425(G8425,G14537,G7586);
  nand GNAME8426(G8426,G8196,G7587);
  nand GNAME8427(G8427,G7584,G36574);
  nand GNAME8428(G8428,G7185,G7585);
  nand GNAME8429(G8429,G7189,G7588);
  nand GNAME8430(G8430,G14536,G7586);
  nand GNAME8431(G8431,G8208,G7587);
  nand GNAME8432(G8432,G7584,G36575);
  nand GNAME8433(G8433,G7183,G7585);
  nand GNAME8434(G8434,G7187,G7588);
  nand GNAME8435(G8435,G14535,G7586);
  nand GNAME8436(G8436,G8220,G7587);
  nand GNAME8437(G8437,G7584,G36576);
  nand GNAME8438(G8438,G7181,G7585);
  nand GNAME8439(G8439,G7185,G7588);
  nand GNAME8440(G8440,G14534,G7586);
  nand GNAME8441(G8441,G8232,G7587);
  nand GNAME8442(G8442,G7584,G36577);
  nand GNAME8443(G8443,G7179,G7585);
  nand GNAME8444(G8444,G7183,G7588);
  nand GNAME8445(G8445,G14533,G7586);
  nand GNAME8446(G8446,G8243,G7587);
  nand GNAME8447(G8447,G7584,G36578);
  nand GNAME8448(G8448,G7177,G7585);
  nand GNAME8449(G8449,G7181,G7588);
  nand GNAME8450(G8450,G14531,G7586);
  nand GNAME8451(G8451,G7566,G7587);
  nand GNAME8452(G8452,G7584,G36579);
  nand GNAME8453(G8453,G7175,G7585);
  nand GNAME8454(G8454,G7179,G7588);
  nand GNAME8455(G8455,G14530,G7586);
  nand GNAME8456(G8456,G7567,G7587);
  nand GNAME8457(G8457,G7584,G36580);
  nand GNAME8458(G8458,G7173,G7585);
  nand GNAME8459(G8459,G7177,G7588);
  nand GNAME8460(G8460,G14529,G7586);
  nand GNAME8461(G8461,G7568,G7587);
  nand GNAME8462(G8462,G7584,G36581);
  nand GNAME8463(G8463,G7171,G7585);
  nand GNAME8464(G8464,G7175,G7588);
  nand GNAME8465(G8465,G14528,G7586);
  nand GNAME8466(G8466,G7569,G7587);
  nand GNAME8467(G8467,G7584,G36582);
  nand GNAME8468(G8468,G7169,G7585);
  nand GNAME8469(G8469,G7173,G7588);
  nand GNAME8470(G8470,G14527,G7586);
  nand GNAME8471(G8471,G7570,G7587);
  nand GNAME8472(G8472,G7584,G36583);
  nand GNAME8473(G8473,G7167,G7585);
  nand GNAME8474(G8474,G7171,G7588);
  nand GNAME8475(G8475,G14526,G7586);
  nand GNAME8476(G8476,G7571,G7587);
  nand GNAME8477(G8477,G7584,G36584);
  nand GNAME8478(G8478,G7165,G7585);
  nand GNAME8479(G8479,G7169,G7588);
  nand GNAME8480(G8480,G14525,G7586);
  nand GNAME8481(G8481,G7572,G7587);
  nand GNAME8482(G8482,G7584,G36585);
  nand GNAME8483(G8483,G7163,G7585);
  nand GNAME8484(G8484,G7167,G7588);
  nand GNAME8485(G8485,G14524,G7586);
  nand GNAME8486(G8486,G7573,G7587);
  nand GNAME8487(G8487,G7584,G36586);
  nand GNAME8488(G8488,G7161,G7585);
  nand GNAME8489(G8489,G7165,G7588);
  nand GNAME8490(G8490,G14523,G7586);
  nand GNAME8491(G8491,G7574,G7587);
  nand GNAME8492(G8492,G7584,G36587);
  nand GNAME8493(G8493,G7163,G7588);
  nand GNAME8494(G8494,G14522,G7586);
  nand GNAME8495(G8495,G7575,G7587);
  nand GNAME8496(G8496,G7578,G7587);
  nand GNAME8497(G8497,G7584,G36589);
  nand GNAME8498(G8498,G7579,G7587);
  nand GNAME8499(G8499,G7584,G36590);
  nand GNAME8500(G8500,G8000,G9559);
  nand GNAME8501(G8501,G8500,G7664);
  nand GNAME8502(G8502,G7580,G8345,G7540);
  nand GNAME8503(G8503,G8501,G7583);
  nand GNAME8504(G8504,G8503,G7593,G8502);
  not GNAME8505(G8505,G7608);
  nor GNAME8506(G8506,G7595,G9568);
  or GNAME8507(G8507,G8506,G7556);
  nand GNAME8508(G8508,G7217,G7591);
  nand GNAME8509(G8509,G14517,G7592);
  nand GNAME8510(G8510,G36685,G7594);
  nand GNAME8511(G8511,G8005,G7597);
  nand GNAME8512(G8512,G7590,G36591);
  nand GNAME8513(G8513,G7555,G7601);
  nand GNAME8514(G8514,G7215,G7591);
  nand GNAME8515(G8515,G7219,G7598);
  nand GNAME8516(G8516,G36695,G7594);
  nand GNAME8517(G8517,G8027,G7597);
  nand GNAME8518(G8518,G7213,G7591);
  nand GNAME8519(G8519,G7217,G7598);
  nand GNAME8520(G8520,G14466,G7592);
  nand GNAME8521(G8521,G36680,G7594);
  nand GNAME8522(G8522,G8040,G7597);
  nand GNAME8523(G8523,G7590,G36593);
  nand GNAME8524(G8524,G7211,G7591);
  nand GNAME8525(G8525,G7215,G7598);
  nand GNAME8526(G8526,G14469,G7592);
  nand GNAME8527(G8527,G14937,G7594);
  nand GNAME8528(G8528,G8052,G7597);
  nand GNAME8529(G8529,G7590,G36594);
  nand GNAME8530(G8530,G7209,G7591);
  nand GNAME8531(G8531,G7213,G7598);
  nand GNAME8532(G8532,G14521,G7592);
  nand GNAME8533(G8533,G14941,G7594);
  nand GNAME8534(G8534,G8064,G7597);
  nand GNAME8535(G8535,G7590,G36595);
  nand GNAME8536(G8536,G7207,G7591);
  nand GNAME8537(G8537,G7211,G7598);
  nand GNAME8538(G8538,G14520,G7592);
  nand GNAME8539(G8539,G14933,G7594);
  nand GNAME8540(G8540,G8076,G7597);
  nand GNAME8541(G8541,G7590,G36596);
  nand GNAME8542(G8542,G7205,G7591);
  nand GNAME8543(G8543,G7209,G7598);
  nand GNAME8544(G8544,G14470,G7592);
  nand GNAME8545(G8545,G14919,G7594);
  nand GNAME8546(G8546,G8088,G7597);
  nand GNAME8547(G8547,G7590,G36597);
  nand GNAME8548(G8548,G7203,G7591);
  nand GNAME8549(G8549,G7207,G7598);
  nand GNAME8550(G8550,G14471,G7592);
  nand GNAME8551(G8551,G14929,G7594);
  nand GNAME8552(G8552,G8100,G7597);
  nand GNAME8553(G8553,G7590,G36598);
  nand GNAME8554(G8554,G7201,G7591);
  nand GNAME8555(G8555,G7205,G7598);
  nand GNAME8556(G8556,G14519,G7592);
  nand GNAME8557(G8557,G14923,G7594);
  nand GNAME8558(G8558,G8112,G7597);
  nand GNAME8559(G8559,G7590,G36599);
  nand GNAME8560(G8560,G7199,G7591);
  nand GNAME8561(G8561,G7203,G7598);
  nand GNAME8562(G8562,G14518,G7592);
  nand GNAME8563(G8563,G14925,G7594);
  nand GNAME8564(G8564,G8124,G7597);
  nand GNAME8565(G8565,G7590,G36600);
  nand GNAME8566(G8566,G7197,G7591);
  nand GNAME8567(G8567,G7201,G7598);
  nand GNAME8568(G8568,G14463,G7592);
  nand GNAME8569(G8569,G14924,G7594);
  nand GNAME8570(G8570,G8136,G7597);
  nand GNAME8571(G8571,G7590,G36601);
  nand GNAME8572(G8572,G7195,G7591);
  nand GNAME8573(G8573,G7199,G7598);
  nand GNAME8574(G8574,G14464,G7592);
  nand GNAME8575(G8575,G14920,G7594);
  nand GNAME8576(G8576,G8148,G7597);
  nand GNAME8577(G8577,G7590,G36602);
  nand GNAME8578(G8578,G7193,G7591);
  nand GNAME8579(G8579,G7197,G7598);
  nand GNAME8580(G8580,G14539,G7592);
  nand GNAME8581(G8581,G14935,G7594);
  nand GNAME8582(G8582,G8160,G7597);
  nand GNAME8583(G8583,G7590,G36603);
  nand GNAME8584(G8584,G7191,G7591);
  nand GNAME8585(G8585,G7195,G7598);
  nand GNAME8586(G8586,G14538,G7592);
  nand GNAME8587(G8587,G14936,G7594);
  nand GNAME8588(G8588,G8172,G7597);
  nand GNAME8589(G8589,G7590,G36604);
  nand GNAME8590(G8590,G7189,G7591);
  nand GNAME8591(G8591,G7193,G7598);
  nand GNAME8592(G8592,G14465,G7592);
  nand GNAME8593(G8593,G14942,G7594);
  nand GNAME8594(G8594,G8184,G7597);
  nand GNAME8595(G8595,G7590,G36605);
  nand GNAME8596(G8596,G7187,G7591);
  nand GNAME8597(G8597,G7191,G7598);
  nand GNAME8598(G8598,G14537,G7592);
  nand GNAME8599(G8599,G14932,G7594);
  nand GNAME8600(G8600,G8196,G7597);
  nand GNAME8601(G8601,G7590,G36606);
  nand GNAME8602(G8602,G7185,G7591);
  nand GNAME8603(G8603,G7189,G7598);
  nand GNAME8604(G8604,G14536,G7592);
  nand GNAME8605(G8605,G14918,G7594);
  nand GNAME8606(G8606,G8208,G7597);
  nand GNAME8607(G8607,G7590,G36607);
  nand GNAME8608(G8608,G7183,G7591);
  nand GNAME8609(G8609,G7187,G7598);
  nand GNAME8610(G8610,G14535,G7592);
  nand GNAME8611(G8611,G14930,G7594);
  nand GNAME8612(G8612,G8220,G7597);
  nand GNAME8613(G8613,G7590,G36608);
  nand GNAME8614(G8614,G7181,G7591);
  nand GNAME8615(G8615,G7185,G7598);
  nand GNAME8616(G8616,G14534,G7592);
  nand GNAME8617(G8617,G14922,G7594);
  nand GNAME8618(G8618,G8232,G7597);
  nand GNAME8619(G8619,G7590,G36609);
  nand GNAME8620(G8620,G7179,G7591);
  nand GNAME8621(G8621,G7183,G7598);
  nand GNAME8622(G8622,G14533,G7592);
  nand GNAME8623(G8623,G14926,G7594);
  nand GNAME8624(G8624,G8243,G7597);
  nand GNAME8625(G8625,G7590,G36610);
  nand GNAME8626(G8626,G7177,G7591);
  nand GNAME8627(G8627,G7181,G7598);
  nand GNAME8628(G8628,G14531,G7592);
  nand GNAME8629(G8629,G14931,G7594);
  nand GNAME8630(G8630,G7566,G7597);
  nand GNAME8631(G8631,G7590,G36611);
  nand GNAME8632(G8632,G7175,G7591);
  nand GNAME8633(G8633,G7179,G7598);
  nand GNAME8634(G8634,G14530,G7592);
  nand GNAME8635(G8635,G14939,G7594);
  nand GNAME8636(G8636,G7567,G7597);
  nand GNAME8637(G8637,G7590,G36612);
  nand GNAME8638(G8638,G7173,G7591);
  nand GNAME8639(G8639,G7177,G7598);
  nand GNAME8640(G8640,G14529,G7592);
  nand GNAME8641(G8641,G14928,G7594);
  nand GNAME8642(G8642,G7568,G7597);
  nand GNAME8643(G8643,G7590,G36613);
  nand GNAME8644(G8644,G7171,G7591);
  nand GNAME8645(G8645,G7175,G7598);
  nand GNAME8646(G8646,G14528,G7592);
  nand GNAME8647(G8647,G14917,G7594);
  nand GNAME8648(G8648,G7569,G7597);
  nand GNAME8649(G8649,G7590,G36614);
  nand GNAME8650(G8650,G7169,G7591);
  nand GNAME8651(G8651,G7173,G7598);
  nand GNAME8652(G8652,G14527,G7592);
  nand GNAME8653(G8653,G14921,G7594);
  nand GNAME8654(G8654,G7570,G7597);
  nand GNAME8655(G8655,G7590,G36615);
  nand GNAME8656(G8656,G7167,G7591);
  nand GNAME8657(G8657,G7171,G7598);
  nand GNAME8658(G8658,G14526,G7592);
  nand GNAME8659(G8659,G14927,G7594);
  nand GNAME8660(G8660,G7571,G7597);
  nand GNAME8661(G8661,G7590,G36616);
  nand GNAME8662(G8662,G7165,G7591);
  nand GNAME8663(G8663,G7169,G7598);
  nand GNAME8664(G8664,G14525,G7592);
  nand GNAME8665(G8665,G14938,G7594);
  nand GNAME8666(G8666,G7572,G7597);
  nand GNAME8667(G8667,G7590,G36617);
  nand GNAME8668(G8668,G7163,G7591);
  nand GNAME8669(G8669,G7167,G7598);
  nand GNAME8670(G8670,G14524,G7592);
  nand GNAME8671(G8671,G14934,G7594);
  nand GNAME8672(G8672,G7573,G7597);
  nand GNAME8673(G8673,G7590,G36618);
  nand GNAME8674(G8674,G7161,G7591);
  nand GNAME8675(G8675,G7165,G7598);
  nand GNAME8676(G8676,G14523,G7592);
  nand GNAME8677(G8677,G14940,G7594);
  nand GNAME8678(G8678,G7574,G7597);
  nand GNAME8679(G8679,G7590,G36619);
  nand GNAME8680(G8680,G7163,G7598);
  nand GNAME8681(G8681,G14522,G7592);
  nand GNAME8682(G8682,G7575,G7597);
  nand GNAME8683(G8683,G7577,G7871);
  nand GNAME8684(G8684,G14967,G7594);
  nand GNAME8685(G8685,G7578,G7597);
  nand GNAME8686(G8686,G7590,G36621);
  nand GNAME8687(G8687,G7579,G7597);
  nand GNAME8688(G8688,G7590,G36622);
  or GNAME8689(G8689,G7551,G7535);
  nand GNAME8690(G8690,G8689,G9537);
  nand GNAME8691(G8691,G7866,G8690);
  nand GNAME8692(G8692,G7607,G8505);
  nand GNAME8693(G8693,G14533,G7606);
  nand GNAME8694(G8694,G9524,G14027);
  nand GNAME8695(G8695,G9523,G7665);
  nand GNAME8696(G8696,G7610,G36623);
  nand GNAME8697(G8697,G14534,G7606);
  nand GNAME8698(G8698,G9524,G14105);
  nand GNAME8699(G8699,G9523,G7688);
  nand GNAME8700(G8700,G7610,G36624);
  nand GNAME8701(G8701,G14535,G7606);
  nand GNAME8702(G8702,G9524,G14107);
  nand GNAME8703(G8703,G9523,G7687);
  nand GNAME8704(G8704,G7610,G36625);
  nand GNAME8705(G8705,G14536,G7606);
  nand GNAME8706(G8706,G9524,G14109);
  nand GNAME8707(G8707,G9523,G7686);
  nand GNAME8708(G8708,G7610,G36626);
  nand GNAME8709(G8709,G14537,G7606);
  nand GNAME8710(G8710,G9524,G14111);
  nand GNAME8711(G8711,G9523,G7685);
  nand GNAME8712(G8712,G7610,G36627);
  nand GNAME8713(G8713,G14465,G7606);
  nand GNAME8714(G8714,G9524,G14113);
  nand GNAME8715(G8715,G9523,G7684);
  nand GNAME8716(G8716,G7610,G36628);
  nand GNAME8717(G8717,G14538,G7606);
  nand GNAME8718(G8718,G9524,G14115);
  nand GNAME8719(G8719,G9523,G7683);
  nand GNAME8720(G8720,G7610,G36629);
  nand GNAME8721(G8721,G14539,G7606);
  nand GNAME8722(G8722,G9524,G14117);
  nand GNAME8723(G8723,G9523,G7682);
  nand GNAME8724(G8724,G7610,G36630);
  nand GNAME8725(G8725,G14464,G7606);
  nand GNAME8726(G8726,G9524,G14119);
  nand GNAME8727(G8727,G9523,G7681);
  nand GNAME8728(G8728,G7610,G36631);
  nand GNAME8729(G8729,G14463,G7606);
  nand GNAME8730(G8730,G9524,G14121);
  nand GNAME8731(G8731,G9523,G7680);
  nand GNAME8732(G8732,G7610,G36632);
  nand GNAME8733(G8733,G14518,G7606);
  nand GNAME8734(G8734,G9524,G14087);
  nand GNAME8735(G8735,G9523,G7679);
  nand GNAME8736(G8736,G7610,G36633);
  nand GNAME8737(G8737,G14519,G7606);
  nand GNAME8738(G8738,G9524,G14089);
  nand GNAME8739(G8739,G9523,G7678);
  nand GNAME8740(G8740,G7610,G36634);
  nand GNAME8741(G8741,G14471,G7606);
  nand GNAME8742(G8742,G9524,G14091);
  nand GNAME8743(G8743,G9523,G7677);
  nand GNAME8744(G8744,G7610,G36635);
  nand GNAME8745(G8745,G14470,G7606);
  nand GNAME8746(G8746,G9524,G14093);
  nand GNAME8747(G8747,G9523,G7676);
  nand GNAME8748(G8748,G7610,G36636);
  nand GNAME8749(G8749,G14520,G7606);
  nand GNAME8750(G8750,G9524,G14095);
  nand GNAME8751(G8751,G9523,G7675);
  nand GNAME8752(G8752,G7610,G36637);
  nand GNAME8753(G8753,G14521,G7606);
  nand GNAME8754(G8754,G9524,G14097);
  nand GNAME8755(G8755,G9523,G7674);
  nand GNAME8756(G8756,G7610,G36638);
  nand GNAME8757(G8757,G14469,G7606);
  nand GNAME8758(G8758,G9524,G14099);
  nand GNAME8759(G8759,G9523,G7673);
  nand GNAME8760(G8760,G7610,G36639);
  nand GNAME8761(G8761,G14466,G7606);
  nand GNAME8762(G8762,G9524,G14101);
  nand GNAME8763(G8763,G9523,G7672);
  nand GNAME8764(G8764,G7610,G36640);
  nand GNAME8765(G8765,G14532,G7606);
  nand GNAME8766(G8766,G9524,G14067);
  nand GNAME8767(G8767,G9523,G7671);
  nand GNAME8768(G8768,G7610,G36641);
  nand GNAME8769(G8769,G14517,G7606);
  nand GNAME8770(G8770,G9524,G14028);
  nand GNAME8771(G8771,G9523,G7669);
  nand GNAME8772(G8772,G7610,G36642);
  nand GNAME8773(G8773,G9853,G7617);
  nand GNAME8774(G8774,G7863,G7618);
  or GNAME8775(G8775,G14993,G7619);
  nand GNAME8776(G8776,G9696,G9697,G8774,G8775);
  nand GNAME8777(G8777,G7616,G7543,G7615);
  nand GNAME8778(G8778,G7595,G7617);
  nand GNAME8779(G8779,G8777,G8778);
  nand GNAME8780(G8780,G14993,G7663,G9562);
  nand GNAME8781(G8781,G8779,G9853);
  nand GNAME8782(G8782,G7551,G14239);
  nand GNAME8783(G8783,G8773,G9559,G7599,G7614);
  nand GNAME8784(G8784,G9856,G9857,G7659,G9568);
  nand GNAME8785(G8785,G8776,G7659);
  nand GNAME8786(G8786,G8785,G8783,G8784);
  nor GNAME8787(G8787,G7612,G7659);
  or GNAME8788(G8788,G7317,G7604,G7614,G8787);
  nand GNAME8789(G8789,G14239,G7538,G7612);
  nand GNAME8790(G8790,G8788,G36675);
  nand GNAME8791(G8791,G36705,G8786);
  nand GNAME8792(G8792,G7191,G7626);
  nand GNAME8793(G8793,G7187,G7627);
  nand GNAME8794(G8794,G7547,G14932);
  nand GNAME8795(G8795,G8794,G8792,G8793);
  nand GNAME8796(G8796,G7846,G7596);
  nand GNAME8797(G8797,G8796,G7663);
  or GNAME8798(G8798,G7666,G7544);
  nand GNAME8799(G8799,G7845,G8797,G8798,G7555);
  nand GNAME8800(G8800,G8799,G7865);
  nand GNAME8801(G8801,G7864,G7623);
  nand GNAME8802(G8802,G8800,G8801);
  nand GNAME8803(G8803,G9568,G9565);
  nand GNAME8804(G8804,G8803,G7551);
  nand GNAME8805(G8805,G7545,G8799);
  nand GNAME8806(G8806,G7547,G7623);
  nand GNAME8807(G8807,G8806,G8804,G8805);
  nand GNAME8808(G8808,G8807,G7538);
  nand GNAME8809(G8809,G36705,G7659);
  nand GNAME8810(G8810,G8196,G7622);
  nand GNAME8811(G8811,G7630,G14932);
  nand GNAME8812(G8812,G7722,G7624);
  nand GNAME8813(G8813,G14537,G7625);
  nand GNAME8814(G8814,G8795,G7628);
  nand GNAME8815(G8815,G7317,G36676);
  nand GNAME8816(G8816,G7169,G7626);
  nand GNAME8817(G8817,G7165,G7627);
  nand GNAME8818(G8818,G7547,G14938);
  nand GNAME8819(G8819,G8818,G8816,G8817);
  nand GNAME8820(G8820,G7608,G7865);
  nand GNAME8821(G8821,G8820,G7593);
  nand GNAME8822(G8822,G7572,G7629);
  nand GNAME8823(G8823,G14525,G7625);
  nand GNAME8824(G8824,G7630,G14938);
  nand GNAME8825(G8825,G8819,G7628);
  nand GNAME8826(G8826,G7317,G36677);
  nand GNAME8827(G8827,G7209,G7626);
  nand GNAME8828(G8828,G7205,G7627);
  nand GNAME8829(G8829,G7547,G14919);
  nand GNAME8830(G8830,G8829,G8827,G8828);
  nand GNAME8831(G8831,G8088,G7622);
  nand GNAME8832(G8832,G7630,G14919);
  nand GNAME8833(G8833,G7736,G7624);
  nand GNAME8834(G8834,G14470,G7625);
  nand GNAME8835(G8835,G8830,G7628);
  nand GNAME8836(G8836,G7317,G36678);
  nand GNAME8837(G8837,G7185,G7626);
  nand GNAME8838(G8838,G7181,G7627);
  nand GNAME8839(G8839,G7547,G14922);
  nand GNAME8840(G8840,G8839,G8837,G8838);
  nand GNAME8841(G8841,G8232,G7622);
  nand GNAME8842(G8842,G7630,G14922);
  nand GNAME8843(G8843,G7730,G7624);
  nand GNAME8844(G8844,G14534,G7625);
  nand GNAME8845(G8845,G8840,G7628);
  nand GNAME8846(G8846,G7317,G36679);
  nand GNAME8847(G8847,G7217,G7626);
  nand GNAME8848(G8848,G7213,G7627);
  nand GNAME8849(G8849,G7547,G36680);
  nand GNAME8850(G8850,G8849,G8847,G8848);
  nand GNAME8851(G8851,G8040,G7622);
  nand GNAME8852(G8852,G7630,G36680);
  nand GNAME8853(G8853,G7735,G7624);
  nand GNAME8854(G8854,G14466,G7625);
  nand GNAME8855(G8855,G8850,G7628);
  nand GNAME8856(G8856,G7317,G36680);
  nand GNAME8857(G8857,G7199,G7626);
  nand GNAME8858(G8858,G7195,G7627);
  nand GNAME8859(G8859,G7547,G14920);
  nand GNAME8860(G8860,G8859,G8857,G8858);
  nand GNAME8861(G8861,G8148,G7622);
  nand GNAME8862(G8862,G7630,G14920);
  nand GNAME8863(G8863,G7723,G7624);
  nand GNAME8864(G8864,G14464,G7625);
  nand GNAME8865(G8865,G8860,G7628);
  nand GNAME8866(G8866,G7317,G36681);
  nand GNAME8867(G8867,G7177,G7626);
  nand GNAME8868(G8868,G7173,G7627);
  nand GNAME8869(G8869,G7547,G14928);
  nand GNAME8870(G8870,G8869,G8867,G8868);
  nand GNAME8871(G8871,G7568,G7629);
  nand GNAME8872(G8872,G14529,G7625);
  nand GNAME8873(G8873,G7630,G14928);
  nand GNAME8874(G8874,G8870,G7628);
  nand GNAME8875(G8875,G7317,G36682);
  nand GNAME8876(G8876,G7195,G7626);
  nand GNAME8877(G8877,G7191,G7627);
  nand GNAME8878(G8878,G7547,G14936);
  nand GNAME8879(G8879,G8878,G8876,G8877);
  nand GNAME8880(G8880,G8172,G7622);
  nand GNAME8881(G8881,G7630,G14936);
  nand GNAME8882(G8882,G7725,G7624);
  nand GNAME8883(G8883,G14538,G7625);
  nand GNAME8884(G8884,G8879,G7628);
  nand GNAME8885(G8885,G7317,G36683);
  nand GNAME8886(G8886,G7181,G7626);
  nand GNAME8887(G8887,G7177,G7627);
  nand GNAME8888(G8888,G7547,G14931);
  nand GNAME8889(G8889,G8888,G8886,G8887);
  nand GNAME8890(G8890,G7566,G7629);
  nand GNAME8891(G8891,G14531,G7625);
  nand GNAME8892(G8892,G7630,G14931);
  nand GNAME8893(G8893,G8889,G7628);
  nand GNAME8894(G8894,G7317,G36684);
  and GNAME8895(G8895,G7547,G7628);
  or GNAME8896(G8896,G8895,G7630);
  nand GNAME8897(G8897,G8005,G7622);
  nand GNAME8898(G8898,G7628,G7217,G7627);
  nand GNAME8899(G8899,G8896,G36685);
  nand GNAME8900(G8900,G7721,G7624);
  nand GNAME8901(G8901,G14517,G7625);
  nand GNAME8902(G8902,G7317,G36685);
  nand GNAME8903(G8903,G7203,G7626);
  nand GNAME8904(G8904,G7199,G7627);
  nand GNAME8905(G8905,G7547,G14925);
  nand GNAME8906(G8906,G8905,G8903,G8904);
  nand GNAME8907(G8907,G8124,G7622);
  nand GNAME8908(G8908,G7630,G14925);
  nand GNAME8909(G8909,G7740,G7624);
  nand GNAME8910(G8910,G14518,G7625);
  nand GNAME8911(G8911,G8906,G7628);
  nand GNAME8912(G8912,G7317,G36686);
  nand GNAME8913(G8913,G7213,G7626);
  nand GNAME8914(G8914,G7209,G7627);
  nand GNAME8915(G8915,G7547,G14941);
  nand GNAME8916(G8916,G8915,G8913,G8914);
  nand GNAME8917(G8917,G8064,G7622);
  nand GNAME8918(G8918,G7630,G14941);
  nand GNAME8919(G8919,G7734,G7624);
  nand GNAME8920(G8920,G14521,G7625);
  nand GNAME8921(G8921,G8916,G7628);
  nand GNAME8922(G8922,G7317,G36687);
  nand GNAME8923(G8923,G7173,G7626);
  nand GNAME8924(G8924,G7169,G7627);
  nand GNAME8925(G8925,G7547,G14921);
  nand GNAME8926(G8926,G8925,G8923,G8924);
  nand GNAME8927(G8927,G7570,G7629);
  nand GNAME8928(G8928,G14527,G7625);
  nand GNAME8929(G8929,G7630,G14921);
  nand GNAME8930(G8930,G8926,G7628);
  nand GNAME8931(G8931,G7317,G36688);
  nand GNAME8932(G8932,G7187,G7626);
  nand GNAME8933(G8933,G7183,G7627);
  nand GNAME8934(G8934,G7547,G14930);
  nand GNAME8935(G8935,G8934,G8932,G8933);
  nand GNAME8936(G8936,G8220,G7622);
  nand GNAME8937(G8937,G7630,G14930);
  nand GNAME8938(G8938,G7728,G7624);
  nand GNAME8939(G8939,G14535,G7625);
  nand GNAME8940(G8940,G8935,G7628);
  nand GNAME8941(G8941,G7317,G36689);
  nand GNAME8942(G8942,G7211,G7626);
  nand GNAME8943(G8943,G7207,G7627);
  nand GNAME8944(G8944,G7547,G14933);
  nand GNAME8945(G8945,G8944,G8942,G8943);
  nand GNAME8946(G8946,G8076,G7622);
  nand GNAME8947(G8947,G7630,G14933);
  nand GNAME8948(G8948,G7738,G7624);
  nand GNAME8949(G8949,G14520,G7625);
  nand GNAME8950(G8950,G8945,G7628);
  nand GNAME8951(G8951,G7317,G36690);
  nand GNAME8952(G8952,G7189,G7626);
  nand GNAME8953(G8953,G7185,G7627);
  nand GNAME8954(G8954,G7547,G14918);
  nand GNAME8955(G8955,G8954,G8952,G8953);
  nand GNAME8956(G8956,G8208,G7622);
  nand GNAME8957(G8957,G7630,G14918);
  nand GNAME8958(G8958,G7726,G7624);
  nand GNAME8959(G8959,G14536,G7625);
  nand GNAME8960(G8960,G8955,G7628);
  nand GNAME8961(G8961,G7317,G36691);
  nand GNAME8962(G8962,G7171,G7626);
  nand GNAME8963(G8963,G7167,G7627);
  nand GNAME8964(G8964,G7547,G14927);
  nand GNAME8965(G8965,G8964,G8962,G8963);
  nand GNAME8966(G8966,G7571,G7629);
  nand GNAME8967(G8967,G14526,G7625);
  nand GNAME8968(G8968,G7630,G14927);
  nand GNAME8969(G8969,G8965,G7628);
  nand GNAME8970(G8970,G7317,G36692);
  nand GNAME8971(G8971,G7197,G7626);
  nand GNAME8972(G8972,G7193,G7627);
  nand GNAME8973(G8973,G7547,G14935);
  nand GNAME8974(G8974,G8973,G8971,G8972);
  nand GNAME8975(G8975,G8160,G7622);
  nand GNAME8976(G8976,G7630,G14935);
  nand GNAME8977(G8977,G7727,G7624);
  nand GNAME8978(G8978,G14539,G7625);
  nand GNAME8979(G8979,G8974,G7628);
  nand GNAME8980(G8980,G7317,G36693);
  nand GNAME8981(G8981,G7179,G7626);
  nand GNAME8982(G8982,G7175,G7627);
  nand GNAME8983(G8983,G7547,G14939);
  nand GNAME8984(G8984,G8983,G8981,G8982);
  nand GNAME8985(G8985,G7567,G7629);
  nand GNAME8986(G8986,G14530,G7625);
  nand GNAME8987(G8987,G7630,G14939);
  nand GNAME8988(G8988,G8984,G7628);
  nand GNAME8989(G8989,G7317,G36694);
  nand GNAME8990(G8990,G7219,G7626);
  nand GNAME8991(G8991,G7215,G7627);
  nand GNAME8992(G8992,G7547,G36695);
  nand GNAME8993(G8993,G8992,G8990,G8991);
  nand GNAME8994(G8994,G8027,G7622);
  nand GNAME8995(G8995,G7630,G36695);
  nand GNAME8996(G8996,G7733,G7624);
  nand GNAME8997(G8997,G14532,G7625);
  nand GNAME8998(G8998,G8993,G7628);
  nand GNAME8999(G8999,G7317,G36695);
  nand GNAME9000(G9000,G7205,G7626);
  nand GNAME9001(G9001,G7201,G7627);
  nand GNAME9002(G9002,G7547,G14923);
  nand GNAME9003(G9003,G9002,G9000,G9001);
  nand GNAME9004(G9004,G8112,G7622);
  nand GNAME9005(G9005,G7630,G14923);
  nand GNAME9006(G9006,G7732,G7624);
  nand GNAME9007(G9007,G14519,G7625);
  nand GNAME9008(G9008,G9003,G7628);
  nand GNAME9009(G9009,G7317,G36696);
  nand GNAME9010(G9010,G7165,G7626);
  nand GNAME9011(G9011,G7161,G7627);
  nand GNAME9012(G9012,G7547,G14940);
  nand GNAME9013(G9013,G9012,G9010,G9011);
  nand GNAME9014(G9014,G7574,G7629);
  nand GNAME9015(G9015,G14523,G7625);
  nand GNAME9016(G9016,G7630,G14940);
  nand GNAME9017(G9017,G9013,G7628);
  nand GNAME9018(G9018,G7317,G36697);
  nand GNAME9019(G9019,G7183,G7626);
  nand GNAME9020(G9020,G7179,G7627);
  nand GNAME9021(G9021,G7547,G14926);
  nand GNAME9022(G9022,G9021,G9019,G9020);
  nand GNAME9023(G9023,G8243,G7622);
  nand GNAME9024(G9024,G7630,G14926);
  nand GNAME9025(G9025,G7729,G7624);
  nand GNAME9026(G9026,G14533,G7625);
  nand GNAME9027(G9027,G9022,G7628);
  nand GNAME9028(G9028,G7317,G36698);
  nand GNAME9029(G9029,G7215,G7626);
  nand GNAME9030(G9030,G7211,G7627);
  nand GNAME9031(G9031,G7547,G14937);
  nand GNAME9032(G9032,G9031,G9029,G9030);
  nand GNAME9033(G9033,G8052,G7622);
  nand GNAME9034(G9034,G7630,G14937);
  nand GNAME9035(G9035,G7731,G7624);
  nand GNAME9036(G9036,G14469,G7625);
  nand GNAME9037(G9037,G9032,G7628);
  nand GNAME9038(G9038,G7317,G36699);
  nand GNAME9039(G9039,G7201,G7626);
  nand GNAME9040(G9040,G7197,G7627);
  nand GNAME9041(G9041,G7547,G14924);
  nand GNAME9042(G9042,G9041,G9039,G9040);
  nand GNAME9043(G9043,G8136,G7622);
  nand GNAME9044(G9044,G7630,G14924);
  nand GNAME9045(G9045,G7739,G7624);
  nand GNAME9046(G9046,G14463,G7625);
  nand GNAME9047(G9047,G9042,G7628);
  nand GNAME9048(G9048,G7317,G36700);
  nand GNAME9049(G9049,G7175,G7626);
  nand GNAME9050(G9050,G7171,G7627);
  nand GNAME9051(G9051,G7547,G14917);
  nand GNAME9052(G9052,G9051,G9049,G9050);
  nand GNAME9053(G9053,G7569,G7629);
  nand GNAME9054(G9054,G14528,G7625);
  nand GNAME9055(G9055,G7630,G14917);
  nand GNAME9056(G9056,G9052,G7628);
  nand GNAME9057(G9057,G7317,G36701);
  nand GNAME9058(G9058,G7193,G7626);
  nand GNAME9059(G9059,G7189,G7627);
  nand GNAME9060(G9060,G7547,G14942);
  nand GNAME9061(G9061,G9060,G9058,G9059);
  nand GNAME9062(G9062,G8184,G7622);
  nand GNAME9063(G9063,G7630,G14942);
  nand GNAME9064(G9064,G7724,G7624);
  nand GNAME9065(G9065,G14465,G7625);
  nand GNAME9066(G9066,G9061,G7628);
  nand GNAME9067(G9067,G7317,G36702);
  nand GNAME9068(G9068,G7167,G7626);
  nand GNAME9069(G9069,G7163,G7627);
  nand GNAME9070(G9070,G7547,G14934);
  nand GNAME9071(G9071,G9070,G9068,G9069);
  nand GNAME9072(G9072,G7573,G7629);
  nand GNAME9073(G9073,G14524,G7625);
  nand GNAME9074(G9074,G7630,G14934);
  nand GNAME9075(G9075,G9071,G7628);
  nand GNAME9076(G9076,G7317,G36703);
  nand GNAME9077(G9077,G7207,G7626);
  nand GNAME9078(G9078,G7203,G7627);
  nand GNAME9079(G9079,G7547,G14929);
  nand GNAME9080(G9080,G9079,G9077,G9078);
  nand GNAME9081(G9081,G8100,G7622);
  nand GNAME9082(G9082,G7630,G14929);
  nand GNAME9083(G9083,G7737,G7624);
  nand GNAME9084(G9084,G14471,G7625);
  nand GNAME9085(G9085,G9080,G7628);
  nand GNAME9086(G9086,G7317,G36704);
  nand GNAME9087(G9087,G9522,G7632);
  nand GNAME9088(G9088,G9087,G7841);
  nand GNAME9089(G9089,G9522,G7631);
  nand GNAME9090(G9090,G7562,G7659);
  nand GNAME9091(G9091,G9089,G9090);
  nand GNAME9092(G9092,G9091,G36600);
  nand GNAME9093(G9093,G9088,G36568);
  nand GNAME9094(G9094,G9091,G36599);
  nand GNAME9095(G9095,G9088,G36567);
  nand GNAME9096(G9096,G9091,G36598);
  nand GNAME9097(G9097,G9088,G36566);
  nand GNAME9098(G9098,G9091,G36597);
  nand GNAME9099(G9099,G9088,G36565);
  nand GNAME9100(G9100,G9091,G36596);
  nand GNAME9101(G9101,G9088,G36564);
  nand GNAME9102(G9102,G9091,G36595);
  nand GNAME9103(G9103,G9088,G36563);
  nand GNAME9104(G9104,G9091,G36594);
  nand GNAME9105(G9105,G9088,G36562);
  nand GNAME9106(G9106,G9091,G36593);
  nand GNAME9107(G9107,G9088,G36561);
  nand GNAME9108(G9108,G9091,G36610);
  nand GNAME9109(G9109,G9088,G36578);
  nand GNAME9110(G9110,G9091,G36609);
  nand GNAME9111(G9111,G9088,G36577);
  nand GNAME9112(G9112,G9091,G36608);
  nand GNAME9113(G9113,G9088,G36576);
  nand GNAME9114(G9114,G9091,G36607);
  nand GNAME9115(G9115,G9088,G36575);
  nand GNAME9116(G9116,G9091,G36606);
  nand GNAME9117(G9117,G9088,G36574);
  nand GNAME9118(G9118,G9091,G36605);
  nand GNAME9119(G9119,G9088,G36573);
  nand GNAME9120(G9120,G9091,G36604);
  nand GNAME9121(G9121,G9088,G36572);
  nand GNAME9122(G9122,G9091,G36603);
  nand GNAME9123(G9123,G9088,G36571);
  nand GNAME9124(G9124,G9091,G36602);
  nand GNAME9125(G9125,G9088,G36570);
  nand GNAME9126(G9126,G9091,G36601);
  nand GNAME9127(G9127,G9088,G36569);
  nand GNAME9128(G9128,G9091,G36592);
  nand GNAME9129(G9129,G9088,G36560);
  nand GNAME9130(G9130,G9091,G36591);
  nand GNAME9131(G9131,G9088,G36559);
  or GNAME9132(G9132,G7659,G9241);
  or GNAME9133(G9133,G7581,G7580,G7541);
  nand GNAME9134(G9134,G9171,G7740);
  nand GNAME9135(G9135,G7201,G9132);
  nand GNAME9136(G9136,G36600,G7648);
  nand GNAME9137(G9137,G36568,G7649);
  nand GNAME9138(G9138,G9171,G7732);
  nand GNAME9139(G9139,G7203,G9132);
  nand GNAME9140(G9140,G36599,G7648);
  nand GNAME9141(G9141,G36567,G7649);
  nand GNAME9142(G9142,G9171,G7737);
  nand GNAME9143(G9143,G7205,G9132);
  nand GNAME9144(G9144,G36598,G7648);
  nand GNAME9145(G9145,G36566,G7649);
  nand GNAME9146(G9146,G9171,G7736);
  nand GNAME9147(G9147,G7207,G9132);
  nand GNAME9148(G9148,G36597,G7648);
  nand GNAME9149(G9149,G36565,G7649);
  nand GNAME9150(G9150,G9171,G7738);
  nand GNAME9151(G9151,G7209,G9132);
  nand GNAME9152(G9152,G36596,G7648);
  nand GNAME9153(G9153,G36564,G7649);
  nand GNAME9154(G9154,G9171,G7734);
  nand GNAME9155(G9155,G7211,G9132);
  nand GNAME9156(G9156,G36595,G7648);
  nand GNAME9157(G9157,G36563,G7649);
  nand GNAME9158(G9158,G36610,G7648);
  nand GNAME9159(G9159,G36578,G7649);
  nand GNAME9160(G9160,G7163,G7646);
  nand GNAME9161(G9161,G7639,G7574);
  nand GNAME9162(G9162,G7161,G7647);
  nand GNAME9163(G9163,G7640,G7575);
  nand GNAME9164(G9164,G7157,G7659);
  nand GNAME9165(G9165,G7159,G7659);
  nand GNAME9166(G9166,G9171,G7731);
  nand GNAME9167(G9167,G7213,G9132);
  nand GNAME9168(G9168,G36594,G7648);
  nand GNAME9169(G9169,G36562,G7649);
  nand GNAME9170(G9170,G7161,G7659);
  or GNAME9171(G9171,G7639,G7640);
  nand GNAME9172(G9172,G7163,G9132);
  nand GNAME9173(G9173,G9171,G7574);
  nand GNAME9174(G9174,G7165,G9132);
  nand GNAME9175(G9175,G9171,G7573);
  nand GNAME9176(G9176,G7167,G9132);
  nand GNAME9177(G9177,G9171,G7572);
  nand GNAME9178(G9178,G7169,G9132);
  nand GNAME9179(G9179,G9171,G7571);
  nand GNAME9180(G9180,G7171,G9132);
  nand GNAME9181(G9181,G9171,G7570);
  nand GNAME9182(G9182,G7173,G9132);
  nand GNAME9183(G9183,G9171,G7569);
  nand GNAME9184(G9184,G7175,G9132);
  nand GNAME9185(G9185,G9171,G7568);
  nand GNAME9186(G9186,G7177,G9132);
  nand GNAME9187(G9187,G9171,G7567);
  nand GNAME9188(G9188,G7179,G9132);
  nand GNAME9189(G9189,G9171,G7566);
  nand GNAME9190(G9190,G9171,G7735);
  nand GNAME9191(G9191,G7215,G9132);
  nand GNAME9192(G9192,G36593,G7648);
  nand GNAME9193(G9193,G36561,G7649);
  nand GNAME9194(G9194,G9171,G7729);
  nand GNAME9195(G9195,G7181,G9132);
  nand GNAME9196(G9196,G9171,G7730);
  nand GNAME9197(G9197,G7183,G9132);
  nand GNAME9198(G9198,G36609,G7648);
  nand GNAME9199(G9199,G36577,G7649);
  nand GNAME9200(G9200,G9171,G7728);
  nand GNAME9201(G9201,G7185,G9132);
  nand GNAME9202(G9202,G36608,G7648);
  nand GNAME9203(G9203,G36576,G7649);
  nand GNAME9204(G9204,G9171,G7726);
  nand GNAME9205(G9205,G7187,G9132);
  nand GNAME9206(G9206,G36607,G7648);
  nand GNAME9207(G9207,G36575,G7649);
  nand GNAME9208(G9208,G9171,G7722);
  nand GNAME9209(G9209,G7189,G9132);
  nand GNAME9210(G9210,G36606,G7648);
  nand GNAME9211(G9211,G36574,G7649);
  nand GNAME9212(G9212,G9171,G7724);
  nand GNAME9213(G9213,G7191,G9132);
  nand GNAME9214(G9214,G36605,G7648);
  nand GNAME9215(G9215,G36573,G7649);
  nand GNAME9216(G9216,G9171,G7725);
  nand GNAME9217(G9217,G7193,G9132);
  nand GNAME9218(G9218,G36604,G7648);
  nand GNAME9219(G9219,G36572,G7649);
  nand GNAME9220(G9220,G9171,G7727);
  nand GNAME9221(G9221,G7195,G9132);
  nand GNAME9222(G9222,G36603,G7648);
  nand GNAME9223(G9223,G36571,G7649);
  nand GNAME9224(G9224,G9171,G7723);
  nand GNAME9225(G9225,G7197,G9132);
  nand GNAME9226(G9226,G36602,G7648);
  nand GNAME9227(G9227,G36570,G7649);
  nand GNAME9228(G9228,G9171,G7739);
  nand GNAME9229(G9229,G7199,G9132);
  nand GNAME9230(G9230,G36601,G7648);
  nand GNAME9231(G9231,G36569,G7649);
  nand GNAME9232(G9232,G9171,G7733);
  nand GNAME9233(G9233,G7217,G9132);
  nand GNAME9234(G9234,G36592,G7648);
  nand GNAME9235(G9235,G36560,G7649);
  nand GNAME9236(G9236,G9171,G7721);
  nand GNAME9237(G9237,G7219,G9132);
  nand GNAME9238(G9238,G36591,G7648);
  nand GNAME9239(G9239,G36559,G7649);
  or GNAME9240(G9240,G7649,G7648);
  or GNAME9241(G9241,G7646,G7647);
  nand GNAME9242(G9242,G9241,G7740);
  nand GNAME9243(G9243,G9240,G7679);
  nand GNAME9244(G9244,G7201,G9171);
  nand GNAME9245(G9245,G9241,G7732);
  nand GNAME9246(G9246,G9240,G7678);
  nand GNAME9247(G9247,G7203,G9171);
  nand GNAME9248(G9248,G9241,G7737);
  nand GNAME9249(G9249,G9240,G7677);
  nand GNAME9250(G9250,G7205,G9171);
  nand GNAME9251(G9251,G9241,G7736);
  nand GNAME9252(G9252,G9240,G7676);
  nand GNAME9253(G9253,G7207,G9171);
  nand GNAME9254(G9254,G9241,G7738);
  nand GNAME9255(G9255,G9240,G7675);
  nand GNAME9256(G9256,G7209,G9171);
  nand GNAME9257(G9257,G9241,G7734);
  nand GNAME9258(G9258,G9240,G7674);
  nand GNAME9259(G9259,G7211,G9171);
  nand GNAME9260(G9260,G7646,G7574);
  nand GNAME9261(G9261,G7163,G7639);
  nand GNAME9262(G9262,G7647,G7575);
  nand GNAME9263(G9263,G7161,G7640);
  nand GNAME9264(G9264,G9241,G7731);
  nand GNAME9265(G9265,G9240,G7673);
  nand GNAME9266(G9266,G7213,G9171);
  nand GNAME9267(G9267,G9241,G7574);
  nand GNAME9268(G9268,G7163,G9171);
  nand GNAME9269(G9269,G9241,G7573);
  nand GNAME9270(G9270,G7165,G9171);
  nand GNAME9271(G9271,G9241,G7572);
  nand GNAME9272(G9272,G7167,G9171);
  nand GNAME9273(G9273,G9241,G7571);
  nand GNAME9274(G9274,G7169,G9171);
  nand GNAME9275(G9275,G9241,G7570);
  nand GNAME9276(G9276,G7171,G9171);
  nand GNAME9277(G9277,G9241,G7569);
  nand GNAME9278(G9278,G7173,G9171);
  nand GNAME9279(G9279,G9241,G7568);
  nand GNAME9280(G9280,G7175,G9171);
  nand GNAME9281(G9281,G9241,G7567);
  nand GNAME9282(G9282,G7177,G9171);
  nand GNAME9283(G9283,G9241,G7566);
  nand GNAME9284(G9284,G7179,G9171);
  nand GNAME9285(G9285,G9241,G7735);
  nand GNAME9286(G9286,G9240,G7672);
  nand GNAME9287(G9287,G7215,G9171);
  nand GNAME9288(G9288,G9241,G7729);
  nand GNAME9289(G9289,G7181,G9171);
  nand GNAME9290(G9290,G9241,G7730);
  nand GNAME9291(G9291,G9240,G7688);
  nand GNAME9292(G9292,G7183,G9171);
  nand GNAME9293(G9293,G9241,G7728);
  nand GNAME9294(G9294,G9240,G7687);
  nand GNAME9295(G9295,G7185,G9171);
  nand GNAME9296(G9296,G9241,G7726);
  nand GNAME9297(G9297,G9240,G7686);
  nand GNAME9298(G9298,G7187,G9171);
  nand GNAME9299(G9299,G9241,G7722);
  nand GNAME9300(G9300,G9240,G7685);
  nand GNAME9301(G9301,G7189,G9171);
  nand GNAME9302(G9302,G9241,G7724);
  nand GNAME9303(G9303,G9240,G7684);
  nand GNAME9304(G9304,G7191,G9171);
  nand GNAME9305(G9305,G9241,G7725);
  nand GNAME9306(G9306,G9240,G7683);
  nand GNAME9307(G9307,G7193,G9171);
  nand GNAME9308(G9308,G9241,G7727);
  nand GNAME9309(G9309,G9240,G7682);
  nand GNAME9310(G9310,G7195,G9171);
  nand GNAME9311(G9311,G9241,G7723);
  nand GNAME9312(G9312,G9240,G7681);
  nand GNAME9313(G9313,G7197,G9171);
  nand GNAME9314(G9314,G9241,G7739);
  nand GNAME9315(G9315,G9240,G7680);
  nand GNAME9316(G9316,G7199,G9171);
  nand GNAME9317(G9317,G9241,G7733);
  nand GNAME9318(G9318,G9240,G7671);
  nand GNAME9319(G9319,G7217,G9171);
  nand GNAME9320(G9320,G9241,G7721);
  nand GNAME9321(G9321,G9240,G7669);
  nand GNAME9322(G9322,G7219,G9171);
  and GNAME9323(G9323,G7663,G9565);
  nand GNAME9324(G9324,G7844,G7654);
  nand GNAME9325(G9325,G7659,G7611);
  not GNAME9326(G9326,G7653);
  nand GNAME9327(G9327,G7652,G9326);
  nand GNAME9328(G9328,G7201,G9327);
  nand GNAME9329(G9329,G9324,G7740);
  nand GNAME9330(G9330,G7203,G9537);
  nand GNAME9331(G9331,G7203,G9327);
  nand GNAME9332(G9332,G9324,G7732);
  nand GNAME9333(G9333,G7205,G9537);
  nand GNAME9334(G9334,G7205,G9327);
  nand GNAME9335(G9335,G9324,G7737);
  nand GNAME9336(G9336,G7207,G9537);
  nand GNAME9337(G9337,G7207,G9327);
  nand GNAME9338(G9338,G9324,G7736);
  nand GNAME9339(G9339,G7209,G9537);
  nand GNAME9340(G9340,G7209,G9327);
  nand GNAME9341(G9341,G9324,G7738);
  nand GNAME9342(G9342,G7211,G9537);
  nand GNAME9343(G9343,G7211,G9327);
  nand GNAME9344(G9344,G9324,G7734);
  nand GNAME9345(G9345,G7213,G9537);
  nand GNAME9346(G9346,G7157,G9327);
  nand GNAME9347(G9347,G9324,G7579);
  nand GNAME9348(G9348,G7159,G9327);
  nand GNAME9349(G9349,G9324,G7578);
  nand GNAME9350(G9350,G7213,G9327);
  nand GNAME9351(G9351,G9324,G7731);
  nand GNAME9352(G9352,G7215,G9537);
  nand GNAME9353(G9353,G7161,G9327);
  nand GNAME9354(G9354,G9324,G7575);
  nand GNAME9355(G9355,G7163,G9537);
  nand GNAME9356(G9356,G7163,G9327);
  nand GNAME9357(G9357,G9324,G7574);
  nand GNAME9358(G9358,G7165,G9537);
  nand GNAME9359(G9359,G7165,G9327);
  nand GNAME9360(G9360,G9324,G7573);
  nand GNAME9361(G9361,G7167,G9537);
  nand GNAME9362(G9362,G7167,G9327);
  nand GNAME9363(G9363,G9324,G7572);
  nand GNAME9364(G9364,G7169,G9537);
  nand GNAME9365(G9365,G7169,G9327);
  nand GNAME9366(G9366,G9324,G7571);
  nand GNAME9367(G9367,G7171,G9537);
  nand GNAME9368(G9368,G7171,G9327);
  nand GNAME9369(G9369,G9324,G7570);
  nand GNAME9370(G9370,G7173,G9537);
  nand GNAME9371(G9371,G7173,G9327);
  nand GNAME9372(G9372,G9324,G7569);
  nand GNAME9373(G9373,G7175,G9537);
  nand GNAME9374(G9374,G7175,G9327);
  nand GNAME9375(G9375,G9324,G7568);
  nand GNAME9376(G9376,G7177,G9537);
  nand GNAME9377(G9377,G7177,G9327);
  nand GNAME9378(G9378,G9324,G7567);
  nand GNAME9379(G9379,G7179,G9537);
  nand GNAME9380(G9380,G7179,G9327);
  nand GNAME9381(G9381,G9324,G7566);
  nand GNAME9382(G9382,G7181,G9537);
  nand GNAME9383(G9383,G7215,G9327);
  nand GNAME9384(G9384,G9324,G7735);
  nand GNAME9385(G9385,G7217,G9537);
  nand GNAME9386(G9386,G7181,G9327);
  nand GNAME9387(G9387,G9324,G7729);
  nand GNAME9388(G9388,G7183,G9537);
  nand GNAME9389(G9389,G7183,G9327);
  nand GNAME9390(G9390,G9324,G7730);
  nand GNAME9391(G9391,G7185,G9537);
  nand GNAME9392(G9392,G7185,G9327);
  nand GNAME9393(G9393,G9324,G7728);
  nand GNAME9394(G9394,G7187,G9537);
  nand GNAME9395(G9395,G7187,G9327);
  nand GNAME9396(G9396,G9324,G7726);
  nand GNAME9397(G9397,G7189,G9537);
  nand GNAME9398(G9398,G7189,G9327);
  nand GNAME9399(G9399,G9324,G7722);
  nand GNAME9400(G9400,G7191,G9537);
  nand GNAME9401(G9401,G7191,G9327);
  nand GNAME9402(G9402,G9324,G7724);
  nand GNAME9403(G9403,G7193,G9537);
  nand GNAME9404(G9404,G7193,G9327);
  nand GNAME9405(G9405,G9324,G7725);
  nand GNAME9406(G9406,G7195,G9537);
  nand GNAME9407(G9407,G7195,G9327);
  nand GNAME9408(G9408,G9324,G7727);
  nand GNAME9409(G9409,G7197,G9537);
  nand GNAME9410(G9410,G7197,G9327);
  nand GNAME9411(G9411,G9324,G7723);
  nand GNAME9412(G9412,G7199,G9537);
  nand GNAME9413(G9413,G7199,G9327);
  nand GNAME9414(G9414,G9324,G7739);
  nand GNAME9415(G9415,G7201,G9537);
  nand GNAME9416(G9416,G7217,G9327);
  nand GNAME9417(G9417,G9324,G7733);
  nand GNAME9418(G9418,G7219,G9537);
  nand GNAME9419(G9419,G7219,G9327);
  nand GNAME9420(G9420,G9324,G7721);
  or GNAME9421(G9421,G791,G7844);
  nand GNAME9422(G9422,G9421,G7654);
  nand GNAME9423(G9423,G7655,G7201);
  nand GNAME9424(G9424,G7201,G9422);
  nand GNAME9425(G9425,G7653,G7740);
  nand GNAME9426(G9426,G7655,G7203);
  nand GNAME9427(G9427,G7203,G9422);
  nand GNAME9428(G9428,G7653,G7732);
  nand GNAME9429(G9429,G7655,G7205);
  nand GNAME9430(G9430,G7205,G9422);
  nand GNAME9431(G9431,G7653,G7737);
  nand GNAME9432(G9432,G7655,G7207);
  nand GNAME9433(G9433,G7207,G9422);
  nand GNAME9434(G9434,G7653,G7736);
  nand GNAME9435(G9435,G7655,G7209);
  nand GNAME9436(G9436,G7209,G9422);
  nand GNAME9437(G9437,G7653,G7738);
  nand GNAME9438(G9438,G7655,G7211);
  nand GNAME9439(G9439,G7211,G9422);
  nand GNAME9440(G9440,G7653,G7734);
  nand GNAME9441(G9441,G7655,G14914);
  nand GNAME9442(G9442,G7157,G9422);
  nand GNAME9443(G9443,G7653,G7579);
  nand GNAME9444(G9444,G7655,G14913);
  nand GNAME9445(G9445,G7159,G9422);
  nand GNAME9446(G9446,G7653,G7578);
  nand GNAME9447(G9447,G7655,G7213);
  nand GNAME9448(G9448,G7213,G9422);
  nand GNAME9449(G9449,G7653,G7731);
  nand GNAME9450(G9450,G7655,G7161);
  nand GNAME9451(G9451,G7161,G9422);
  nand GNAME9452(G9452,G7653,G7575);
  nand GNAME9453(G9453,G7655,G7163);
  nand GNAME9454(G9454,G7163,G9422);
  nand GNAME9455(G9455,G7653,G7574);
  nand GNAME9456(G9456,G7655,G7165);
  nand GNAME9457(G9457,G7165,G9422);
  nand GNAME9458(G9458,G7653,G7573);
  nand GNAME9459(G9459,G7655,G7167);
  nand GNAME9460(G9460,G7167,G9422);
  nand GNAME9461(G9461,G7653,G7572);
  nand GNAME9462(G9462,G7655,G7169);
  nand GNAME9463(G9463,G7169,G9422);
  nand GNAME9464(G9464,G7653,G7571);
  nand GNAME9465(G9465,G7655,G7171);
  nand GNAME9466(G9466,G7171,G9422);
  nand GNAME9467(G9467,G7653,G7570);
  nand GNAME9468(G9468,G7655,G7173);
  nand GNAME9469(G9469,G7173,G9422);
  nand GNAME9470(G9470,G7653,G7569);
  nand GNAME9471(G9471,G7655,G7175);
  nand GNAME9472(G9472,G7175,G9422);
  nand GNAME9473(G9473,G7653,G7568);
  nand GNAME9474(G9474,G7655,G7177);
  nand GNAME9475(G9475,G7177,G9422);
  nand GNAME9476(G9476,G7653,G7567);
  nand GNAME9477(G9477,G7655,G7179);
  nand GNAME9478(G9478,G7179,G9422);
  nand GNAME9479(G9479,G7653,G7566);
  nand GNAME9480(G9480,G7655,G7215);
  nand GNAME9481(G9481,G7215,G9422);
  nand GNAME9482(G9482,G7653,G7735);
  nand GNAME9483(G9483,G7655,G7181);
  nand GNAME9484(G9484,G7181,G9422);
  nand GNAME9485(G9485,G7653,G7729);
  nand GNAME9486(G9486,G7655,G7183);
  nand GNAME9487(G9487,G7183,G9422);
  nand GNAME9488(G9488,G7653,G7730);
  nand GNAME9489(G9489,G7655,G7185);
  nand GNAME9490(G9490,G7185,G9422);
  nand GNAME9491(G9491,G7653,G7728);
  nand GNAME9492(G9492,G7655,G7187);
  nand GNAME9493(G9493,G7187,G9422);
  nand GNAME9494(G9494,G7653,G7726);
  nand GNAME9495(G9495,G7655,G7189);
  nand GNAME9496(G9496,G7189,G9422);
  nand GNAME9497(G9497,G7653,G7722);
  nand GNAME9498(G9498,G7655,G7191);
  nand GNAME9499(G9499,G7191,G9422);
  nand GNAME9500(G9500,G7653,G7724);
  nand GNAME9501(G9501,G7655,G7193);
  nand GNAME9502(G9502,G7193,G9422);
  nand GNAME9503(G9503,G7653,G7725);
  nand GNAME9504(G9504,G7655,G7195);
  nand GNAME9505(G9505,G7195,G9422);
  nand GNAME9506(G9506,G7653,G7727);
  nand GNAME9507(G9507,G7655,G7197);
  nand GNAME9508(G9508,G7197,G9422);
  nand GNAME9509(G9509,G7653,G7723);
  nand GNAME9510(G9510,G7655,G7199);
  nand GNAME9511(G9511,G7199,G9422);
  nand GNAME9512(G9512,G7653,G7739);
  nand GNAME9513(G9513,G7655,G7217);
  nand GNAME9514(G9514,G7217,G9422);
  nand GNAME9515(G9515,G7653,G7733);
  nand GNAME9516(G9516,G7655,G7219);
  nand GNAME9517(G9517,G7219,G9422);
  nand GNAME9518(G9518,G7653,G7721);
  nand GNAME9519(G9519,G7545,G7621);
  nand GNAME9520(G9520,G7609,G8692,G7670);
  or GNAME9521(G9521,G7546,G7580,G7581);
  nand GNAME9522(G9522,G7607,G7848,G7861);
  nand GNAME9523(G9523,G9525,G9630,G9631);
  nand GNAME9524(G9524,G7872,G9520);
  or GNAME9525(G9525,G7317,G7670,G7610,G9537);
  nand GNAME9526(G9526,G7533,G36488);
  nand GNAME9527(G9527,G14406,G36494);
  nand GNAME9528(G9528,G7533,G36489);
  nand GNAME9529(G9529,G14375,G36494);
  nand GNAME9530(G9530,G9528,G9529);
  nand GNAME9531(G9531,G7533,G36487);
  nand GNAME9532(G9532,G14407,G36494);
  or GNAME9533(G9533,G36675,G7534);
  or GNAME9534(G9534,G7537,G7658,G7536);
  nand GNAME9535(G9535,G7533,G36486);
  nand GNAME9536(G9536,G14374,G36494);
  not GNAME9537(G9537,G7659);
  nand GNAME9538(G9538,G7868,G36495);
  nand GNAME9539(G9539,G7982,G7835);
  nand GNAME9540(G9540,G7868,G36496);
  nand GNAME9541(G9541,G7983,G7835);
  nand GNAME9542(G9542,G7533,G36492,G36493);
  nand GNAME9543(G9543,G36494,G14377,G14404);
  nand GNAME9544(G9544,G9542,G9543);
  nand GNAME9545(G9545,G7533,G7531,G36493);
  nand GNAME9546(G9546,G36494,G7530,G14404);
  nand GNAME9547(G9547,G9545,G9546);
  nand GNAME9548(G9548,G7533,G7532,G36492);
  or GNAME9549(G9549,G7533,G14404,G7530);
  nand GNAME9550(G9550,G9548,G9549);
  or GNAME9551(G9551,G36494,G36493,G36492);
  or GNAME9552(G9552,G7533,G14377,G14404);
  nand GNAME9553(G9553,G9551,G9552);
  or GNAME9554(G9554,G36494,G36491,G36490);
  or GNAME9555(G9555,G7533,G14376,G14405);
  not GNAME9556(G9556,G7662);
  nand GNAME9557(G9557,G7533,G36484);
  nand GNAME9558(G9558,G14408,G36494);
  not GNAME9559(G9559,G7663);
  nand GNAME9560(G9560,G7533,G36485);
  nand GNAME9561(G9561,G14373,G36494);
  not GNAME9562(G9562,G7664);
  nand GNAME9563(G9563,G7533,G36483);
  nand GNAME9564(G9564,G14409,G36494);
  not GNAME9565(G9565,G7666);
  nand GNAME9566(G9566,G7533,G36482);
  nand GNAME9567(G9567,G14372,G36494);
  not GNAME9568(G9568,G7665);
  nand GNAME9569(G9569,G7981,G36496);
  nand GNAME9570(G9570,G7539,G7983);
  not GNAME9571(G9571,G7667);
  nand GNAME9572(G9572,G7981,G36495);
  nand GNAME9573(G9573,G7539,G7982);
  not GNAME9574(G9574,G7668);
  nand GNAME9575(G9575,G7533,G36463);
  nand GNAME9576(G9576,G36463,G36494);
  nand GNAME9577(G9577,G7533,G36491);
  nand GNAME9578(G9578,G14405,G36494);
  not GNAME9579(G9579,G7670);
  nand GNAME9580(G9580,G7528,G7548);
  or GNAME9581(G9581,G7528,G14376,G7533);
  nand GNAME9582(G9582,G7529,G7549);
  or GNAME9583(G9583,G7529,G36490,G36494);
  nand GNAME9584(G9584,G7533,G36464);
  nand GNAME9585(G9585,G14397,G36494);
  nand GNAME9586(G9586,G7533,G36465);
  nand GNAME9587(G9587,G14378,G36494);
  nand GNAME9588(G9588,G7533,G36466);
  nand GNAME9589(G9589,G14379,G36494);
  nand GNAME9590(G9590,G7533,G36467);
  nand GNAME9591(G9591,G14402,G36494);
  nand GNAME9592(G9592,G7533,G36468);
  nand GNAME9593(G9593,G14401,G36494);
  nand GNAME9594(G9594,G7533,G36469);
  nand GNAME9595(G9595,G14380,G36494);
  nand GNAME9596(G9596,G7533,G36470);
  nand GNAME9597(G9597,G14381,G36494);
  nand GNAME9598(G9598,G7533,G36471);
  nand GNAME9599(G9599,G14400,G36494);
  nand GNAME9600(G9600,G7533,G36472);
  nand GNAME9601(G9601,G14399,G36494);
  nand GNAME9602(G9602,G7533,G36473);
  nand GNAME9603(G9603,G14367,G36494);
  nand GNAME9604(G9604,G7533,G36474);
  nand GNAME9605(G9605,G14368,G36494);
  nand GNAME9606(G9606,G7533,G36475);
  nand GNAME9607(G9607,G14414,G36494);
  nand GNAME9608(G9608,G7533,G36476);
  nand GNAME9609(G9609,G14413,G36494);
  nand GNAME9610(G9610,G7533,G36477);
  nand GNAME9611(G9611,G14369,G36494);
  nand GNAME9612(G9612,G7533,G36478);
  nand GNAME9613(G9613,G14370,G36494);
  nand GNAME9614(G9614,G7533,G36479);
  nand GNAME9615(G9615,G14412,G36494);
  nand GNAME9616(G9616,G7533,G36480);
  nand GNAME9617(G9617,G14411,G36494);
  nand GNAME9618(G9618,G7533,G36481);
  nand GNAME9619(G9619,G14371,G36494);
  nand GNAME9620(G9620,G7553,G36556);
  nand GNAME9621(G9621,G7869,G7836);
  nand GNAME9622(G9622,G7991,G9562);
  nand GNAME9623(G9623,G7561,G9568);
  nand GNAME9624(G9624,G7584,G36588);
  nand GNAME9625(G9625,G7870,G7836);
  nand GNAME9626(G9626,G7590,G36592);
  nand GNAME9627(G9627,G7871,G8513,G14532);
  nand GNAME9628(G9628,G7590,G36620);
  nand GNAME9629(G9629,G7871,G7836);
  nand GNAME9630(G9630,G7605,G7670);
  nand GNAME9631(G9631,G9579,G8692,G7609);
  nand GNAME9632(G9632,G7867,G36643);
  nand GNAME9633(G9633,G7219,G7605);
  nand GNAME9634(G9634,G7867,G36644);
  nand GNAME9635(G9635,G7217,G7605);
  nand GNAME9636(G9636,G7867,G36645);
  nand GNAME9637(G9637,G7215,G7605);
  nand GNAME9638(G9638,G7867,G36646);
  nand GNAME9639(G9639,G7213,G7605);
  nand GNAME9640(G9640,G7867,G36647);
  nand GNAME9641(G9641,G7211,G7605);
  nand GNAME9642(G9642,G7867,G36648);
  nand GNAME9643(G9643,G7209,G7605);
  nand GNAME9644(G9644,G7867,G36649);
  nand GNAME9645(G9645,G7207,G7605);
  nand GNAME9646(G9646,G7867,G36650);
  nand GNAME9647(G9647,G7205,G7605);
  nand GNAME9648(G9648,G7867,G36651);
  nand GNAME9649(G9649,G7203,G7605);
  nand GNAME9650(G9650,G7867,G36652);
  nand GNAME9651(G9651,G7201,G7605);
  nand GNAME9652(G9652,G7867,G36653);
  nand GNAME9653(G9653,G7199,G7605);
  nand GNAME9654(G9654,G7867,G36654);
  nand GNAME9655(G9655,G7197,G7605);
  nand GNAME9656(G9656,G7867,G36655);
  nand GNAME9657(G9657,G7195,G7605);
  nand GNAME9658(G9658,G7867,G36656);
  nand GNAME9659(G9659,G7193,G7605);
  nand GNAME9660(G9660,G7867,G36657);
  nand GNAME9661(G9661,G7191,G7605);
  nand GNAME9662(G9662,G7867,G36658);
  nand GNAME9663(G9663,G7189,G7605);
  nand GNAME9664(G9664,G7867,G36659);
  nand GNAME9665(G9665,G7187,G7605);
  nand GNAME9666(G9666,G7867,G36660);
  nand GNAME9667(G9667,G7185,G7605);
  nand GNAME9668(G9668,G7867,G36661);
  nand GNAME9669(G9669,G7183,G7605);
  nand GNAME9670(G9670,G7867,G36662);
  nand GNAME9671(G9671,G7181,G7605);
  nand GNAME9672(G9672,G7867,G36663);
  nand GNAME9673(G9673,G7179,G7605);
  nand GNAME9674(G9674,G7867,G36664);
  nand GNAME9675(G9675,G7177,G7605);
  nand GNAME9676(G9676,G7867,G36665);
  nand GNAME9677(G9677,G7175,G7605);
  nand GNAME9678(G9678,G7867,G36666);
  nand GNAME9679(G9679,G7173,G7605);
  nand GNAME9680(G9680,G7867,G36667);
  nand GNAME9681(G9681,G7171,G7605);
  nand GNAME9682(G9682,G7867,G36668);
  nand GNAME9683(G9683,G7169,G7605);
  nand GNAME9684(G9684,G7867,G36669);
  nand GNAME9685(G9685,G7167,G7605);
  nand GNAME9686(G9686,G7867,G36670);
  nand GNAME9687(G9687,G7165,G7605);
  nand GNAME9688(G9688,G7867,G36671);
  nand GNAME9689(G9689,G7163,G7605);
  nand GNAME9690(G9690,G7867,G36672);
  nand GNAME9691(G9691,G7161,G7605);
  nand GNAME9692(G9692,G7867,G36673);
  nand GNAME9693(G9693,G7159,G7605);
  nand GNAME9694(G9694,G7867,G36674);
  nand GNAME9695(G9695,G7157,G7605);
  nand GNAME9696(G9696,G7613,G9559,G7600);
  or GNAME9697(G9697,G7613,G7620);
  nand GNAME9698(G9698,G7866,G814);
  nand GNAME9699(G9699,G7671,G7839);
  not GNAME9700(G9700,G7733);
  nand GNAME9701(G9701,G7988,G9700);
  nand GNAME9702(G9702,G7217,G7733);
  nand GNAME9703(G9703,G9701,G9702);
  nand GNAME9704(G9704,G7866,G800);
  nand GNAME9705(G9705,G7673,G7839);
  not GNAME9706(G9706,G7731);
  nand GNAME9707(G9707,G8038,G9706);
  nand GNAME9708(G9708,G7213,G7731);
  nand GNAME9709(G9709,G9707,G9708);
  nand GNAME9710(G9710,G7866,G795);
  nand GNAME9711(G9711,G7678,G7839);
  not GNAME9712(G9712,G7732);
  nand GNAME9713(G9713,G8098,G9712);
  nand GNAME9714(G9714,G7203,G7732);
  nand GNAME9715(G9715,G9713,G9714);
  nand GNAME9716(G9716,G7866,G799);
  nand GNAME9717(G9717,G7674,G7839);
  not GNAME9718(G9718,G7734);
  nand GNAME9719(G9719,G8050,G9718);
  nand GNAME9720(G9720,G7211,G7734);
  nand GNAME9721(G9721,G9719,G9720);
  nand GNAME9722(G9722,G7866,G803);
  nand GNAME9723(G9723,G7672,G7839);
  not GNAME9724(G9724,G7735);
  nand GNAME9725(G9725,G8020,G9724);
  nand GNAME9726(G9726,G7215,G7735);
  nand GNAME9727(G9727,G9725,G9726);
  nand GNAME9728(G9728,G7866,G798);
  nand GNAME9729(G9729,G7675,G7839);
  not GNAME9730(G9730,G7738);
  nand GNAME9731(G9731,G8062,G9730);
  nand GNAME9732(G9732,G7209,G7738);
  nand GNAME9733(G9733,G9731,G9732);
  nand GNAME9734(G9734,G7866,G797);
  nand GNAME9735(G9735,G7676,G7839);
  not GNAME9736(G9736,G7736);
  nand GNAME9737(G9737,G8074,G9736);
  nand GNAME9738(G9738,G7207,G7736);
  nand GNAME9739(G9739,G9737,G9738);
  nand GNAME9740(G9740,G7866,G796);
  nand GNAME9741(G9741,G7677,G7839);
  not GNAME9742(G9742,G7737);
  nand GNAME9743(G9743,G8086,G9742);
  nand GNAME9744(G9744,G7205,G7737);
  nand GNAME9745(G9745,G9743,G9744);
  nand GNAME9746(G9746,G7866,G824);
  nand GNAME9747(G9747,G7680,G7839);
  not GNAME9748(G9748,G7739);
  nand GNAME9749(G9749,G8122,G9748);
  nand GNAME9750(G9750,G7199,G7739);
  nand GNAME9751(G9751,G9749,G9750);
  nand GNAME9752(G9752,G7866,G794);
  nand GNAME9753(G9753,G7679,G7839);
  not GNAME9754(G9754,G7740);
  nand GNAME9755(G9755,G8110,G9754);
  nand GNAME9756(G9756,G7201,G7740);
  nand GNAME9757(G9757,G9755,G9756);
  nand GNAME9758(G9758,G7177,G7567);
  or GNAME9759(G9759,G7567,G7177);
  nand GNAME9760(G9760,G9758,G9759);
  nand GNAME9761(G9761,G7171,G7570);
  or GNAME9762(G9762,G7570,G7171);
  nand GNAME9763(G9763,G9761,G9762);
  nand GNAME9764(G9764,G7159,G7578);
  or GNAME9765(G9765,G7578,G7159);
  nand GNAME9766(G9766,G9764,G9765);
  nand GNAME9767(G9767,G7173,G7569);
  or GNAME9768(G9768,G7569,G7173);
  nand GNAME9769(G9769,G9767,G9768);
  nand GNAME9770(G9770,G7161,G7575);
  or GNAME9771(G9771,G7161,G7575);
  nand GNAME9772(G9772,G9770,G9771);
  nand GNAME9773(G9773,G7169,G7571);
  or GNAME9774(G9774,G7571,G7169);
  nand GNAME9775(G9775,G9773,G9774);
  nand GNAME9776(G9776,G7165,G7573);
  or GNAME9777(G9777,G7573,G7165);
  nand GNAME9778(G9778,G9776,G9777);
  nand GNAME9779(G9779,G7179,G7566);
  or GNAME9780(G9780,G7566,G7179);
  nand GNAME9781(G9781,G9779,G9780);
  nand GNAME9782(G9782,G7175,G7568);
  or GNAME9783(G9783,G7568,G7175);
  nand GNAME9784(G9784,G9782,G9783);
  nand GNAME9785(G9785,G7157,G7579);
  or GNAME9786(G9786,G7579,G7157);
  nand GNAME9787(G9787,G9785,G9786);
  nand GNAME9788(G9788,G7163,G7574);
  or GNAME9789(G9789,G7163,G7574);
  nand GNAME9790(G9790,G9788,G9789);
  nand GNAME9791(G9791,G7866,G823);
  nand GNAME9792(G9792,G7681,G7839);
  not GNAME9793(G9793,G7723);
  nand GNAME9794(G9794,G8134,G9793);
  nand GNAME9795(G9795,G7197,G7723);
  nand GNAME9796(G9796,G9794,G9795);
  nand GNAME9797(G9797,G7167,G7572);
  or GNAME9798(G9798,G7572,G7167);
  nand GNAME9799(G9799,G9797,G9798);
  nand GNAME9800(G9800,G7866,G819);
  nand GNAME9801(G9801,G7685,G7839);
  not GNAME9802(G9802,G7722);
  nand GNAME9803(G9803,G8182,G9802);
  nand GNAME9804(G9804,G7189,G7722);
  nand GNAME9805(G9805,G9803,G9804);
  nand GNAME9806(G9806,G7866,G820);
  nand GNAME9807(G9807,G7684,G7839);
  not GNAME9808(G9808,G7724);
  nand GNAME9809(G9809,G8170,G9808);
  nand GNAME9810(G9810,G7191,G7724);
  nand GNAME9811(G9811,G9809,G9810);
  nand GNAME9812(G9812,G7866,G821);
  nand GNAME9813(G9813,G7683,G7839);
  not GNAME9814(G9814,G7725);
  nand GNAME9815(G9815,G8158,G9814);
  nand GNAME9816(G9816,G7193,G7725);
  nand GNAME9817(G9817,G9815,G9816);
  nand GNAME9818(G9818,G7866,G817);
  nand GNAME9819(G9819,G7687,G7839);
  not GNAME9820(G9820,G7728);
  nand GNAME9821(G9821,G8206,G9820);
  nand GNAME9822(G9822,G7185,G7728);
  nand GNAME9823(G9823,G9821,G9822);
  nand GNAME9824(G9824,G7866,G818);
  nand GNAME9825(G9825,G7686,G7839);
  not GNAME9826(G9826,G7726);
  nand GNAME9827(G9827,G8194,G9826);
  nand GNAME9828(G9828,G7187,G7726);
  nand GNAME9829(G9829,G9827,G9828);
  nand GNAME9830(G9830,G7866,G822);
  nand GNAME9831(G9831,G7682,G7839);
  not GNAME9832(G9832,G7727);
  nand GNAME9833(G9833,G8146,G9832);
  nand GNAME9834(G9834,G7195,G7727);
  nand GNAME9835(G9835,G9833,G9834);
  nand GNAME9836(G9836,G7866,G815);
  nand GNAME9837(G9837,G7665,G7839);
  not GNAME9838(G9838,G7729);
  nand GNAME9839(G9839,G8230,G9838);
  nand GNAME9840(G9840,G7181,G7729);
  nand GNAME9841(G9841,G9839,G9840);
  nand GNAME9842(G9842,G7866,G816);
  nand GNAME9843(G9843,G7688,G7839);
  not GNAME9844(G9844,G7730);
  nand GNAME9845(G9845,G8218,G9844);
  nand GNAME9846(G9846,G7183,G7730);
  nand GNAME9847(G9847,G9845,G9846);
  nand GNAME9848(G9848,G7866,G825);
  nand GNAME9849(G9849,G7669,G7839);
  not GNAME9850(G9850,G7721);
  nand GNAME9851(G9851,G8025,G9850);
  nand GNAME9852(G9852,G7219,G7721);
  nand GNAME9853(G9853,G9851,G9852);
  nand GNAME9854(G9854,G14239,G9559);
  nand GNAME9855(G9855,G7613,G7663);
  nand GNAME9856(G9856,G9565,G9854,G9855);
  nand GNAME9857(G9857,G7666,G8782,G8780,G8781);
  nand GNAME9858(G9858,G14518,G14239);
  nand GNAME9859(G9859,G7613,G7201);
  nand GNAME9860(G9860,G14519,G14239);
  nand GNAME9861(G9861,G7613,G7203);
  nand GNAME9862(G9862,G14471,G14239);
  nand GNAME9863(G9863,G7613,G7205);
  nand GNAME9864(G9864,G14470,G14239);
  nand GNAME9865(G9865,G7613,G7207);
  nand GNAME9866(G9866,G14520,G14239);
  nand GNAME9867(G9867,G7613,G7209);
  nand GNAME9868(G9868,G14521,G14239);
  nand GNAME9869(G9869,G7613,G7211);
  nand GNAME9870(G9870,G14239,G14468);
  nand GNAME9871(G9871,G7613,G7157);
  nand GNAME9872(G9872,G14239,G14467);
  nand GNAME9873(G9873,G7613,G7159);
  nand GNAME9874(G9874,G14469,G14239);
  nand GNAME9875(G9875,G7613,G7213);
  nand GNAME9876(G9876,G14522,G14239);
  nand GNAME9877(G9877,G7613,G7161);
  nand GNAME9878(G9878,G14523,G14239);
  nand GNAME9879(G9879,G7613,G7163);
  nand GNAME9880(G9880,G14524,G14239);
  nand GNAME9881(G9881,G7613,G7165);
  nand GNAME9882(G9882,G14525,G14239);
  nand GNAME9883(G9883,G7613,G7167);
  nand GNAME9884(G9884,G14526,G14239);
  nand GNAME9885(G9885,G7613,G7169);
  nand GNAME9886(G9886,G14527,G14239);
  nand GNAME9887(G9887,G7613,G7171);
  nand GNAME9888(G9888,G14528,G14239);
  nand GNAME9889(G9889,G7613,G7173);
  nand GNAME9890(G9890,G14529,G14239);
  nand GNAME9891(G9891,G7613,G7175);
  nand GNAME9892(G9892,G14530,G14239);
  nand GNAME9893(G9893,G7613,G7177);
  nand GNAME9894(G9894,G14531,G14239);
  nand GNAME9895(G9895,G7613,G7179);
  nand GNAME9896(G9896,G14466,G14239);
  nand GNAME9897(G9897,G7613,G7215);
  nand GNAME9898(G9898,G14533,G14239);
  nand GNAME9899(G9899,G7613,G7181);
  nand GNAME9900(G9900,G14534,G14239);
  nand GNAME9901(G9901,G7613,G7183);
  nand GNAME9902(G9902,G14535,G14239);
  nand GNAME9903(G9903,G7613,G7185);
  nand GNAME9904(G9904,G14536,G14239);
  nand GNAME9905(G9905,G7613,G7187);
  nand GNAME9906(G9906,G14537,G14239);
  nand GNAME9907(G9907,G7613,G7189);
  nand GNAME9908(G9908,G14465,G14239);
  nand GNAME9909(G9909,G7613,G7191);
  nand GNAME9910(G9910,G14538,G14239);
  nand GNAME9911(G9911,G7613,G7193);
  nand GNAME9912(G9912,G14539,G14239);
  nand GNAME9913(G9913,G7613,G7195);
  nand GNAME9914(G9914,G14464,G14239);
  nand GNAME9915(G9915,G7613,G7197);
  nand GNAME9916(G9916,G14463,G14239);
  nand GNAME9917(G9917,G7613,G7199);
  nand GNAME9918(G9918,G14532,G14239);
  nand GNAME9919(G9919,G7613,G7217);
  nand GNAME9920(G9920,G14517,G14239);
  nand GNAME9921(G9921,G7613,G7219);
  not GNAME9922(G9922,G7538);
  nand GNAME9923(G9923,G15012,G7761);
  or GNAME9924(G9924,G7730,G15011);
  nand GNAME9925(G9925,G9926,G9928,G9927);
  nand GNAME9926(G9926,G15011,G7730);
  or GNAME9927(G9927,G7763,G15010);
  nand GNAME9928(G9928,G9929,G9931,G9930);
  nand GNAME9929(G9929,G15010,G7763);
  or GNAME9930(G9930,G7726,G15009);
  nand GNAME9931(G9931,G15071,G15069,G15070);
  not GNAME9932(G9932,G36133);
  not GNAME9933(G9933,G36623);
  and GNAME9934(G9934,G10071,G10072);
  and GNAME9935(G9935,G10067,G10069);
  and GNAME9936(G9936,G10064,G10066);
  and GNAME9937(G9937,G10062,G10063);
  and GNAME9938(G9938,G10057,G10059);
  nand GNAME9939(G9939,G10076,G10111,G10112);
  not GNAME9940(G9940,G36152);
  nand GNAME9941(G9941,G36397,G36152);
  not GNAME9942(G9942,G36396);
  not GNAME9943(G9943,G36150);
  not GNAME9944(G9944,G36395);
  not GNAME9945(G9945,G36149);
  not GNAME9946(G9946,G36394);
  not GNAME9947(G9947,G36145);
  not GNAME9948(G9948,G36390);
  not GNAME9949(G9949,G36144);
  not GNAME9950(G9950,G36389);
  not GNAME9951(G9951,G36388);
  not GNAME9952(G9952,G36143);
  not GNAME9953(G9953,G36386);
  not GNAME9954(G9954,G36140);
  not GNAME9955(G9955,G36385);
  not GNAME9956(G9956,G36139);
  not GNAME9957(G9957,G36384);
  not GNAME9958(G9958,G36381);
  not GNAME9959(G9959,G36136);
  nor GNAME9960(G9960,G10145,G9966);
  not GNAME9961(G9961,G36380);
  not GNAME9962(G9962,G36135);
  and GNAME9963(G9963,G10051,G10052);
  not GNAME9964(G9964,G36379);
  not GNAME9965(G9965,G36134);
  and GNAME9966(G9966,G10045,G10060);
  or GNAME9967(G9967,G10044,G9968);
  and GNAME9968(G9968,G10042,G10043);
  and GNAME9969(G9969,G10035,G10036);
  and GNAME9970(G9970,G10032,G10033);
  or GNAME9971(G9971,G10034,G9970);
  nand GNAME9972(G9972,G10143,G10144);
  nand GNAME9973(G9973,G10080,G10081);
  nand GNAME9974(G9974,G10085,G10086);
  nand GNAME9975(G9975,G10090,G10091);
  nand GNAME9976(G9976,G10092,G10093);
  nand GNAME9977(G9977,G10094,G10095);
  nand GNAME9978(G9978,G10096,G10097);
  nand GNAME9979(G9979,G10101,G10102);
  nand GNAME9980(G9980,G10106,G10107);
  nand GNAME9981(G9981,G10119,G10120);
  nand GNAME9982(G9982,G10124,G10125);
  nand GNAME9983(G9983,G10129,G10130);
  nand GNAME9984(G9984,G10134,G10135);
  nand GNAME9985(G9985,G10139,G10140);
  nand GNAME9986(G9986,G10024,G10025);
  nand GNAME9987(G9987,G10021,G10022);
  nand GNAME9988(G9988,G10026,G10019);
  and GNAME9989(G9989,G10016,G10014);
  and GNAME9990(G9990,G10027,G10012);
  and GNAME9991(G9991,G10008,G10009);
  nand GNAME9992(G9992,G10005,G10006);
  or GNAME9993(G9993,G10003,G9994);
  nor GNAME9994(G9994,G9941,G9942);
  not GNAME9995(G9995,G36378);
  not GNAME9996(G9996,G36133);
  and GNAME9997(G9997,G10047,G10048);
  nand GNAME9998(G9998,G10039,G10040);
  or GNAME9999(G9999,G10037,G9969);
  not GNAME10000(G10000,G9960);
  not GNAME10001(G10001,G9941);
  or GNAME10002(G10002,G10001,G36396);
  and GNAME10003(G10003,G10002,G36151);
  nand GNAME10004(G10004,G9944,G9943);
  nand GNAME10005(G10005,G9993,G10004);
  or GNAME10006(G10006,G9943,G9944);
  nand GNAME10007(G10007,G9946,G9945);
  nand GNAME10008(G10008,G9992,G10007);
  or GNAME10009(G10009,G9945,G9946);
  not GNAME10010(G10010,G9991);
  or GNAME10011(G10011,G36148,G36393);
  nand GNAME10012(G10012,G10010,G10011);
  not GNAME10013(G10013,G9990);
  nand GNAME10014(G10014,G36147,G36392);
  or GNAME10015(G10015,G36392,G36147);
  nand GNAME10016(G10016,G10013,G10015);
  not GNAME10017(G10017,G9989);
  or GNAME10018(G10018,G36391,G36146);
  nand GNAME10019(G10019,G10017,G10018);
  nand GNAME10020(G10020,G9948,G9947);
  nand GNAME10021(G10021,G9988,G10020);
  or GNAME10022(G10022,G9947,G9948);
  nand GNAME10023(G10023,G9950,G9949);
  nand GNAME10024(G10024,G9987,G10023);
  or GNAME10025(G10025,G9949,G9950);
  nand GNAME10026(G10026,G36146,G36391);
  nand GNAME10027(G10027,G36393,G36148);
  nand GNAME10028(G10028,G36137,G36382);
  and GNAME10029(G10029,G36138,G36383);
  and GNAME10030(G10030,G36142,G36387);
  nand GNAME10031(G10031,G9951,G9952);
  nand GNAME10032(G10032,G9986,G10031);
  or GNAME10033(G10033,G9951,G9952);
  nor GNAME10034(G10034,G36387,G36142);
  nand GNAME10035(G10035,G10147,G9971);
  or GNAME10036(G10036,G36141,G36386);
  and GNAME10037(G10037,G36141,G36386);
  nand GNAME10038(G10038,G9955,G9954);
  nand GNAME10039(G10039,G9999,G10038);
  or GNAME10040(G10040,G9954,G9955);
  nand GNAME10041(G10041,G9957,G9956);
  nand GNAME10042(G10042,G9998,G10041);
  or GNAME10043(G10043,G9956,G9957);
  nor GNAME10044(G10044,G36383,G36138);
  nand GNAME10045(G10045,G10146,G9967);
  or GNAME10046(G10046,G9958,G9959);
  nand GNAME10047(G10047,G10046,G9960);
  nand GNAME10048(G10048,G9958,G9959);
  not GNAME10049(G10049,G9997);
  or GNAME10050(G10050,G9961,G9962);
  nand GNAME10051(G10051,G10049,G10050);
  nand GNAME10052(G10052,G9961,G9962);
  not GNAME10053(G10053,G9963);
  nand GNAME10054(G10054,G9965,G9964);
  nand GNAME10055(G10055,G10054,G9963);
  or GNAME10056(G10056,G9964,G9965);
  nand GNAME10057(G10057,G10113,G10114,G10055,G10056);
  nand GNAME10058(G10058,G10053,G10056);
  nand GNAME10059(G10059,G10115,G10058,G10054);
  or GNAME10060(G10060,G36382,G36137);
  nand GNAME10061(G10061,G10028,G10060);
  nand GNAME10062(G10062,G10061,G10146,G9967);
  nand GNAME10063(G10063,G10028,G9966);
  or GNAME10064(G10064,G10029,G9967);
  or GNAME10065(G10065,G10029,G10044);
  nand GNAME10066(G10066,G10065,G9968);
  nand GNAME10067(G10067,G10141,G10142,G10147,G9971);
  nand GNAME10068(G10068,G36141,G36386);
  nand GNAME10069(G10069,G10068,G9969);
  or GNAME10070(G10070,G10030,G10034);
  nand GNAME10071(G10071,G10070,G9970);
  or GNAME10072(G10072,G10030,G9971);
  nand GNAME10073(G10073,G10018,G10026);
  nand GNAME10074(G10074,G10014,G10015);
  nand GNAME10075(G10075,G10011,G10027);
  nand GNAME10076(G10076,G9942,G10110);
  or GNAME10077(G10077,G36143,G9951);
  or GNAME10078(G10078,G36388,G9952);
  and GNAME10079(G10079,G10077,G10078);
  nand GNAME10080(G10080,G9986,G10077,G10078);
  or GNAME10081(G10081,G10079,G9986);
  or GNAME10082(G10082,G36144,G9950);
  or GNAME10083(G10083,G36389,G9949);
  and GNAME10084(G10084,G10082,G10083);
  nand GNAME10085(G10085,G9987,G10082,G10083);
  or GNAME10086(G10086,G10084,G9987);
  or GNAME10087(G10087,G36145,G9948);
  or GNAME10088(G10088,G36390,G9947);
  and GNAME10089(G10089,G10087,G10088);
  nand GNAME10090(G10090,G9988,G10087,G10088);
  or GNAME10091(G10091,G10089,G9988);
  nand GNAME10092(G10092,G10017,G10073);
  nand GNAME10093(G10093,G9989,G10018,G10026);
  nand GNAME10094(G10094,G10013,G10074);
  nand GNAME10095(G10095,G9990,G10014,G10015);
  nand GNAME10096(G10096,G10010,G10075);
  nand GNAME10097(G10097,G9991,G10011,G10027);
  or GNAME10098(G10098,G36149,G9946);
  or GNAME10099(G10099,G36394,G9945);
  and GNAME10100(G10100,G10098,G10099);
  nand GNAME10101(G10101,G9992,G10098,G10099);
  or GNAME10102(G10102,G10100,G9992);
  or GNAME10103(G10103,G36150,G9944);
  or GNAME10104(G10104,G36395,G9943);
  and GNAME10105(G10105,G10103,G10104);
  nand GNAME10106(G10106,G9993,G10103,G10104);
  or GNAME10107(G10107,G10105,G9993);
  nand GNAME10108(G10108,G9941,G36151);
  or GNAME10109(G10109,G36151,G9941);
  nand GNAME10110(G10110,G10108,G10109);
  or GNAME10111(G10111,G36151,G10001,G9942);
  nand GNAME10112(G10112,G36151,G9994);
  or GNAME10113(G10113,G36133,G9995);
  or GNAME10114(G10114,G36378,G9996);
  nand GNAME10115(G10115,G10113,G10114);
  or GNAME10116(G10116,G36379,G9965);
  or GNAME10117(G10117,G36134,G9964);
  nand GNAME10118(G10118,G10116,G10117);
  nand GNAME10119(G10119,G10053,G10118);
  nand GNAME10120(G10120,G9963,G10116,G10117);
  or GNAME10121(G10121,G36380,G9962);
  or GNAME10122(G10122,G36135,G9961);
  nand GNAME10123(G10123,G10121,G10122);
  nand GNAME10124(G10124,G10049,G10123);
  nand GNAME10125(G10125,G9997,G10121,G10122);
  or GNAME10126(G10126,G36381,G9959);
  or GNAME10127(G10127,G36136,G9958);
  nand GNAME10128(G10128,G10126,G10127);
  nand GNAME10129(G10129,G10000,G10126,G10127);
  nand GNAME10130(G10130,G9960,G10128);
  or GNAME10131(G10131,G36139,G9957);
  or GNAME10132(G10132,G36384,G9956);
  and GNAME10133(G10133,G10131,G10132);
  nand GNAME10134(G10134,G9998,G10131,G10132);
  or GNAME10135(G10135,G10133,G9998);
  or GNAME10136(G10136,G36140,G9955);
  or GNAME10137(G10137,G36385,G9954);
  and GNAME10138(G10138,G10136,G10137);
  nand GNAME10139(G10139,G9999,G10136,G10137);
  or GNAME10140(G10140,G10138,G9999);
  or GNAME10141(G10141,G36141,G9953);
  nand GNAME10142(G10142,G9953,G36141);
  or GNAME10143(G10143,G36397,G9940);
  nand GNAME10144(G10144,G9940,G36397);
  not GNAME10145(G10145,G10028);
  not GNAME10146(G10146,G10029);
  not GNAME10147(G10147,G10030);
  nand GNAME10148(G10148,G10284,G10282);
  nand GNAME10149(G10149,G10285,G10243);
  not GNAME10150(G10150,G36642);
  nor GNAME10151(G10151,G9972,G10150);
  not GNAME10152(G10152,G36641);
  not GNAME10153(G10153,G9980);
  not GNAME10154(G10154,G36640);
  not GNAME10155(G10155,G9979);
  not GNAME10156(G10156,G36639);
  not GNAME10157(G10157,G9978);
  not GNAME10158(G10158,G36638);
  not GNAME10159(G10159,G9977);
  not GNAME10160(G10160,G36637);
  not GNAME10161(G10161,G9976);
  not GNAME10162(G10162,G36636);
  not GNAME10163(G10163,G9975);
  not GNAME10164(G10164,G36635);
  not GNAME10165(G10165,G9974);
  not GNAME10166(G10166,G36634);
  not GNAME10167(G10167,G9973);
  not GNAME10168(G10168,G36633);
  not GNAME10169(G10169,G9934);
  not GNAME10170(G10170,G36632);
  not GNAME10171(G10171,G9935);
  not GNAME10172(G10172,G36631);
  not GNAME10173(G10173,G9985);
  not GNAME10174(G10174,G36630);
  not GNAME10175(G10175,G9984);
  not GNAME10176(G10176,G36629);
  not GNAME10177(G10177,G9936);
  not GNAME10178(G10178,G36628);
  not GNAME10179(G10179,G9937);
  not GNAME10180(G10180,G36627);
  not GNAME10181(G10181,G9983);
  not GNAME10182(G10182,G36626);
  not GNAME10183(G10183,G9982);
  not GNAME10184(G10184,G36625);
  not GNAME10185(G10185,G36624);
  and GNAME10186(G10186,G10279,G10329);
  not GNAME10187(G10187,G9981);
  nand GNAME10188(G10188,G10319,G10320);
  and GNAME10189(G10189,G10286,G10263);
  and GNAME10190(G10190,G10289,G10290);
  and GNAME10191(G10191,G10293,G10294);
  and GNAME10192(G10192,G10297,G10298);
  and GNAME10193(G10193,G10301,G10302);
  and GNAME10194(G10194,G10305,G10306);
  and GNAME10195(G10195,G10309,G10310);
  and GNAME10196(G10196,G10313,G10314);
  and GNAME10197(G10197,G10317,G10318);
  and GNAME10198(G10198,G10324,G10325);
  and GNAME10199(G10199,G10328,G10329);
  and GNAME10200(G10200,G10332,G10333);
  and GNAME10201(G10201,G10336,G10337);
  and GNAME10202(G10202,G10340,G10341);
  and GNAME10203(G10203,G10344,G10345);
  and GNAME10204(G10204,G10348,G10349);
  and GNAME10205(G10205,G10352,G10353);
  and GNAME10206(G10206,G10356,G10357);
  and GNAME10207(G10207,G10260,G10290);
  and GNAME10208(G10208,G10287,G10288);
  and GNAME10209(G10209,G10258,G10294);
  and GNAME10210(G10210,G10291,G10292);
  and GNAME10211(G10211,G10256,G10298);
  and GNAME10212(G10212,G10295,G10296);
  and GNAME10213(G10213,G10254,G10302);
  and GNAME10214(G10214,G10299,G10300);
  and GNAME10215(G10215,G10252,G10306);
  and GNAME10216(G10216,G10303,G10304);
  and GNAME10217(G10217,G10250,G10310);
  and GNAME10218(G10218,G10307,G10308);
  and GNAME10219(G10219,G10248,G10314);
  and GNAME10220(G10220,G10311,G10312);
  and GNAME10221(G10221,G10245,G10246);
  and GNAME10222(G10222,G10315,G10316);
  not GNAME10223(G10223,G9939);
  not GNAME10224(G10224,G9938);
  not GNAME10225(G10225,G36623);
  and GNAME10226(G10226,G10326,G10327);
  and GNAME10227(G10227,G10277,G10333);
  and GNAME10228(G10228,G10330,G10331);
  and GNAME10229(G10229,G10275,G10337);
  and GNAME10230(G10230,G10334,G10335);
  and GNAME10231(G10231,G10273,G10341);
  and GNAME10232(G10232,G10338,G10339);
  and GNAME10233(G10233,G10271,G10345);
  and GNAME10234(G10234,G10342,G10343);
  and GNAME10235(G10235,G10269,G10349);
  and GNAME10236(G10236,G10346,G10347);
  and GNAME10237(G10237,G10267,G10353);
  and GNAME10238(G10238,G10350,G10351);
  and GNAME10239(G10239,G10265,G10357);
  and GNAME10240(G10240,G10354,G10355);
  and GNAME10241(G10241,G10262,G10263);
  and GNAME10242(G10242,G10358,G10359);
  not GNAME10243(G10243,G10151);
  or GNAME10244(G10244,G10151,G36641);
  nand GNAME10245(G10245,G10223,G10244);
  or GNAME10246(G10246,G10243,G10152);
  nor GNAME10247(G10247,G36640,G10153);
  or GNAME10248(G10248,G10221,G10247);
  nor GNAME10249(G10249,G36639,G10155);
  or GNAME10250(G10250,G10219,G10249);
  nor GNAME10251(G10251,G36638,G10157);
  or GNAME10252(G10252,G10217,G10251);
  nor GNAME10253(G10253,G36637,G10159);
  or GNAME10254(G10254,G10215,G10253);
  nor GNAME10255(G10255,G36636,G10161);
  or GNAME10256(G10256,G10213,G10255);
  nor GNAME10257(G10257,G36635,G10163);
  or GNAME10258(G10258,G10211,G10257);
  nor GNAME10259(G10259,G36634,G10165);
  or GNAME10260(G10260,G10209,G10259);
  nor GNAME10261(G10261,G36633,G10167);
  or GNAME10262(G10262,G10207,G10261);
  or GNAME10263(G10263,G9973,G10168);
  nor GNAME10264(G10264,G36632,G10169);
  or GNAME10265(G10265,G10241,G10264);
  nor GNAME10266(G10266,G36631,G10171);
  or GNAME10267(G10267,G10239,G10266);
  nor GNAME10268(G10268,G36630,G10173);
  or GNAME10269(G10269,G10237,G10268);
  nor GNAME10270(G10270,G36629,G10175);
  or GNAME10271(G10271,G10235,G10270);
  nor GNAME10272(G10272,G36628,G10177);
  or GNAME10273(G10273,G10233,G10272);
  nor GNAME10274(G10274,G36627,G10179);
  or GNAME10275(G10275,G10231,G10274);
  nor GNAME10276(G10276,G36626,G10181);
  or GNAME10277(G10277,G10229,G10276);
  nor GNAME10278(G10278,G36625,G10183);
  or GNAME10279(G10279,G10227,G10278);
  nor GNAME10280(G10280,G36624,G10187);
  or GNAME10281(G10281,G10186,G10280);
  nand GNAME10282(G10282,G10323,G10281,G10325);
  nand GNAME10283(G10283,G10325,G10186);
  nand GNAME10284(G10284,G10321,G10322,G10283,G10324);
  nand GNAME10285(G10285,G10150,G9972);
  or GNAME10286(G10286,G36633,G10167);
  nand GNAME10287(G10287,G10189,G10207);
  or GNAME10288(G10288,G10207,G10189);
  or GNAME10289(G10289,G36634,G10165);
  or GNAME10290(G10290,G9974,G10166);
  nand GNAME10291(G10291,G10190,G10209);
  or GNAME10292(G10292,G10209,G10190);
  or GNAME10293(G10293,G36635,G10163);
  or GNAME10294(G10294,G9975,G10164);
  nand GNAME10295(G10295,G10191,G10211);
  or GNAME10296(G10296,G10211,G10191);
  or GNAME10297(G10297,G36636,G10161);
  or GNAME10298(G10298,G9976,G10162);
  nand GNAME10299(G10299,G10192,G10213);
  or GNAME10300(G10300,G10213,G10192);
  or GNAME10301(G10301,G36637,G10159);
  or GNAME10302(G10302,G9977,G10160);
  nand GNAME10303(G10303,G10193,G10215);
  or GNAME10304(G10304,G10215,G10193);
  or GNAME10305(G10305,G36638,G10157);
  or GNAME10306(G10306,G9978,G10158);
  nand GNAME10307(G10307,G10194,G10217);
  or GNAME10308(G10308,G10217,G10194);
  or GNAME10309(G10309,G36639,G10155);
  or GNAME10310(G10310,G9979,G10156);
  nand GNAME10311(G10311,G10195,G10219);
  or GNAME10312(G10312,G10219,G10195);
  or GNAME10313(G10313,G36640,G10153);
  or GNAME10314(G10314,G9980,G10154);
  nand GNAME10315(G10315,G10196,G10221);
  or GNAME10316(G10316,G10221,G10196);
  or GNAME10317(G10317,G36641,G10223);
  or GNAME10318(G10318,G9939,G10152);
  nand GNAME10319(G10319,G10151,G10197);
  or GNAME10320(G10320,G10151,G10197);
  or GNAME10321(G10321,G36623,G10224);
  or GNAME10322(G10322,G9938,G10225);
  nand GNAME10323(G10323,G10321,G10322);
  or GNAME10324(G10324,G36624,G10187);
  or GNAME10325(G10325,G9981,G10185);
  nand GNAME10326(G10326,G10186,G10198);
  or GNAME10327(G10327,G10186,G10198);
  or GNAME10328(G10328,G36625,G10183);
  or GNAME10329(G10329,G9982,G10184);
  nand GNAME10330(G10330,G10199,G10227);
  or GNAME10331(G10331,G10227,G10199);
  or GNAME10332(G10332,G36626,G10181);
  or GNAME10333(G10333,G9983,G10182);
  nand GNAME10334(G10334,G10200,G10229);
  or GNAME10335(G10335,G10229,G10200);
  or GNAME10336(G10336,G36627,G10179);
  or GNAME10337(G10337,G9937,G10180);
  nand GNAME10338(G10338,G10201,G10231);
  or GNAME10339(G10339,G10231,G10201);
  or GNAME10340(G10340,G36628,G10177);
  or GNAME10341(G10341,G9936,G10178);
  nand GNAME10342(G10342,G10202,G10233);
  or GNAME10343(G10343,G10233,G10202);
  or GNAME10344(G10344,G36629,G10175);
  or GNAME10345(G10345,G9984,G10176);
  nand GNAME10346(G10346,G10203,G10235);
  or GNAME10347(G10347,G10235,G10203);
  or GNAME10348(G10348,G36630,G10173);
  or GNAME10349(G10349,G9985,G10174);
  nand GNAME10350(G10350,G10204,G10237);
  or GNAME10351(G10351,G10237,G10204);
  or GNAME10352(G10352,G36631,G10171);
  or GNAME10353(G10353,G9935,G10172);
  nand GNAME10354(G10354,G10205,G10239);
  or GNAME10355(G10355,G10239,G10205);
  or GNAME10356(G10356,G36632,G10169);
  or GNAME10357(G10357,G9934,G10170);
  nand GNAME10358(G10358,G10206,G10241);
  or GNAME10359(G10359,G10241,G10206);
  not GNAME10360(G10360,G36378);
  and GNAME10361(G10361,G10585,G10586);
  and GNAME10362(G10362,G10581,G10583);
  and GNAME10363(G10363,G10579,G10580);
  and GNAME10364(G10364,G10575,G10577);
  and GNAME10365(G10365,G10573,G10574);
  and GNAME10366(G10366,G10568,G10570);
  nand GNAME10367(G10367,G10590,G10678,G10679);
  not GNAME10368(G10368,G921);
  nand GNAME10369(G10369,G32,G921);
  not GNAME10370(G10370,G31);
  not GNAME10371(G10371,G909);
  not GNAME10372(G10372,G30);
  not GNAME10373(G10373,G898);
  not GNAME10374(G10374,G29);
  not GNAME10375(G10375,G892);
  not GNAME10376(G10376,G25);
  not GNAME10377(G10377,G891);
  not GNAME10378(G10378,G24);
  not GNAME10379(G10379,G23);
  not GNAME10380(G10380,G890);
  not GNAME10381(G10381,G17);
  not GNAME10382(G10382,G21);
  not GNAME10383(G10383,G917);
  not GNAME10384(G10384,G20);
  not GNAME10385(G10385,G916);
  not GNAME10386(G10386,G19);
  not GNAME10387(G10387,G913);
  not GNAME10388(G10388,G16);
  not GNAME10389(G10389,G912);
  not GNAME10390(G10390,G15);
  not GNAME10391(G10391,G911);
  not GNAME10392(G10392,G14);
  not GNAME10393(G10393,G910);
  not GNAME10394(G10394,G13);
  not GNAME10395(G10395,G908);
  not GNAME10396(G10396,G12);
  not GNAME10397(G10397,G907);
  not GNAME10398(G10398,G11);
  not GNAME10399(G10399,G906);
  not GNAME10400(G10400,G10);
  not GNAME10401(G10401,G905);
  not GNAME10402(G10402,G9);
  not GNAME10403(G10403,G904);
  not GNAME10404(G10404,G8);
  not GNAME10405(G10405,G903);
  not GNAME10406(G10406,G7);
  not GNAME10407(G10407,G902);
  not GNAME10408(G10408,G6);
  not GNAME10409(G10409,G4);
  not GNAME10410(G10410,G900);
  nor GNAME10411(G10411,G10716,G10418);
  not GNAME10412(G10412,G3);
  not GNAME10413(G10413,G899);
  and GNAME10414(G10414,G10562,G10563);
  not GNAME10415(G10415,G2);
  not GNAME10416(G10416,G897);
  and GNAME10417(G10417,G10554,G10555);
  nor GNAME10418(G10418,G10556,G10417);
  and GNAME10419(G10419,G10520,G10521);
  and GNAME10420(G10420,G10517,G10518);
  or GNAME10421(G10421,G10519,G10420);
  and GNAME10422(G10422,G10510,G10511);
  and GNAME10423(G10423,G10507,G10508);
  or GNAME10424(G10424,G10509,G10423);
  nand GNAME10425(G10425,G10714,G10715);
  nand GNAME10426(G10426,G10594,G10595);
  nand GNAME10427(G10427,G10599,G10600);
  nand GNAME10428(G10428,G10604,G10605);
  nand GNAME10429(G10429,G10606,G10607);
  nand GNAME10430(G10430,G10608,G10609);
  nand GNAME10431(G10431,G10610,G10611);
  nand GNAME10432(G10432,G10615,G10616);
  nand GNAME10433(G10433,G10623,G10624);
  nand GNAME10434(G10434,G10628,G10629);
  nand GNAME10435(G10435,G10633,G10634);
  nand GNAME10436(G10436,G10638,G10639);
  nand GNAME10437(G10437,G10643,G10644);
  nand GNAME10438(G10438,G10648,G10649);
  nand GNAME10439(G10439,G10653,G10654);
  nand GNAME10440(G10440,G10658,G10659);
  nand GNAME10441(G10441,G10663,G10664);
  nand GNAME10442(G10442,G10668,G10669);
  nand GNAME10443(G10443,G10673,G10674);
  nand GNAME10444(G10444,G10683,G10684);
  nand GNAME10445(G10445,G10688,G10689);
  nand GNAME10446(G10446,G10693,G10694);
  nand GNAME10447(G10447,G10698,G10699);
  nand GNAME10448(G10448,G10705,G10706);
  nand GNAME10449(G10449,G10710,G10711);
  nand GNAME10450(G10450,G10499,G10500);
  nand GNAME10451(G10451,G10496,G10497);
  nand GNAME10452(G10452,G10501,G10494);
  and GNAME10453(G10453,G10491,G10489);
  and GNAME10454(G10454,G10502,G10487);
  and GNAME10455(G10455,G10483,G10484);
  nand GNAME10456(G10456,G10480,G10481);
  not GNAME10457(G10457,G1);
  not GNAME10458(G10458,G896);
  or GNAME10459(G10459,G10478,G10468);
  and GNAME10460(G10460,G10558,G10559);
  nand GNAME10461(G10461,G10551,G10552);
  nand GNAME10462(G10462,G10548,G10549);
  nand GNAME10463(G10463,G10545,G10546);
  nand GNAME10464(G10464,G10542,G10543);
  nand GNAME10465(G10465,G10539,G10540);
  nand GNAME10466(G10466,G10536,G10537);
  nand GNAME10467(G10467,G10533,G10534);
  nor GNAME10468(G10468,G10369,G10370);
  nand GNAME10469(G10469,G10530,G10531);
  nand GNAME10470(G10470,G10527,G10528);
  nand GNAME10471(G10471,G10524,G10525);
  or GNAME10472(G10472,G10522,G10419);
  nand GNAME10473(G10473,G10514,G10515);
  or GNAME10474(G10474,G10512,G10422);
  not GNAME10475(G10475,G10411);
  not GNAME10476(G10476,G10369);
  or GNAME10477(G10477,G10476,G31);
  and GNAME10478(G10478,G10477,G920);
  nand GNAME10479(G10479,G10372,G10371);
  nand GNAME10480(G10480,G10459,G10479);
  or GNAME10481(G10481,G10371,G10372);
  nand GNAME10482(G10482,G10374,G10373);
  nand GNAME10483(G10483,G10456,G10482);
  or GNAME10484(G10484,G10373,G10374);
  not GNAME10485(G10485,G10455);
  or GNAME10486(G10486,G895,G28);
  nand GNAME10487(G10487,G10485,G10486);
  not GNAME10488(G10488,G10454);
  nand GNAME10489(G10489,G894,G27);
  or GNAME10490(G10490,G27,G894);
  nand GNAME10491(G10491,G10488,G10490);
  not GNAME10492(G10492,G10453);
  or GNAME10493(G10493,G26,G893);
  nand GNAME10494(G10494,G10492,G10493);
  nand GNAME10495(G10495,G10376,G10375);
  nand GNAME10496(G10496,G10452,G10495);
  or GNAME10497(G10497,G10375,G10376);
  nand GNAME10498(G10498,G10378,G10377);
  nand GNAME10499(G10499,G10451,G10498);
  or GNAME10500(G10500,G10377,G10378);
  nand GNAME10501(G10501,G893,G26);
  nand GNAME10502(G10502,G28,G895);
  nand GNAME10503(G10503,G901,G5);
  and GNAME10504(G10504,G915,G18);
  and GNAME10505(G10505,G919,G22);
  nand GNAME10506(G10506,G10379,G10380);
  nand GNAME10507(G10507,G10450,G10506);
  or GNAME10508(G10508,G10379,G10380);
  nor GNAME10509(G10509,G22,G919);
  nand GNAME10510(G10510,G10718,G10424);
  or GNAME10511(G10511,G918,G21);
  and GNAME10512(G10512,G918,G21);
  nand GNAME10513(G10513,G10384,G10383);
  nand GNAME10514(G10514,G10474,G10513);
  or GNAME10515(G10515,G10383,G10384);
  nand GNAME10516(G10516,G10386,G10385);
  nand GNAME10517(G10517,G10473,G10516);
  or GNAME10518(G10518,G10385,G10386);
  nor GNAME10519(G10519,G18,G915);
  nand GNAME10520(G10520,G10717,G10421);
  or GNAME10521(G10521,G914,G17);
  and GNAME10522(G10522,G914,G17);
  nand GNAME10523(G10523,G10388,G10387);
  nand GNAME10524(G10524,G10472,G10523);
  or GNAME10525(G10525,G10387,G10388);
  nand GNAME10526(G10526,G10390,G10389);
  nand GNAME10527(G10527,G10471,G10526);
  or GNAME10528(G10528,G10389,G10390);
  nand GNAME10529(G10529,G10392,G10391);
  nand GNAME10530(G10530,G10470,G10529);
  or GNAME10531(G10531,G10391,G10392);
  nand GNAME10532(G10532,G10394,G10393);
  nand GNAME10533(G10533,G10469,G10532);
  or GNAME10534(G10534,G10393,G10394);
  nand GNAME10535(G10535,G10396,G10395);
  nand GNAME10536(G10536,G10467,G10535);
  or GNAME10537(G10537,G10395,G10396);
  nand GNAME10538(G10538,G10398,G10397);
  nand GNAME10539(G10539,G10466,G10538);
  or GNAME10540(G10540,G10397,G10398);
  nand GNAME10541(G10541,G10400,G10399);
  nand GNAME10542(G10542,G10465,G10541);
  or GNAME10543(G10543,G10399,G10400);
  nand GNAME10544(G10544,G10402,G10401);
  nand GNAME10545(G10545,G10464,G10544);
  or GNAME10546(G10546,G10401,G10402);
  nand GNAME10547(G10547,G10404,G10403);
  nand GNAME10548(G10548,G10463,G10547);
  or GNAME10549(G10549,G10403,G10404);
  nand GNAME10550(G10550,G10406,G10405);
  nand GNAME10551(G10551,G10462,G10550);
  or GNAME10552(G10552,G10405,G10406);
  nand GNAME10553(G10553,G10408,G10407);
  nand GNAME10554(G10554,G10461,G10553);
  or GNAME10555(G10555,G10407,G10408);
  nor GNAME10556(G10556,G901,G5);
  or GNAME10557(G10557,G10409,G10410);
  nand GNAME10558(G10558,G10557,G10411);
  nand GNAME10559(G10559,G10409,G10410);
  not GNAME10560(G10560,G10460);
  or GNAME10561(G10561,G10412,G10413);
  nand GNAME10562(G10562,G10560,G10561);
  nand GNAME10563(G10563,G10412,G10413);
  not GNAME10564(G10564,G10414);
  nand GNAME10565(G10565,G10416,G10415);
  nand GNAME10566(G10566,G10565,G10414);
  or GNAME10567(G10567,G10415,G10416);
  nand GNAME10568(G10568,G10617,G10618,G10566,G10567);
  nand GNAME10569(G10569,G10564,G10567);
  nand GNAME10570(G10570,G10619,G10569,G10565);
  or GNAME10571(G10571,G5,G901);
  nand GNAME10572(G10572,G10503,G10571);
  nand GNAME10573(G10573,G10572,G10417);
  nand GNAME10574(G10574,G10503,G10418);
  nand GNAME10575(G10575,G10700,G10701,G10717,G10421);
  nand GNAME10576(G10576,G914,G17);
  nand GNAME10577(G10577,G10576,G10419);
  or GNAME10578(G10578,G10504,G10519);
  nand GNAME10579(G10579,G10578,G10420);
  or GNAME10580(G10580,G10504,G10421);
  nand GNAME10581(G10581,G10712,G10713,G10718,G10424);
  nand GNAME10582(G10582,G918,G21);
  nand GNAME10583(G10583,G10582,G10422);
  or GNAME10584(G10584,G10505,G10509);
  nand GNAME10585(G10585,G10584,G10423);
  or GNAME10586(G10586,G10505,G10424);
  nand GNAME10587(G10587,G10493,G10501);
  nand GNAME10588(G10588,G10489,G10490);
  nand GNAME10589(G10589,G10486,G10502);
  nand GNAME10590(G10590,G10370,G10677);
  or GNAME10591(G10591,G890,G10379);
  or GNAME10592(G10592,G23,G10380);
  and GNAME10593(G10593,G10591,G10592);
  nand GNAME10594(G10594,G10450,G10591,G10592);
  or GNAME10595(G10595,G10593,G10450);
  or GNAME10596(G10596,G891,G10378);
  or GNAME10597(G10597,G24,G10377);
  and GNAME10598(G10598,G10596,G10597);
  nand GNAME10599(G10599,G10451,G10596,G10597);
  or GNAME10600(G10600,G10598,G10451);
  or GNAME10601(G10601,G892,G10376);
  or GNAME10602(G10602,G25,G10375);
  and GNAME10603(G10603,G10601,G10602);
  nand GNAME10604(G10604,G10452,G10601,G10602);
  or GNAME10605(G10605,G10603,G10452);
  nand GNAME10606(G10606,G10492,G10587);
  nand GNAME10607(G10607,G10453,G10493,G10501);
  nand GNAME10608(G10608,G10488,G10588);
  nand GNAME10609(G10609,G10454,G10489,G10490);
  nand GNAME10610(G10610,G10485,G10589);
  nand GNAME10611(G10611,G10455,G10486,G10502);
  or GNAME10612(G10612,G898,G10374);
  or GNAME10613(G10613,G29,G10373);
  and GNAME10614(G10614,G10612,G10613);
  nand GNAME10615(G10615,G10456,G10612,G10613);
  or GNAME10616(G10616,G10614,G10456);
  or GNAME10617(G10617,G896,G10457);
  or GNAME10618(G10618,G1,G10458);
  nand GNAME10619(G10619,G10617,G10618);
  or GNAME10620(G10620,G2,G10416);
  or GNAME10621(G10621,G897,G10415);
  nand GNAME10622(G10622,G10620,G10621);
  nand GNAME10623(G10623,G10564,G10622);
  nand GNAME10624(G10624,G10414,G10620,G10621);
  or GNAME10625(G10625,G909,G10372);
  or GNAME10626(G10626,G30,G10371);
  and GNAME10627(G10627,G10625,G10626);
  nand GNAME10628(G10628,G10459,G10625,G10626);
  or GNAME10629(G10629,G10627,G10459);
  or GNAME10630(G10630,G3,G10413);
  or GNAME10631(G10631,G899,G10412);
  nand GNAME10632(G10632,G10630,G10631);
  nand GNAME10633(G10633,G10560,G10632);
  nand GNAME10634(G10634,G10460,G10630,G10631);
  or GNAME10635(G10635,G4,G10410);
  or GNAME10636(G10636,G900,G10409);
  nand GNAME10637(G10637,G10635,G10636);
  nand GNAME10638(G10638,G10475,G10635,G10636);
  nand GNAME10639(G10639,G10411,G10637);
  or GNAME10640(G10640,G902,G10408);
  or GNAME10641(G10641,G6,G10407);
  and GNAME10642(G10642,G10640,G10641);
  nand GNAME10643(G10643,G10461,G10640,G10641);
  or GNAME10644(G10644,G10642,G10461);
  or GNAME10645(G10645,G903,G10406);
  or GNAME10646(G10646,G7,G10405);
  and GNAME10647(G10647,G10645,G10646);
  nand GNAME10648(G10648,G10462,G10645,G10646);
  or GNAME10649(G10649,G10647,G10462);
  or GNAME10650(G10650,G904,G10404);
  or GNAME10651(G10651,G8,G10403);
  and GNAME10652(G10652,G10650,G10651);
  nand GNAME10653(G10653,G10463,G10650,G10651);
  or GNAME10654(G10654,G10652,G10463);
  or GNAME10655(G10655,G905,G10402);
  or GNAME10656(G10656,G9,G10401);
  and GNAME10657(G10657,G10655,G10656);
  nand GNAME10658(G10658,G10464,G10655,G10656);
  or GNAME10659(G10659,G10657,G10464);
  or GNAME10660(G10660,G906,G10400);
  or GNAME10661(G10661,G10,G10399);
  and GNAME10662(G10662,G10660,G10661);
  nand GNAME10663(G10663,G10465,G10660,G10661);
  or GNAME10664(G10664,G10662,G10465);
  or GNAME10665(G10665,G907,G10398);
  or GNAME10666(G10666,G11,G10397);
  and GNAME10667(G10667,G10665,G10666);
  nand GNAME10668(G10668,G10466,G10665,G10666);
  or GNAME10669(G10669,G10667,G10466);
  or GNAME10670(G10670,G908,G10396);
  or GNAME10671(G10671,G12,G10395);
  and GNAME10672(G10672,G10670,G10671);
  nand GNAME10673(G10673,G10467,G10670,G10671);
  or GNAME10674(G10674,G10672,G10467);
  nand GNAME10675(G10675,G10369,G920);
  or GNAME10676(G10676,G920,G10369);
  nand GNAME10677(G10677,G10675,G10676);
  or GNAME10678(G10678,G920,G10476,G10370);
  nand GNAME10679(G10679,G920,G10468);
  or GNAME10680(G10680,G910,G10394);
  or GNAME10681(G10681,G13,G10393);
  and GNAME10682(G10682,G10680,G10681);
  nand GNAME10683(G10683,G10469,G10680,G10681);
  or GNAME10684(G10684,G10682,G10469);
  or GNAME10685(G10685,G911,G10392);
  or GNAME10686(G10686,G14,G10391);
  and GNAME10687(G10687,G10685,G10686);
  nand GNAME10688(G10688,G10470,G10685,G10686);
  or GNAME10689(G10689,G10687,G10470);
  or GNAME10690(G10690,G912,G10390);
  or GNAME10691(G10691,G15,G10389);
  and GNAME10692(G10692,G10690,G10691);
  nand GNAME10693(G10693,G10471,G10690,G10691);
  or GNAME10694(G10694,G10692,G10471);
  or GNAME10695(G10695,G913,G10388);
  or GNAME10696(G10696,G16,G10387);
  and GNAME10697(G10697,G10695,G10696);
  nand GNAME10698(G10698,G10472,G10695,G10696);
  or GNAME10699(G10699,G10697,G10472);
  or GNAME10700(G10700,G914,G10381);
  nand GNAME10701(G10701,G10381,G914);
  or GNAME10702(G10702,G916,G10386);
  or GNAME10703(G10703,G19,G10385);
  and GNAME10704(G10704,G10702,G10703);
  nand GNAME10705(G10705,G10473,G10702,G10703);
  or GNAME10706(G10706,G10704,G10473);
  or GNAME10707(G10707,G917,G10384);
  or GNAME10708(G10708,G20,G10383);
  and GNAME10709(G10709,G10707,G10708);
  nand GNAME10710(G10710,G10474,G10707,G10708);
  or GNAME10711(G10711,G10709,G10474);
  or GNAME10712(G10712,G918,G10382);
  nand GNAME10713(G10713,G10382,G918);
  or GNAME10714(G10714,G32,G10368);
  nand GNAME10715(G10715,G10368,G32);
  not GNAME10716(G10716,G10503);
  not GNAME10717(G10717,G10504);
  not GNAME10718(G10718,G10505);
  nand GNAME10719(G10719,G10939,G10937);
  nand GNAME10720(G10720,G10940,G10874);
  not GNAME10721(G10721,G36398);
  nor GNAME10722(G10722,G36153,G10721);
  not GNAME10723(G10723,G36399);
  not GNAME10724(G10724,G36155);
  not GNAME10725(G10725,G36400);
  not GNAME10726(G10726,G36156);
  not GNAME10727(G10727,G36401);
  not GNAME10728(G10728,G36157);
  not GNAME10729(G10729,G36402);
  not GNAME10730(G10730,G36158);
  not GNAME10731(G10731,G36403);
  not GNAME10732(G10732,G36159);
  not GNAME10733(G10733,G36404);
  not GNAME10734(G10734,G36160);
  not GNAME10735(G10735,G36405);
  not GNAME10736(G10736,G36161);
  not GNAME10737(G10737,G36406);
  not GNAME10738(G10738,G36162);
  not GNAME10739(G10739,G36407);
  not GNAME10740(G10740,G36163);
  not GNAME10741(G10741,G36408);
  not GNAME10742(G10742,G36164);
  not GNAME10743(G10743,G36409);
  not GNAME10744(G10744,G36165);
  not GNAME10745(G10745,G36410);
  not GNAME10746(G10746,G36166);
  not GNAME10747(G10747,G36411);
  not GNAME10748(G10748,G36167);
  not GNAME10749(G10749,G36412);
  not GNAME10750(G10750,G36168);
  not GNAME10751(G10751,G36413);
  not GNAME10752(G10752,G36169);
  not GNAME10753(G10753,G36414);
  not GNAME10754(G10754,G36170);
  not GNAME10755(G10755,G36415);
  not GNAME10756(G10756,G36171);
  not GNAME10757(G10757,G36416);
  not GNAME10758(G10758,G36172);
  not GNAME10759(G10759,G36417);
  not GNAME10760(G10760,G36173);
  not GNAME10761(G10761,G36418);
  not GNAME10762(G10762,G36174);
  not GNAME10763(G10763,G36419);
  not GNAME10764(G10764,G36175);
  not GNAME10765(G10765,G36420);
  not GNAME10766(G10766,G36176);
  not GNAME10767(G10767,G36421);
  not GNAME10768(G10768,G36177);
  not GNAME10769(G10769,G36422);
  not GNAME10770(G10770,G36178);
  not GNAME10771(G10771,G36423);
  not GNAME10772(G10772,G36179);
  not GNAME10773(G10773,G36424);
  not GNAME10774(G10774,G36180);
  not GNAME10775(G10775,G36425);
  not GNAME10776(G10776,G36181);
  not GNAME10777(G10777,G36426);
  not GNAME10778(G10778,G36182);
  not GNAME10779(G10779,G36427);
  not GNAME10780(G10780,G36428);
  and GNAME10781(G10781,G10934,G10980);
  not GNAME10782(G10782,G36183);
  nand GNAME10783(G10783,G11021,G11022);
  and GNAME10784(G10784,G10941,G10894);
  and GNAME10785(G10785,G10944,G10945);
  and GNAME10786(G10786,G10948,G10949);
  and GNAME10787(G10787,G10952,G10953);
  and GNAME10788(G10788,G10956,G10957);
  and GNAME10789(G10789,G10960,G10961);
  and GNAME10790(G10790,G10964,G10965);
  and GNAME10791(G10791,G10971,G10972);
  and GNAME10792(G10792,G10975,G10976);
  and GNAME10793(G10793,G10979,G10980);
  and GNAME10794(G10794,G10983,G10984);
  and GNAME10795(G10795,G10987,G10988);
  and GNAME10796(G10796,G10991,G10992);
  and GNAME10797(G10797,G10995,G10996);
  and GNAME10798(G10798,G10999,G11000);
  and GNAME10799(G10799,G11003,G11004);
  and GNAME10800(G10800,G11007,G11008);
  and GNAME10801(G10801,G11011,G11012);
  and GNAME10802(G10802,G11015,G11016);
  and GNAME10803(G10803,G11019,G11020);
  and GNAME10804(G10804,G11023,G11024);
  and GNAME10805(G10805,G11027,G11028);
  and GNAME10806(G10806,G11031,G11032);
  and GNAME10807(G10807,G11035,G11036);
  and GNAME10808(G10808,G11039,G11040);
  and GNAME10809(G10809,G11043,G11044);
  and GNAME10810(G10810,G11047,G11048);
  and GNAME10811(G10811,G11051,G11052);
  and GNAME10812(G10812,G11055,G11056);
  and GNAME10813(G10813,G11059,G11060);
  and GNAME10814(G10814,G10891,G10945);
  and GNAME10815(G10815,G10942,G10943);
  and GNAME10816(G10816,G10889,G10949);
  and GNAME10817(G10817,G10946,G10947);
  and GNAME10818(G10818,G10887,G10953);
  and GNAME10819(G10819,G10950,G10951);
  and GNAME10820(G10820,G10885,G10957);
  and GNAME10821(G10821,G10954,G10955);
  and GNAME10822(G10822,G10883,G10961);
  and GNAME10823(G10823,G10958,G10959);
  and GNAME10824(G10824,G10881,G10965);
  and GNAME10825(G10825,G10962,G10963);
  and GNAME10826(G10826,G10879,G10976);
  and GNAME10827(G10827,G10966,G10967);
  not GNAME10828(G10828,G36184);
  not GNAME10829(G10829,G36429);
  and GNAME10830(G10830,G10973,G10974);
  and GNAME10831(G10831,G10876,G10877);
  and GNAME10832(G10832,G10977,G10978);
  and GNAME10833(G10833,G10932,G10984);
  and GNAME10834(G10834,G10981,G10982);
  and GNAME10835(G10835,G10930,G10988);
  and GNAME10836(G10836,G10985,G10986);
  and GNAME10837(G10837,G10928,G10992);
  and GNAME10838(G10838,G10989,G10990);
  and GNAME10839(G10839,G10926,G10996);
  and GNAME10840(G10840,G10993,G10994);
  and GNAME10841(G10841,G10924,G11000);
  and GNAME10842(G10842,G10997,G10998);
  and GNAME10843(G10843,G10922,G11004);
  and GNAME10844(G10844,G11001,G11002);
  and GNAME10845(G10845,G10920,G11008);
  and GNAME10846(G10846,G11005,G11006);
  and GNAME10847(G10847,G10918,G11012);
  and GNAME10848(G10848,G11009,G11010);
  and GNAME10849(G10849,G10916,G11016);
  and GNAME10850(G10850,G11013,G11014);
  and GNAME10851(G10851,G10914,G11024);
  and GNAME10852(G10852,G11017,G11018);
  not GNAME10853(G10853,G36154);
  and GNAME10854(G10854,G10912,G11028);
  and GNAME10855(G10855,G11025,G11026);
  and GNAME10856(G10856,G10910,G11032);
  and GNAME10857(G10857,G11029,G11030);
  and GNAME10858(G10858,G10908,G11036);
  and GNAME10859(G10859,G11033,G11034);
  and GNAME10860(G10860,G10906,G11040);
  and GNAME10861(G10861,G11037,G11038);
  and GNAME10862(G10862,G10904,G11044);
  and GNAME10863(G10863,G11041,G11042);
  and GNAME10864(G10864,G10902,G11048);
  and GNAME10865(G10865,G11045,G11046);
  and GNAME10866(G10866,G10900,G11052);
  and GNAME10867(G10867,G11049,G11050);
  and GNAME10868(G10868,G10898,G11056);
  and GNAME10869(G10869,G11053,G11054);
  and GNAME10870(G10870,G10896,G11060);
  and GNAME10871(G10871,G11057,G11058);
  and GNAME10872(G10872,G10893,G10894);
  and GNAME10873(G10873,G11061,G11062);
  not GNAME10874(G10874,G10722);
  or GNAME10875(G10875,G10722,G36399);
  nand GNAME10876(G10876,G10853,G10875);
  or GNAME10877(G10877,G10874,G10723);
  nor GNAME10878(G10878,G36400,G10724);
  or GNAME10879(G10879,G10831,G10878);
  nor GNAME10880(G10880,G36401,G10726);
  or GNAME10881(G10881,G10826,G10880);
  nor GNAME10882(G10882,G36402,G10728);
  or GNAME10883(G10883,G10824,G10882);
  nor GNAME10884(G10884,G36403,G10730);
  or GNAME10885(G10885,G10822,G10884);
  nor GNAME10886(G10886,G36404,G10732);
  or GNAME10887(G10887,G10820,G10886);
  nor GNAME10888(G10888,G36405,G10734);
  or GNAME10889(G10889,G10818,G10888);
  nor GNAME10890(G10890,G36406,G10736);
  or GNAME10891(G10891,G10816,G10890);
  nor GNAME10892(G10892,G36407,G10738);
  or GNAME10893(G10893,G10814,G10892);
  or GNAME10894(G10894,G36162,G10739);
  nor GNAME10895(G10895,G36408,G10740);
  or GNAME10896(G10896,G10872,G10895);
  nor GNAME10897(G10897,G36409,G10742);
  or GNAME10898(G10898,G10870,G10897);
  nor GNAME10899(G10899,G36410,G10744);
  or GNAME10900(G10900,G10868,G10899);
  nor GNAME10901(G10901,G36411,G10746);
  or GNAME10902(G10902,G10866,G10901);
  nor GNAME10903(G10903,G36412,G10748);
  or GNAME10904(G10904,G10864,G10903);
  nor GNAME10905(G10905,G36413,G10750);
  or GNAME10906(G10906,G10862,G10905);
  nor GNAME10907(G10907,G36414,G10752);
  or GNAME10908(G10908,G10860,G10907);
  nor GNAME10909(G10909,G36415,G10754);
  or GNAME10910(G10910,G10858,G10909);
  nor GNAME10911(G10911,G36416,G10756);
  or GNAME10912(G10912,G10856,G10911);
  nor GNAME10913(G10913,G36417,G10758);
  or GNAME10914(G10914,G10854,G10913);
  nor GNAME10915(G10915,G36418,G10760);
  or GNAME10916(G10916,G10851,G10915);
  nor GNAME10917(G10917,G36419,G10762);
  or GNAME10918(G10918,G10849,G10917);
  nor GNAME10919(G10919,G36420,G10764);
  or GNAME10920(G10920,G10847,G10919);
  nor GNAME10921(G10921,G36421,G10766);
  or GNAME10922(G10922,G10845,G10921);
  nor GNAME10923(G10923,G36422,G10768);
  or GNAME10924(G10924,G10843,G10923);
  nor GNAME10925(G10925,G36423,G10770);
  or GNAME10926(G10926,G10841,G10925);
  nor GNAME10927(G10927,G36424,G10772);
  or GNAME10928(G10928,G10839,G10927);
  nor GNAME10929(G10929,G36425,G10774);
  or GNAME10930(G10930,G10837,G10929);
  nor GNAME10931(G10931,G36426,G10776);
  or GNAME10932(G10932,G10835,G10931);
  nor GNAME10933(G10933,G36427,G10778);
  or GNAME10934(G10934,G10833,G10933);
  nor GNAME10935(G10935,G36428,G10782);
  or GNAME10936(G10936,G10781,G10935);
  nand GNAME10937(G10937,G10970,G10936,G10972);
  nand GNAME10938(G10938,G10972,G10781);
  nand GNAME10939(G10939,G10968,G10969,G10938,G10971);
  nand GNAME10940(G10940,G10721,G36153);
  or GNAME10941(G10941,G36407,G10738);
  nand GNAME10942(G10942,G10784,G10814);
  or GNAME10943(G10943,G10814,G10784);
  or GNAME10944(G10944,G36406,G10736);
  or GNAME10945(G10945,G36161,G10737);
  nand GNAME10946(G10946,G10785,G10816);
  or GNAME10947(G10947,G10816,G10785);
  or GNAME10948(G10948,G36405,G10734);
  or GNAME10949(G10949,G36160,G10735);
  nand GNAME10950(G10950,G10786,G10818);
  or GNAME10951(G10951,G10818,G10786);
  or GNAME10952(G10952,G36404,G10732);
  or GNAME10953(G10953,G36159,G10733);
  nand GNAME10954(G10954,G10787,G10820);
  or GNAME10955(G10955,G10820,G10787);
  or GNAME10956(G10956,G36403,G10730);
  or GNAME10957(G10957,G36158,G10731);
  nand GNAME10958(G10958,G10788,G10822);
  or GNAME10959(G10959,G10822,G10788);
  or GNAME10960(G10960,G36402,G10728);
  or GNAME10961(G10961,G36157,G10729);
  nand GNAME10962(G10962,G10789,G10824);
  or GNAME10963(G10963,G10824,G10789);
  or GNAME10964(G10964,G36401,G10726);
  or GNAME10965(G10965,G36156,G10727);
  nand GNAME10966(G10966,G10790,G10826);
  or GNAME10967(G10967,G10826,G10790);
  or GNAME10968(G10968,G36429,G10828);
  or GNAME10969(G10969,G36184,G10829);
  nand GNAME10970(G10970,G10968,G10969);
  or GNAME10971(G10971,G36428,G10782);
  or GNAME10972(G10972,G36183,G10780);
  nand GNAME10973(G10973,G10781,G10791);
  or GNAME10974(G10974,G10781,G10791);
  or GNAME10975(G10975,G36400,G10724);
  or GNAME10976(G10976,G36155,G10725);
  nand GNAME10977(G10977,G10792,G10831);
  or GNAME10978(G10978,G10831,G10792);
  or GNAME10979(G10979,G36427,G10778);
  or GNAME10980(G10980,G36182,G10779);
  nand GNAME10981(G10981,G10793,G10833);
  or GNAME10982(G10982,G10833,G10793);
  or GNAME10983(G10983,G36426,G10776);
  or GNAME10984(G10984,G36181,G10777);
  nand GNAME10985(G10985,G10794,G10835);
  or GNAME10986(G10986,G10835,G10794);
  or GNAME10987(G10987,G36425,G10774);
  or GNAME10988(G10988,G36180,G10775);
  nand GNAME10989(G10989,G10795,G10837);
  or GNAME10990(G10990,G10837,G10795);
  or GNAME10991(G10991,G36424,G10772);
  or GNAME10992(G10992,G36179,G10773);
  nand GNAME10993(G10993,G10796,G10839);
  or GNAME10994(G10994,G10839,G10796);
  or GNAME10995(G10995,G36423,G10770);
  or GNAME10996(G10996,G36178,G10771);
  nand GNAME10997(G10997,G10797,G10841);
  or GNAME10998(G10998,G10841,G10797);
  or GNAME10999(G10999,G36422,G10768);
  or GNAME11000(G11000,G36177,G10769);
  nand GNAME11001(G11001,G10798,G10843);
  or GNAME11002(G11002,G10843,G10798);
  or GNAME11003(G11003,G36421,G10766);
  or GNAME11004(G11004,G36176,G10767);
  nand GNAME11005(G11005,G10799,G10845);
  or GNAME11006(G11006,G10845,G10799);
  or GNAME11007(G11007,G36420,G10764);
  or GNAME11008(G11008,G36175,G10765);
  nand GNAME11009(G11009,G10800,G10847);
  or GNAME11010(G11010,G10847,G10800);
  or GNAME11011(G11011,G36419,G10762);
  or GNAME11012(G11012,G36174,G10763);
  nand GNAME11013(G11013,G10801,G10849);
  or GNAME11014(G11014,G10849,G10801);
  or GNAME11015(G11015,G36418,G10760);
  or GNAME11016(G11016,G36173,G10761);
  nand GNAME11017(G11017,G10802,G10851);
  or GNAME11018(G11018,G10851,G10802);
  or GNAME11019(G11019,G36399,G10853);
  or GNAME11020(G11020,G36154,G10723);
  nand GNAME11021(G11021,G10722,G10803);
  or GNAME11022(G11022,G10722,G10803);
  or GNAME11023(G11023,G36417,G10758);
  or GNAME11024(G11024,G36172,G10759);
  nand GNAME11025(G11025,G10804,G10854);
  or GNAME11026(G11026,G10854,G10804);
  or GNAME11027(G11027,G36416,G10756);
  or GNAME11028(G11028,G36171,G10757);
  nand GNAME11029(G11029,G10805,G10856);
  or GNAME11030(G11030,G10856,G10805);
  or GNAME11031(G11031,G36415,G10754);
  or GNAME11032(G11032,G36170,G10755);
  nand GNAME11033(G11033,G10806,G10858);
  or GNAME11034(G11034,G10858,G10806);
  or GNAME11035(G11035,G36414,G10752);
  or GNAME11036(G11036,G36169,G10753);
  nand GNAME11037(G11037,G10807,G10860);
  or GNAME11038(G11038,G10860,G10807);
  or GNAME11039(G11039,G36413,G10750);
  or GNAME11040(G11040,G36168,G10751);
  nand GNAME11041(G11041,G10808,G10862);
  or GNAME11042(G11042,G10862,G10808);
  or GNAME11043(G11043,G36412,G10748);
  or GNAME11044(G11044,G36167,G10749);
  nand GNAME11045(G11045,G10809,G10864);
  or GNAME11046(G11046,G10864,G10809);
  or GNAME11047(G11047,G36411,G10746);
  or GNAME11048(G11048,G36166,G10747);
  nand GNAME11049(G11049,G10810,G10866);
  or GNAME11050(G11050,G10866,G10810);
  or GNAME11051(G11051,G36410,G10744);
  or GNAME11052(G11052,G36165,G10745);
  nand GNAME11053(G11053,G10811,G10868);
  or GNAME11054(G11054,G10868,G10811);
  or GNAME11055(G11055,G36409,G10742);
  or GNAME11056(G11056,G36164,G10743);
  nand GNAME11057(G11057,G10812,G10870);
  or GNAME11058(G11058,G10870,G10812);
  or GNAME11059(G11059,G36408,G10740);
  or GNAME11060(G11060,G36163,G10741);
  nand GNAME11061(G11061,G10813,G10872);
  or GNAME11062(G11062,G10872,G10813);
  and GNAME11063(G11063,G11341,G11342);
  and GNAME11064(G11064,G11337,G11339);
  and GNAME11065(G11065,G11333,G11334);
  and GNAME11066(G11066,G11330,G11331);
  and GNAME11067(G11067,G11326,G11328);
  and GNAME11068(G11068,G11323,G11325);
  and GNAME11069(G11069,G11235,G11237);
  and GNAME11070(G11070,G11229,G11230);
  and GNAME11071(G11071,G11225,G11227);
  not GNAME11072(G11072,G1209);
  not GNAME11073(G11073,G1274);
  not GNAME11074(G11074,G1273);
  not GNAME11075(G11075,G1272);
  not GNAME11076(G11076,G1271);
  not GNAME11077(G11077,G1270);
  not GNAME11078(G11078,G1269);
  not GNAME11079(G11079,G1268);
  not GNAME11080(G11080,G1267);
  not GNAME11081(G11081,G1266);
  not GNAME11082(G11082,G1265);
  and GNAME11083(G11083,G11223,G11198);
  or GNAME11084(G11084,G11195,G11083);
  not GNAME11085(G11085,G1243);
  not GNAME11086(G11086,G1264);
  not GNAME11087(G11087,G1263);
  not GNAME11088(G11088,G1262);
  not GNAME11089(G11089,G1261);
  not GNAME11090(G11090,G1260);
  not GNAME11091(G11091,G1259);
  not GNAME11092(G11092,G1258);
  not GNAME11093(G11093,G1257);
  not GNAME11094(G11094,G1256);
  not GNAME11095(G11095,G1255);
  not GNAME11096(G11096,G1254);
  not GNAME11097(G11097,G1253);
  not GNAME11098(G11098,G1252);
  not GNAME11099(G11099,G1251);
  not GNAME11100(G11100,G1250);
  not GNAME11101(G11101,G1249);
  not GNAME11102(G11102,G1248);
  not GNAME11103(G11103,G1247);
  not GNAME11104(G11104,G1246);
  not GNAME11105(G11105,G1245);
  nor GNAME11106(G11106,G11319,G11107);
  and GNAME11107(G11107,G11318,G11317);
  and GNAME11108(G11108,G11233,G11204);
  or GNAME11109(G11109,G11201,G11108);
  and GNAME11110(G11110,G11259,G11258);
  nor GNAME11111(G11111,G11260,G11110);
  and GNAME11112(G11112,G11335,G11220);
  or GNAME11113(G11113,G11244,G11112);
  and GNAME11114(G11114,G11381,G11382);
  and GNAME11115(G11115,G11386,G11387);
  and GNAME11116(G11116,G11391,G11392);
  nand GNAME11117(G11117,G11503,G11504);
  nand GNAME11118(G11118,G11393,G11394);
  nand GNAME11119(G11119,G11395,G11396);
  nand GNAME11120(G11120,G11397,G11398);
  nand GNAME11121(G11121,G11399,G11400);
  nand GNAME11122(G11122,G11467,G11468);
  nand GNAME11123(G11123,G11469,G11470);
  nand GNAME11124(G11124,G11471,G11472);
  nand GNAME11125(G11125,G11473,G11474);
  nand GNAME11126(G11126,G11475,G11476);
  nand GNAME11127(G11127,G11477,G11478);
  nand GNAME11128(G11128,G11479,G11480);
  nand GNAME11129(G11129,G11481,G11482);
  nand GNAME11130(G11130,G11483,G11484);
  nand GNAME11131(G11131,G11485,G11486);
  nand GNAME11132(G11132,G11487,G11488);
  nand GNAME11133(G11133,G11489,G11490);
  nand GNAME11134(G11134,G11491,G11492);
  nand GNAME11135(G11135,G11493,G11494);
  nand GNAME11136(G11136,G11495,G11496);
  nand GNAME11137(G11137,G11497,G11498);
  nand GNAME11138(G11138,G11499,G11500);
  nand GNAME11139(G11139,G11501,G11502);
  not GNAME11140(G11140,G1231);
  not GNAME11141(G11141,G1233);
  not GNAME11142(G11142,G1234);
  not GNAME11143(G11143,G1235);
  not GNAME11144(G11144,G1237);
  not GNAME11145(G11145,G1238);
  not GNAME11146(G11146,G1239);
  nand GNAME11147(G11147,G11215,G11194);
  nand GNAME11148(G11148,G11221,G11192);
  nand GNAME11149(G11149,G11209,G11200);
  not GNAME11150(G11150,G1211);
  not GNAME11151(G11151,G1210);
  not GNAME11152(G11152,G1225);
  not GNAME11153(G11153,G1226);
  not GNAME11154(G11154,G1229);
  not GNAME11155(G11155,G1230);
  not GNAME11156(G11156,G1228);
  not GNAME11157(G11157,G1227);
  not GNAME11158(G11158,G1224);
  not GNAME11159(G11159,G1223);
  not GNAME11160(G11160,G1222);
  not GNAME11161(G11161,G1221);
  not GNAME11162(G11162,G1220);
  not GNAME11163(G11163,G1219);
  not GNAME11164(G11164,G1218);
  not GNAME11165(G11165,G1217);
  not GNAME11166(G11166,G1216);
  not GNAME11167(G11167,G1215);
  not GNAME11168(G11168,G1214);
  not GNAME11169(G11169,G1213);
  not GNAME11170(G11170,G1212);
  nand GNAME11171(G11171,G11314,G11313);
  nand GNAME11172(G11172,G11310,G11309);
  nand GNAME11173(G11173,G11306,G11305);
  nand GNAME11174(G11174,G11302,G11301);
  nand GNAME11175(G11175,G11298,G11297);
  nand GNAME11176(G11176,G11294,G11293);
  nand GNAME11177(G11177,G11290,G11289);
  nand GNAME11178(G11178,G11286,G11285);
  nand GNAME11179(G11179,G11282,G11281);
  nand GNAME11180(G11180,G11278,G11277);
  nand GNAME11181(G11181,G11231,G11191);
  nand GNAME11182(G11182,G11274,G11273);
  nand GNAME11183(G11183,G11270,G11269);
  nand GNAME11184(G11184,G11266,G11265);
  nand GNAME11185(G11185,G11262,G11240);
  or GNAME11186(G11186,G11111,G11241);
  nand GNAME11187(G11187,G11255,G11254);
  nand GNAME11188(G11188,G11251,G11243);
  nand GNAME11189(G11189,G11205,G11191);
  or GNAME11190(G11190,G11116,G11081);
  or GNAME11191(G11191,G11114,G11073);
  or GNAME11192(G11192,G11115,G11077);
  nand GNAME11193(G11193,G11080,G11369,G11370);
  nand GNAME11194(G11194,G11390,G1267);
  and GNAME11195(G11195,G11079,G11371,G11372);
  nand GNAME11196(G11196,G11389,G1268);
  nand GNAME11197(G11197,G11078,G11373,G11374);
  nand GNAME11198(G11198,G11388,G1269);
  nand GNAME11199(G11199,G11076,G11375,G11376);
  nand GNAME11200(G11200,G11385,G1271);
  and GNAME11201(G11201,G11075,G11377,G11378);
  nand GNAME11202(G11202,G11384,G1272);
  nand GNAME11203(G11203,G11074,G11379,G11380);
  nand GNAME11204(G11204,G11383,G1273);
  nand GNAME11205(G11205,G11073,G11114);
  nand GNAME11206(G11206,G11233,G11204);
  nand GNAME11207(G11207,G11506,G11206);
  nand GNAME11208(G11208,G11207,G11202);
  nand GNAME11209(G11209,G11199,G11208);
  not GNAME11210(G11210,G11149);
  nand GNAME11211(G11211,G11077,G11115);
  nand GNAME11212(G11212,G11223,G11198);
  nand GNAME11213(G11213,G11505,G11212);
  nand GNAME11214(G11214,G11213,G11196);
  nand GNAME11215(G11215,G11193,G11214);
  not GNAME11216(G11216,G11147);
  nand GNAME11217(G11217,G11081,G11116);
  not GNAME11218(G11218,G11247);
  nand GNAME11219(G11219,G11082,G11366,G11367);
  nand GNAME11220(G11220,G11368,G1265);
  nand GNAME11221(G11221,G11149,G11211);
  not GNAME11222(G11222,G11148);
  nand GNAME11223(G11223,G11197,G11148);
  nand GNAME11224(G11224,G11196,G11084);
  nand GNAME11225(G11225,G11224,G11193,G11194);
  nand GNAME11226(G11226,G11193,G11194);
  nand GNAME11227(G11227,G11226,G11196,G11084);
  or GNAME11228(G11228,G11195,G11508);
  nand GNAME11229(G11229,G11228,G11083);
  or GNAME11230(G11230,G11508,G11084);
  nand GNAME11231(G11231,G11205,G1209);
  not GNAME11232(G11232,G11181);
  nand GNAME11233(G11233,G11203,G11181);
  nand GNAME11234(G11234,G11202,G11109);
  nand GNAME11235(G11235,G11234,G11199,G11200);
  nand GNAME11236(G11236,G11199,G11200);
  nand GNAME11237(G11237,G11236,G11202,G11109);
  and GNAME11238(G11238,G11404,G1243);
  nand GNAME11239(G11239,G11091,G11407,G11408);
  nand GNAME11240(G11240,G11424,G1259);
  and GNAME11241(G11241,G11423,G1260);
  nand GNAME11242(G11242,G11087,G11411,G11412);
  nand GNAME11243(G11243,G11416,G1263);
  and GNAME11244(G11244,G11086,G11413,G11414);
  nand GNAME11245(G11245,G11415,G1264);
  nand GNAME11246(G11246,G11147,G11217);
  nand GNAME11247(G11247,G11246,G11190);
  nand GNAME11248(G11248,G11335,G11220);
  nand GNAME11249(G11249,G11507,G11248);
  nand GNAME11250(G11250,G11249,G11245);
  nand GNAME11251(G11251,G11242,G11250);
  not GNAME11252(G11252,G11188);
  nand GNAME11253(G11253,G11088,G11417,G11418);
  nand GNAME11254(G11254,G11419,G1262);
  nand GNAME11255(G11255,G11188,G11253);
  not GNAME11256(G11256,G11187);
  nand GNAME11257(G11257,G11089,G11420,G11421);
  nand GNAME11258(G11258,G11422,G1261);
  nand GNAME11259(G11259,G11187,G11257);
  and GNAME11260(G11260,G11090,G11409,G11410);
  not GNAME11261(G11261,G11186);
  nand GNAME11262(G11262,G11239,G11186);
  not GNAME11263(G11263,G11185);
  nand GNAME11264(G11264,G11092,G11425,G11426);
  nand GNAME11265(G11265,G11427,G1258);
  nand GNAME11266(G11266,G11185,G11264);
  not GNAME11267(G11267,G11184);
  nand GNAME11268(G11268,G11093,G11428,G11429);
  nand GNAME11269(G11269,G11430,G1257);
  nand GNAME11270(G11270,G11184,G11268);
  not GNAME11271(G11271,G11183);
  nand GNAME11272(G11272,G11094,G11431,G11432);
  nand GNAME11273(G11273,G11433,G1256);
  nand GNAME11274(G11274,G11183,G11272);
  not GNAME11275(G11275,G11182);
  nand GNAME11276(G11276,G11095,G11434,G11435);
  nand GNAME11277(G11277,G11436,G1255);
  nand GNAME11278(G11278,G11182,G11276);
  not GNAME11279(G11279,G11180);
  nand GNAME11280(G11280,G11096,G11437,G11438);
  nand GNAME11281(G11281,G11439,G1254);
  nand GNAME11282(G11282,G11180,G11280);
  not GNAME11283(G11283,G11179);
  nand GNAME11284(G11284,G11097,G11440,G11441);
  nand GNAME11285(G11285,G11442,G1253);
  nand GNAME11286(G11286,G11179,G11284);
  not GNAME11287(G11287,G11178);
  nand GNAME11288(G11288,G11098,G11443,G11444);
  nand GNAME11289(G11289,G11445,G1252);
  nand GNAME11290(G11290,G11178,G11288);
  not GNAME11291(G11291,G11177);
  nand GNAME11292(G11292,G11099,G11446,G11447);
  nand GNAME11293(G11293,G11448,G1251);
  nand GNAME11294(G11294,G11177,G11292);
  not GNAME11295(G11295,G11176);
  nand GNAME11296(G11296,G11100,G11449,G11450);
  nand GNAME11297(G11297,G11451,G1250);
  nand GNAME11298(G11298,G11176,G11296);
  not GNAME11299(G11299,G11175);
  nand GNAME11300(G11300,G11101,G11452,G11453);
  nand GNAME11301(G11301,G11454,G1249);
  nand GNAME11302(G11302,G11175,G11300);
  not GNAME11303(G11303,G11174);
  nand GNAME11304(G11304,G11102,G11455,G11456);
  nand GNAME11305(G11305,G11457,G1248);
  nand GNAME11306(G11306,G11174,G11304);
  not GNAME11307(G11307,G11173);
  nand GNAME11308(G11308,G11103,G11458,G11459);
  nand GNAME11309(G11309,G11460,G1247);
  nand GNAME11310(G11310,G11173,G11308);
  not GNAME11311(G11311,G11172);
  nand GNAME11312(G11312,G11104,G11461,G11462);
  nand GNAME11313(G11313,G11463,G1246);
  nand GNAME11314(G11314,G11172,G11312);
  not GNAME11315(G11315,G11171);
  nand GNAME11316(G11316,G11105,G11464,G11465);
  nand GNAME11317(G11317,G11466,G1245);
  nand GNAME11318(G11318,G11171,G11316);
  and GNAME11319(G11319,G11085,G11405,G11406);
  or GNAME11320(G11320,G11238,G11106);
  nand GNAME11321(G11321,G11320,G1241);
  or GNAME11322(G11322,G11106,G1241,G11238);
  nand GNAME11323(G11323,G11403,G11321,G11322);
  nand GNAME11324(G11324,G11321,G11322);
  nand GNAME11325(G11325,G11324,G11401,G11402);
  or GNAME11326(G11326,G11238,G11509);
  or GNAME11327(G11327,G11238,G11319);
  nand GNAME11328(G11328,G11327,G11107);
  or GNAME11329(G11329,G11201,G11510);
  nand GNAME11330(G11330,G11329,G11108);
  or GNAME11331(G11331,G11510,G11109);
  or GNAME11332(G11332,G11241,G11260);
  nand GNAME11333(G11333,G11332,G11110);
  or GNAME11334(G11334,G11241,G11511);
  nand GNAME11335(G11335,G11247,G11219);
  nand GNAME11336(G11336,G11245,G11113);
  nand GNAME11337(G11337,G11336,G11242,G11243);
  nand GNAME11338(G11338,G11242,G11243);
  nand GNAME11339(G11339,G11338,G11245,G11113);
  or GNAME11340(G11340,G11244,G11512);
  nand GNAME11341(G11341,G11340,G11112);
  or GNAME11342(G11342,G11512,G11113);
  not GNAME11343(G11343,G11189);
  nand GNAME11344(G11344,G11219,G11220);
  nand GNAME11345(G11345,G11190,G11217);
  nand GNAME11346(G11346,G11197,G11198);
  nand GNAME11347(G11347,G11192,G11211);
  nand GNAME11348(G11348,G11316,G11317);
  nand GNAME11349(G11349,G11312,G11313);
  nand GNAME11350(G11350,G11308,G11309);
  nand GNAME11351(G11351,G11304,G11305);
  nand GNAME11352(G11352,G11300,G11301);
  nand GNAME11353(G11353,G11296,G11297);
  nand GNAME11354(G11354,G11292,G11293);
  nand GNAME11355(G11355,G11288,G11289);
  nand GNAME11356(G11356,G11284,G11285);
  nand GNAME11357(G11357,G11280,G11281);
  nand GNAME11358(G11358,G11203,G11204);
  nand GNAME11359(G11359,G11276,G11277);
  nand GNAME11360(G11360,G11272,G11273);
  nand GNAME11361(G11361,G11268,G11269);
  nand GNAME11362(G11362,G11264,G11265);
  nand GNAME11363(G11363,G11239,G11240);
  nand GNAME11364(G11364,G11257,G11258);
  nand GNAME11365(G11365,G11253,G11254);
  nand GNAME11366(G11366,G11140,G1209);
  nand GNAME11367(G11367,G11072,G1231);
  nand GNAME11368(G11368,G11366,G11367);
  nand GNAME11369(G11369,G11141,G1209);
  nand GNAME11370(G11370,G11072,G1233);
  nand GNAME11371(G11371,G11142,G1209);
  nand GNAME11372(G11372,G11072,G1234);
  nand GNAME11373(G11373,G11143,G1209);
  nand GNAME11374(G11374,G11072,G1235);
  nand GNAME11375(G11375,G11144,G1209);
  nand GNAME11376(G11376,G11072,G1237);
  nand GNAME11377(G11377,G11145,G1209);
  nand GNAME11378(G11378,G11072,G1238);
  nand GNAME11379(G11379,G11146,G1209);
  nand GNAME11380(G11380,G11072,G1239);
  or GNAME11381(G11381,G1240,G11072);
  nand GNAME11382(G11382,G11072,G1240);
  nand GNAME11383(G11383,G11379,G11380);
  nand GNAME11384(G11384,G11377,G11378);
  nand GNAME11385(G11385,G11375,G11376);
  or GNAME11386(G11386,G1236,G11072);
  nand GNAME11387(G11387,G11072,G1236);
  nand GNAME11388(G11388,G11373,G11374);
  nand GNAME11389(G11389,G11371,G11372);
  nand GNAME11390(G11390,G11369,G11370);
  or GNAME11391(G11391,G1232,G11072);
  nand GNAME11392(G11392,G11072,G1232);
  nand GNAME11393(G11393,G11247,G11344);
  nand GNAME11394(G11394,G11218,G11219,G11220);
  nand GNAME11395(G11395,G11147,G11345);
  nand GNAME11396(G11396,G11216,G11190,G11217);
  nand GNAME11397(G11397,G11148,G11346);
  nand GNAME11398(G11398,G11222,G11197,G11198);
  nand GNAME11399(G11399,G11149,G11347);
  nand GNAME11400(G11400,G11210,G11192,G11211);
  nand GNAME11401(G11401,G11150,G1209);
  nand GNAME11402(G11402,G11072,G1211);
  nand GNAME11403(G11403,G11401,G11402);
  nand GNAME11404(G11404,G11405,G11406);
  nand GNAME11405(G11405,G11151,G1209);
  nand GNAME11406(G11406,G11072,G1210);
  nand GNAME11407(G11407,G11152,G1209);
  nand GNAME11408(G11408,G11072,G1225);
  nand GNAME11409(G11409,G11153,G1209);
  nand GNAME11410(G11410,G11072,G1226);
  nand GNAME11411(G11411,G11154,G1209);
  nand GNAME11412(G11412,G11072,G1229);
  nand GNAME11413(G11413,G11155,G1209);
  nand GNAME11414(G11414,G11072,G1230);
  nand GNAME11415(G11415,G11413,G11414);
  nand GNAME11416(G11416,G11411,G11412);
  nand GNAME11417(G11417,G11156,G1209);
  nand GNAME11418(G11418,G11072,G1228);
  nand GNAME11419(G11419,G11417,G11418);
  nand GNAME11420(G11420,G11157,G1209);
  nand GNAME11421(G11421,G11072,G1227);
  nand GNAME11422(G11422,G11420,G11421);
  nand GNAME11423(G11423,G11409,G11410);
  nand GNAME11424(G11424,G11407,G11408);
  nand GNAME11425(G11425,G11158,G1209);
  nand GNAME11426(G11426,G11072,G1224);
  nand GNAME11427(G11427,G11425,G11426);
  nand GNAME11428(G11428,G11159,G1209);
  nand GNAME11429(G11429,G11072,G1223);
  nand GNAME11430(G11430,G11428,G11429);
  nand GNAME11431(G11431,G11160,G1209);
  nand GNAME11432(G11432,G11072,G1222);
  nand GNAME11433(G11433,G11431,G11432);
  nand GNAME11434(G11434,G11161,G1209);
  nand GNAME11435(G11435,G11072,G1221);
  nand GNAME11436(G11436,G11434,G11435);
  nand GNAME11437(G11437,G11162,G1209);
  nand GNAME11438(G11438,G11072,G1220);
  nand GNAME11439(G11439,G11437,G11438);
  nand GNAME11440(G11440,G11163,G1209);
  nand GNAME11441(G11441,G11072,G1219);
  nand GNAME11442(G11442,G11440,G11441);
  nand GNAME11443(G11443,G11164,G1209);
  nand GNAME11444(G11444,G11072,G1218);
  nand GNAME11445(G11445,G11443,G11444);
  nand GNAME11446(G11446,G11165,G1209);
  nand GNAME11447(G11447,G11072,G1217);
  nand GNAME11448(G11448,G11446,G11447);
  nand GNAME11449(G11449,G11166,G1209);
  nand GNAME11450(G11450,G11072,G1216);
  nand GNAME11451(G11451,G11449,G11450);
  nand GNAME11452(G11452,G11167,G1209);
  nand GNAME11453(G11453,G11072,G1215);
  nand GNAME11454(G11454,G11452,G11453);
  nand GNAME11455(G11455,G11168,G1209);
  nand GNAME11456(G11456,G11072,G1214);
  nand GNAME11457(G11457,G11455,G11456);
  nand GNAME11458(G11458,G11169,G1209);
  nand GNAME11459(G11459,G11072,G1213);
  nand GNAME11460(G11460,G11458,G11459);
  nand GNAME11461(G11461,G11170,G1209);
  nand GNAME11462(G11462,G11072,G1212);
  nand GNAME11463(G11463,G11461,G11462);
  nand GNAME11464(G11464,G11150,G1209);
  nand GNAME11465(G11465,G11072,G1211);
  nand GNAME11466(G11466,G11464,G11465);
  nand GNAME11467(G11467,G11171,G11348);
  nand GNAME11468(G11468,G11315,G11316,G11317);
  nand GNAME11469(G11469,G11172,G11349);
  nand GNAME11470(G11470,G11311,G11312,G11313);
  nand GNAME11471(G11471,G11173,G11350);
  nand GNAME11472(G11472,G11307,G11308,G11309);
  nand GNAME11473(G11473,G11174,G11351);
  nand GNAME11474(G11474,G11303,G11304,G11305);
  nand GNAME11475(G11475,G11175,G11352);
  nand GNAME11476(G11476,G11299,G11300,G11301);
  nand GNAME11477(G11477,G11176,G11353);
  nand GNAME11478(G11478,G11295,G11296,G11297);
  nand GNAME11479(G11479,G11177,G11354);
  nand GNAME11480(G11480,G11291,G11292,G11293);
  nand GNAME11481(G11481,G11178,G11355);
  nand GNAME11482(G11482,G11287,G11288,G11289);
  nand GNAME11483(G11483,G11179,G11356);
  nand GNAME11484(G11484,G11283,G11284,G11285);
  nand GNAME11485(G11485,G11180,G11357);
  nand GNAME11486(G11486,G11279,G11280,G11281);
  nand GNAME11487(G11487,G11181,G11358);
  nand GNAME11488(G11488,G11232,G11203,G11204);
  nand GNAME11489(G11489,G11182,G11359);
  nand GNAME11490(G11490,G11275,G11276,G11277);
  nand GNAME11491(G11491,G11183,G11360);
  nand GNAME11492(G11492,G11271,G11272,G11273);
  nand GNAME11493(G11493,G11184,G11361);
  nand GNAME11494(G11494,G11267,G11268,G11269);
  nand GNAME11495(G11495,G11185,G11362);
  nand GNAME11496(G11496,G11263,G11264,G11265);
  nand GNAME11497(G11497,G11186,G11363);
  nand GNAME11498(G11498,G11261,G11239,G11240);
  nand GNAME11499(G11499,G11187,G11364);
  nand GNAME11500(G11500,G11256,G11257,G11258);
  nand GNAME11501(G11501,G11188,G11365);
  nand GNAME11502(G11502,G11252,G11253,G11254);
  nand GNAME11503(G11503,G11189,G1209);
  nand GNAME11504(G11504,G11072,G11343);
  not GNAME11505(G11505,G11195);
  not GNAME11506(G11506,G11201);
  not GNAME11507(G11507,G11244);
  not GNAME11508(G11508,G11196);
  not GNAME11509(G11509,G11106);
  not GNAME11510(G11510,G11202);
  not GNAME11511(G11511,G11111);
  not GNAME11512(G11512,G11245);
  and GNAME11513(G11513,G11650,G11651);
  and GNAME11514(G11514,G11646,G11648);
  and GNAME11515(G11515,G11643,G11645);
  and GNAME11516(G11516,G11641,G11642);
  and GNAME11517(G11517,G11636,G11638);
  nand GNAME11518(G11518,G11655,G11690,G11691);
  not GNAME11519(G11519,G1722);
  nand GNAME11520(G11520,G1913,G1722);
  not GNAME11521(G11521,G1912);
  not GNAME11522(G11522,G1731);
  not GNAME11523(G11523,G1901);
  not GNAME11524(G11524,G1734);
  not GNAME11525(G11525,G1900);
  not GNAME11526(G11526,G1746);
  not GNAME11527(G11527,G1896);
  not GNAME11528(G11528,G1749);
  not GNAME11529(G11529,G1895);
  not GNAME11530(G11530,G1894);
  not GNAME11531(G11531,G1752);
  not GNAME11532(G11532,G1910);
  not GNAME11533(G11533,G1761);
  not GNAME11534(G11534,G1909);
  not GNAME11535(G11535,G1764);
  not GNAME11536(G11536,G1908);
  not GNAME11537(G11537,G1905);
  not GNAME11538(G11538,G1773);
  nor GNAME11539(G11539,G11724,G11545);
  not GNAME11540(G11540,G1904);
  not GNAME11541(G11541,G1776);
  and GNAME11542(G11542,G11630,G11631);
  not GNAME11543(G11543,G1903);
  not GNAME11544(G11544,G1779);
  and GNAME11545(G11545,G11624,G11639);
  or GNAME11546(G11546,G11623,G11547);
  and GNAME11547(G11547,G11621,G11622);
  and GNAME11548(G11548,G11614,G11615);
  and GNAME11549(G11549,G11611,G11612);
  or GNAME11550(G11550,G11613,G11549);
  nand GNAME11551(G11551,G11722,G11723);
  nand GNAME11552(G11552,G11659,G11660);
  nand GNAME11553(G11553,G11664,G11665);
  nand GNAME11554(G11554,G11669,G11670);
  nand GNAME11555(G11555,G11671,G11672);
  nand GNAME11556(G11556,G11673,G11674);
  nand GNAME11557(G11557,G11675,G11676);
  nand GNAME11558(G11558,G11680,G11681);
  nand GNAME11559(G11559,G11685,G11686);
  nand GNAME11560(G11560,G11698,G11699);
  nand GNAME11561(G11561,G11703,G11704);
  nand GNAME11562(G11562,G11708,G11709);
  nand GNAME11563(G11563,G11713,G11714);
  nand GNAME11564(G11564,G11718,G11719);
  nand GNAME11565(G11565,G11603,G11604);
  nand GNAME11566(G11566,G11600,G11601);
  nand GNAME11567(G11567,G11605,G11598);
  and GNAME11568(G11568,G11595,G11593);
  and GNAME11569(G11569,G11606,G11591);
  and GNAME11570(G11570,G11587,G11588);
  nand GNAME11571(G11571,G11584,G11585);
  or GNAME11572(G11572,G11582,G11573);
  nor GNAME11573(G11573,G11520,G11521);
  not GNAME11574(G11574,G1902);
  not GNAME11575(G11575,G1721);
  and GNAME11576(G11576,G11626,G11627);
  nand GNAME11577(G11577,G11618,G11619);
  or GNAME11578(G11578,G11616,G11548);
  not GNAME11579(G11579,G11539);
  not GNAME11580(G11580,G11520);
  or GNAME11581(G11581,G11580,G1912);
  and GNAME11582(G11582,G11581,G1728);
  nand GNAME11583(G11583,G11523,G11522);
  nand GNAME11584(G11584,G11572,G11583);
  or GNAME11585(G11585,G11522,G11523);
  nand GNAME11586(G11586,G11525,G11524);
  nand GNAME11587(G11587,G11571,G11586);
  or GNAME11588(G11588,G11524,G11525);
  not GNAME11589(G11589,G11570);
  or GNAME11590(G11590,G1737,G1899);
  nand GNAME11591(G11591,G11589,G11590);
  not GNAME11592(G11592,G11569);
  nand GNAME11593(G11593,G1740,G1898);
  or GNAME11594(G11594,G1898,G1740);
  nand GNAME11595(G11595,G11592,G11594);
  not GNAME11596(G11596,G11568);
  or GNAME11597(G11597,G1897,G1743);
  nand GNAME11598(G11598,G11596,G11597);
  nand GNAME11599(G11599,G11527,G11526);
  nand GNAME11600(G11600,G11567,G11599);
  or GNAME11601(G11601,G11526,G11527);
  nand GNAME11602(G11602,G11529,G11528);
  nand GNAME11603(G11603,G11566,G11602);
  or GNAME11604(G11604,G11528,G11529);
  nand GNAME11605(G11605,G1743,G1897);
  nand GNAME11606(G11606,G1899,G1737);
  nand GNAME11607(G11607,G1770,G1906);
  and GNAME11608(G11608,G1767,G1907);
  and GNAME11609(G11609,G1755,G1911);
  nand GNAME11610(G11610,G11530,G11531);
  nand GNAME11611(G11611,G11565,G11610);
  or GNAME11612(G11612,G11530,G11531);
  nor GNAME11613(G11613,G1911,G1755);
  nand GNAME11614(G11614,G11726,G11550);
  or GNAME11615(G11615,G1758,G1910);
  and GNAME11616(G11616,G1758,G1910);
  nand GNAME11617(G11617,G11534,G11533);
  nand GNAME11618(G11618,G11578,G11617);
  or GNAME11619(G11619,G11533,G11534);
  nand GNAME11620(G11620,G11536,G11535);
  nand GNAME11621(G11621,G11577,G11620);
  or GNAME11622(G11622,G11535,G11536);
  nor GNAME11623(G11623,G1907,G1767);
  nand GNAME11624(G11624,G11725,G11546);
  or GNAME11625(G11625,G11537,G11538);
  nand GNAME11626(G11626,G11625,G11539);
  nand GNAME11627(G11627,G11537,G11538);
  not GNAME11628(G11628,G11576);
  or GNAME11629(G11629,G11540,G11541);
  nand GNAME11630(G11630,G11628,G11629);
  nand GNAME11631(G11631,G11540,G11541);
  not GNAME11632(G11632,G11542);
  nand GNAME11633(G11633,G11544,G11543);
  nand GNAME11634(G11634,G11633,G11542);
  or GNAME11635(G11635,G11543,G11544);
  nand GNAME11636(G11636,G11692,G11693,G11634,G11635);
  nand GNAME11637(G11637,G11632,G11635);
  nand GNAME11638(G11638,G11694,G11637,G11633);
  or GNAME11639(G11639,G1906,G1770);
  nand GNAME11640(G11640,G11607,G11639);
  nand GNAME11641(G11641,G11640,G11725,G11546);
  nand GNAME11642(G11642,G11607,G11545);
  or GNAME11643(G11643,G11608,G11546);
  or GNAME11644(G11644,G11608,G11623);
  nand GNAME11645(G11645,G11644,G11547);
  nand GNAME11646(G11646,G11720,G11721,G11726,G11550);
  nand GNAME11647(G11647,G1758,G1910);
  nand GNAME11648(G11648,G11647,G11548);
  or GNAME11649(G11649,G11609,G11613);
  nand GNAME11650(G11650,G11649,G11549);
  or GNAME11651(G11651,G11609,G11550);
  nand GNAME11652(G11652,G11597,G11605);
  nand GNAME11653(G11653,G11593,G11594);
  nand GNAME11654(G11654,G11590,G11606);
  nand GNAME11655(G11655,G11521,G11689);
  or GNAME11656(G11656,G1752,G11530);
  or GNAME11657(G11657,G1894,G11531);
  and GNAME11658(G11658,G11656,G11657);
  nand GNAME11659(G11659,G11565,G11656,G11657);
  or GNAME11660(G11660,G11658,G11565);
  or GNAME11661(G11661,G1749,G11529);
  or GNAME11662(G11662,G1895,G11528);
  and GNAME11663(G11663,G11661,G11662);
  nand GNAME11664(G11664,G11566,G11661,G11662);
  or GNAME11665(G11665,G11663,G11566);
  or GNAME11666(G11666,G1746,G11527);
  or GNAME11667(G11667,G1896,G11526);
  and GNAME11668(G11668,G11666,G11667);
  nand GNAME11669(G11669,G11567,G11666,G11667);
  or GNAME11670(G11670,G11668,G11567);
  nand GNAME11671(G11671,G11596,G11652);
  nand GNAME11672(G11672,G11568,G11597,G11605);
  nand GNAME11673(G11673,G11592,G11653);
  nand GNAME11674(G11674,G11569,G11593,G11594);
  nand GNAME11675(G11675,G11589,G11654);
  nand GNAME11676(G11676,G11570,G11590,G11606);
  or GNAME11677(G11677,G1734,G11525);
  or GNAME11678(G11678,G1900,G11524);
  and GNAME11679(G11679,G11677,G11678);
  nand GNAME11680(G11680,G11571,G11677,G11678);
  or GNAME11681(G11681,G11679,G11571);
  or GNAME11682(G11682,G1731,G11523);
  or GNAME11683(G11683,G1901,G11522);
  and GNAME11684(G11684,G11682,G11683);
  nand GNAME11685(G11685,G11572,G11682,G11683);
  or GNAME11686(G11686,G11684,G11572);
  nand GNAME11687(G11687,G11520,G1728);
  or GNAME11688(G11688,G1728,G11520);
  nand GNAME11689(G11689,G11687,G11688);
  or GNAME11690(G11690,G1728,G11580,G11521);
  nand GNAME11691(G11691,G1728,G11573);
  or GNAME11692(G11692,G1721,G11574);
  or GNAME11693(G11693,G1902,G11575);
  nand GNAME11694(G11694,G11692,G11693);
  or GNAME11695(G11695,G1903,G11544);
  or GNAME11696(G11696,G1779,G11543);
  nand GNAME11697(G11697,G11695,G11696);
  nand GNAME11698(G11698,G11632,G11697);
  nand GNAME11699(G11699,G11542,G11695,G11696);
  or GNAME11700(G11700,G1904,G11541);
  or GNAME11701(G11701,G1776,G11540);
  nand GNAME11702(G11702,G11700,G11701);
  nand GNAME11703(G11703,G11628,G11702);
  nand GNAME11704(G11704,G11576,G11700,G11701);
  or GNAME11705(G11705,G1905,G11538);
  or GNAME11706(G11706,G1773,G11537);
  nand GNAME11707(G11707,G11705,G11706);
  nand GNAME11708(G11708,G11579,G11705,G11706);
  nand GNAME11709(G11709,G11539,G11707);
  or GNAME11710(G11710,G1764,G11536);
  or GNAME11711(G11711,G1908,G11535);
  and GNAME11712(G11712,G11710,G11711);
  nand GNAME11713(G11713,G11577,G11710,G11711);
  or GNAME11714(G11714,G11712,G11577);
  or GNAME11715(G11715,G1761,G11534);
  or GNAME11716(G11716,G1909,G11533);
  and GNAME11717(G11717,G11715,G11716);
  nand GNAME11718(G11718,G11578,G11715,G11716);
  or GNAME11719(G11719,G11717,G11578);
  or GNAME11720(G11720,G1758,G11532);
  nand GNAME11721(G11721,G11532,G1758);
  or GNAME11722(G11722,G1913,G11519);
  nand GNAME11723(G11723,G11519,G1913);
  not GNAME11724(G11724,G11607);
  not GNAME11725(G11725,G11608);
  not GNAME11726(G11726,G11609);
  nand GNAME11727(G11727,G11852,G11851);
  not GNAME11728(G11728,G1729);
  not GNAME11729(G11729,G1870);
  not GNAME11730(G11730,G1735);
  not GNAME11731(G11731,G1866);
  not GNAME11732(G11732,G1741);
  not GNAME11733(G11733,G1864);
  not GNAME11734(G11734,G1747);
  not GNAME11735(G11735,G1862);
  not GNAME11736(G11736,G1753);
  not GNAME11737(G11737,G1891);
  not GNAME11738(G11738,G1759);
  not GNAME11739(G11739,G1889);
  not GNAME11740(G11740,G1765);
  not GNAME11741(G11741,G1887);
  not GNAME11742(G11742,G1771);
  not GNAME11743(G11743,G1885);
  not GNAME11744(G11744,G1777);
  not GNAME11745(G11745,G1883);
  not GNAME11746(G11746,G1782);
  not GNAME11747(G11747,G1880);
  not GNAME11748(G11748,G1580);
  not GNAME11749(G11749,G1878);
  not GNAME11750(G11750,G1582);
  not GNAME11751(G11751,G1876);
  not GNAME11752(G11752,G1584);
  not GNAME11753(G11753,G1874);
  not GNAME11754(G11754,G1586);
  not GNAME11755(G11755,G1872);
  not GNAME11756(G11756,G1588);
  not GNAME11757(G11757,G1869);
  not GNAME11758(G11758,G1591);
  not GNAME11759(G11759,G1892);
  nand GNAME11760(G11760,G11728,G1881);
  nand GNAME11761(G11761,G1724,G11759,G11760);
  or GNAME11762(G11762,G1881,G11728);
  nand GNAME11763(G11763,G11729,G1732);
  nand GNAME11764(G11764,G11763,G11761,G11762);
  or GNAME11765(G11765,G1732,G11729);
  nand GNAME11766(G11766,G11730,G1867);
  nand GNAME11767(G11767,G11766,G11764,G11765);
  or GNAME11768(G11768,G1867,G11730);
  nand GNAME11769(G11769,G11731,G1738);
  nand GNAME11770(G11770,G11769,G11767,G11768);
  or GNAME11771(G11771,G1738,G11731);
  nand GNAME11772(G11772,G11732,G1865);
  nand GNAME11773(G11773,G11772,G11770,G11771);
  or GNAME11774(G11774,G1865,G11732);
  nand GNAME11775(G11775,G11733,G1744);
  nand GNAME11776(G11776,G11775,G11773,G11774);
  or GNAME11777(G11777,G1744,G11733);
  nand GNAME11778(G11778,G11734,G1863);
  nand GNAME11779(G11779,G11778,G11776,G11777);
  or GNAME11780(G11780,G1863,G11734);
  nand GNAME11781(G11781,G11735,G1750);
  nand GNAME11782(G11782,G11781,G11779,G11780);
  or GNAME11783(G11783,G1750,G11735);
  nand GNAME11784(G11784,G11736,G1861);
  nand GNAME11785(G11785,G11784,G11782,G11783);
  or GNAME11786(G11786,G1861,G11736);
  nand GNAME11787(G11787,G11737,G1756);
  nand GNAME11788(G11788,G11787,G11785,G11786);
  or GNAME11789(G11789,G1756,G11737);
  nand GNAME11790(G11790,G11738,G1890);
  nand GNAME11791(G11791,G11790,G11788,G11789);
  or GNAME11792(G11792,G1890,G11738);
  nand GNAME11793(G11793,G11739,G1762);
  nand GNAME11794(G11794,G11793,G11791,G11792);
  or GNAME11795(G11795,G1762,G11739);
  nand GNAME11796(G11796,G11740,G1888);
  nand GNAME11797(G11797,G11796,G11794,G11795);
  or GNAME11798(G11798,G1888,G11740);
  nand GNAME11799(G11799,G11741,G1768);
  nand GNAME11800(G11800,G11799,G11797,G11798);
  or GNAME11801(G11801,G1768,G11741);
  nand GNAME11802(G11802,G11742,G1886);
  nand GNAME11803(G11803,G11802,G11800,G11801);
  or GNAME11804(G11804,G1886,G11742);
  nand GNAME11805(G11805,G11743,G1774);
  nand GNAME11806(G11806,G11805,G11803,G11804);
  or GNAME11807(G11807,G1774,G11743);
  nand GNAME11808(G11808,G11744,G1884);
  nand GNAME11809(G11809,G11808,G11806,G11807);
  or GNAME11810(G11810,G1884,G11744);
  nand GNAME11811(G11811,G11745,G1780);
  nand GNAME11812(G11812,G11811,G11809,G11810);
  or GNAME11813(G11813,G1780,G11745);
  nand GNAME11814(G11814,G11746,G1882);
  nand GNAME11815(G11815,G11814,G11812,G11813);
  or GNAME11816(G11816,G1882,G11746);
  nand GNAME11817(G11817,G11747,G1579);
  nand GNAME11818(G11818,G11817,G11815,G11816);
  or GNAME11819(G11819,G1579,G11747);
  nand GNAME11820(G11820,G11748,G1879);
  nand GNAME11821(G11821,G11820,G11818,G11819);
  or GNAME11822(G11822,G1879,G11748);
  nand GNAME11823(G11823,G11749,G1581);
  nand GNAME11824(G11824,G11823,G11821,G11822);
  or GNAME11825(G11825,G1581,G11749);
  nand GNAME11826(G11826,G11750,G1877);
  nand GNAME11827(G11827,G11826,G11824,G11825);
  or GNAME11828(G11828,G1877,G11750);
  nand GNAME11829(G11829,G11751,G1583);
  nand GNAME11830(G11830,G11829,G11827,G11828);
  or GNAME11831(G11831,G1583,G11751);
  nand GNAME11832(G11832,G11752,G1875);
  nand GNAME11833(G11833,G11832,G11830,G11831);
  or GNAME11834(G11834,G1875,G11752);
  nand GNAME11835(G11835,G11753,G1585);
  nand GNAME11836(G11836,G11835,G11833,G11834);
  or GNAME11837(G11837,G1585,G11753);
  nand GNAME11838(G11838,G11754,G1873);
  nand GNAME11839(G11839,G11838,G11836,G11837);
  or GNAME11840(G11840,G1873,G11754);
  nand GNAME11841(G11841,G11755,G1587);
  nand GNAME11842(G11842,G11841,G11839,G11840);
  or GNAME11843(G11843,G1587,G11755);
  nand GNAME11844(G11844,G11756,G1871);
  nand GNAME11845(G11845,G11844,G11842,G11843);
  or GNAME11846(G11846,G1871,G11756);
  nand GNAME11847(G11847,G11757,G1590);
  nand GNAME11848(G11848,G11847,G11845,G11846);
  or GNAME11849(G11849,G1590,G11757);
  or GNAME11850(G11850,G1868,G11758);
  nand GNAME11851(G11851,G11850,G11848,G11849);
  nand GNAME11852(G11852,G11758,G1868);
  nand GNAME11853(G11853,G11980,G11981);
  and GNAME11854(G11854,G11855,G1308);
  not GNAME11855(G11855,G1340);
  not GNAME11856(G11856,G1307);
  not GNAME11857(G11857,G1338);
  not GNAME11858(G11858,G1305);
  not GNAME11859(G11859,G1336);
  not GNAME11860(G11860,G1303);
  not GNAME11861(G11861,G1334);
  not GNAME11862(G11862,G1301);
  not GNAME11863(G11863,G1332);
  not GNAME11864(G11864,G1299);
  not GNAME11865(G11865,G1330);
  not GNAME11866(G11866,G1297);
  not GNAME11867(G11867,G1328);
  not GNAME11868(G11868,G1295);
  not GNAME11869(G11869,G1326);
  not GNAME11870(G11870,G1293);
  not GNAME11871(G11871,G1324);
  not GNAME11872(G11872,G1291);
  not GNAME11873(G11873,G1322);
  not GNAME11874(G11874,G1289);
  not GNAME11875(G11875,G1320);
  not GNAME11876(G11876,G1287);
  not GNAME11877(G11877,G1318);
  not GNAME11878(G11878,G1285);
  not GNAME11879(G11879,G1316);
  not GNAME11880(G11880,G1283);
  not GNAME11881(G11881,G1314);
  not GNAME11882(G11882,G1281);
  not GNAME11883(G11883,G1312);
  not GNAME11884(G11884,G1279);
  not GNAME11885(G11885,G1310);
  not GNAME11886(G11886,G1277);
  not GNAME11887(G11887,G1309);
  or GNAME11888(G11888,G11854,G1276);
  or GNAME11889(G11889,G1308,G11855);
  nand GNAME11890(G11890,G11856,G1339);
  nand GNAME11891(G11891,G11890,G11888,G11889);
  or GNAME11892(G11892,G1339,G11856);
  nand GNAME11893(G11893,G11857,G1306);
  nand GNAME11894(G11894,G11893,G11891,G11892);
  or GNAME11895(G11895,G1306,G11857);
  nand GNAME11896(G11896,G11858,G1337);
  nand GNAME11897(G11897,G11896,G11894,G11895);
  or GNAME11898(G11898,G1337,G11858);
  nand GNAME11899(G11899,G11859,G1304);
  nand GNAME11900(G11900,G11899,G11897,G11898);
  or GNAME11901(G11901,G1304,G11859);
  nand GNAME11902(G11902,G11860,G1335);
  nand GNAME11903(G11903,G11902,G11900,G11901);
  or GNAME11904(G11904,G1335,G11860);
  nand GNAME11905(G11905,G11861,G1302);
  nand GNAME11906(G11906,G11905,G11903,G11904);
  or GNAME11907(G11907,G1302,G11861);
  nand GNAME11908(G11908,G11862,G1333);
  nand GNAME11909(G11909,G11908,G11906,G11907);
  or GNAME11910(G11910,G1333,G11862);
  nand GNAME11911(G11911,G11863,G1300);
  nand GNAME11912(G11912,G11911,G11909,G11910);
  or GNAME11913(G11913,G1300,G11863);
  nand GNAME11914(G11914,G11864,G1331);
  nand GNAME11915(G11915,G11914,G11912,G11913);
  or GNAME11916(G11916,G1331,G11864);
  nand GNAME11917(G11917,G11865,G1298);
  nand GNAME11918(G11918,G11917,G11915,G11916);
  or GNAME11919(G11919,G1298,G11865);
  nand GNAME11920(G11920,G11866,G1329);
  nand GNAME11921(G11921,G11920,G11918,G11919);
  or GNAME11922(G11922,G1329,G11866);
  nand GNAME11923(G11923,G11867,G1296);
  nand GNAME11924(G11924,G11923,G11921,G11922);
  or GNAME11925(G11925,G1296,G11867);
  nand GNAME11926(G11926,G11868,G1327);
  nand GNAME11927(G11927,G11926,G11924,G11925);
  or GNAME11928(G11928,G1327,G11868);
  nand GNAME11929(G11929,G11869,G1294);
  nand GNAME11930(G11930,G11929,G11927,G11928);
  or GNAME11931(G11931,G1294,G11869);
  nand GNAME11932(G11932,G11870,G1325);
  nand GNAME11933(G11933,G11932,G11930,G11931);
  or GNAME11934(G11934,G1325,G11870);
  nand GNAME11935(G11935,G11871,G1292);
  nand GNAME11936(G11936,G11935,G11933,G11934);
  or GNAME11937(G11937,G1292,G11871);
  nand GNAME11938(G11938,G11872,G1323);
  nand GNAME11939(G11939,G11938,G11936,G11937);
  or GNAME11940(G11940,G1323,G11872);
  nand GNAME11941(G11941,G11873,G1290);
  nand GNAME11942(G11942,G11941,G11939,G11940);
  or GNAME11943(G11943,G1290,G11873);
  nand GNAME11944(G11944,G11874,G1321);
  nand GNAME11945(G11945,G11944,G11942,G11943);
  or GNAME11946(G11946,G1321,G11874);
  nand GNAME11947(G11947,G11875,G1288);
  nand GNAME11948(G11948,G11947,G11945,G11946);
  or GNAME11949(G11949,G1288,G11875);
  nand GNAME11950(G11950,G11876,G1319);
  nand GNAME11951(G11951,G11950,G11948,G11949);
  or GNAME11952(G11952,G1319,G11876);
  nand GNAME11953(G11953,G11877,G1286);
  nand GNAME11954(G11954,G11953,G11951,G11952);
  or GNAME11955(G11955,G1286,G11877);
  nand GNAME11956(G11956,G11878,G1317);
  nand GNAME11957(G11957,G11956,G11954,G11955);
  or GNAME11958(G11958,G1317,G11878);
  nand GNAME11959(G11959,G11879,G1284);
  nand GNAME11960(G11960,G11959,G11957,G11958);
  or GNAME11961(G11961,G1284,G11879);
  nand GNAME11962(G11962,G11880,G1315);
  nand GNAME11963(G11963,G11962,G11960,G11961);
  or GNAME11964(G11964,G1315,G11880);
  nand GNAME11965(G11965,G11881,G1282);
  nand GNAME11966(G11966,G11965,G11963,G11964);
  or GNAME11967(G11967,G1282,G11881);
  nand GNAME11968(G11968,G11882,G1313);
  nand GNAME11969(G11969,G11968,G11966,G11967);
  or GNAME11970(G11970,G1313,G11882);
  nand GNAME11971(G11971,G11883,G1280);
  nand GNAME11972(G11972,G11971,G11969,G11970);
  or GNAME11973(G11973,G1280,G11883);
  nand GNAME11974(G11974,G11884,G1311);
  nand GNAME11975(G11975,G11974,G11972,G11973);
  or GNAME11976(G11976,G1311,G11884);
  nand GNAME11977(G11977,G11885,G1278);
  nand GNAME11978(G11978,G11977,G11975,G11976);
  or GNAME11979(G11979,G1278,G11885);
  nand GNAME11980(G11980,G11983,G11984,G11978,G11979);
  nand GNAME11981(G11981,G11982,G11985,G11986);
  or GNAME11982(G11982,G11886,G11887);
  or GNAME11983(G11983,G1309,G11886);
  or GNAME11984(G11984,G1277,G11887);
  or GNAME11985(G11985,G1275,G1277);
  nand GNAME11986(G11986,G11887,G1275);
  and GNAME11987(G11987,G12006,G12051);
  and GNAME11988(G11988,G12007,G12049);
  and GNAME11989(G11989,G12008,G12048);
  and GNAME11990(G11990,G12009,G12047);
  and GNAME11991(G11991,G12010,G12046);
  and GNAME11992(G11992,G12011,G12045);
  and GNAME11993(G11993,G12012,G12044);
  and GNAME11994(G11994,G12013,G12043);
  and GNAME11995(G11995,G12014,G12042);
  and GNAME11996(G11996,G12015,G12041);
  and GNAME11997(G11997,G12016,G12040);
  and GNAME11998(G11998,G12002,G12039);
  and GNAME11999(G11999,G12003,G12037);
  and GNAME12000(G12000,G12004,G12036);
  and GNAME12001(G12001,G12005,G12035);
  or GNAME12002(G12002,G35974,G35975,G35973);
  or GNAME12003(G12003,G35976,G12002);
  or GNAME12004(G12004,G12058,G35978,G35979);
  or GNAME12005(G12005,G35980,G12004);
  or GNAME12006(G12006,G12054,G35983,G35982);
  or GNAME12007(G12007,G35984,G12006);
  or GNAME12008(G12008,G12082,G35986,G35987);
  or GNAME12009(G12009,G35988,G12008);
  or GNAME12010(G12010,G12078,G35990,G35991);
  or GNAME12011(G12011,G35992,G12010);
  or GNAME12012(G12012,G12072,G35994,G35995);
  or GNAME12013(G12013,G35996,G12012);
  or GNAME12014(G12014,G12068,G35998,G35999);
  or GNAME12015(G12015,G36000,G12014);
  or GNAME12016(G12016,G12015,G36001,G36002);
  nand GNAME12017(G12017,G12073,G12074);
  nand GNAME12018(G12018,G12059,G12060);
  and GNAME12019(G12019,G12050,G12052);
  and GNAME12020(G12020,G12053,G12054);
  and GNAME12021(G12021,G12055,G12056);
  and GNAME12022(G12022,G12057,G12058);
  not GNAME12023(G12023,G36004);
  and GNAME12024(G12024,G12061,G12062);
  and GNAME12025(G12025,G12063,G12064);
  and GNAME12026(G12026,G12065,G12066);
  and GNAME12027(G12027,G12067,G12068);
  and GNAME12028(G12028,G12069,G12070);
  and GNAME12029(G12029,G12071,G12072);
  not GNAME12030(G12030,G35973);
  and GNAME12031(G12031,G12075,G12076);
  and GNAME12032(G12032,G12077,G12078);
  and GNAME12033(G12033,G12079,G12080);
  and GNAME12034(G12034,G12081,G12082);
  nand GNAME12035(G12035,G12004,G35980);
  nand GNAME12036(G12036,G12056,G35979);
  nand GNAME12037(G12037,G12002,G35976);
  or GNAME12038(G12038,G35974,G35973);
  nand GNAME12039(G12039,G12038,G35975);
  nand GNAME12040(G12040,G12064,G36002);
  nand GNAME12041(G12041,G12014,G36000);
  nand GNAME12042(G12042,G12066,G35999);
  nand GNAME12043(G12043,G12012,G35996);
  nand GNAME12044(G12044,G12070,G35995);
  nand GNAME12045(G12045,G12010,G35992);
  nand GNAME12046(G12046,G12076,G35991);
  nand GNAME12047(G12047,G12008,G35988);
  nand GNAME12048(G12048,G12080,G35987);
  nand GNAME12049(G12049,G12006,G35984);
  or GNAME12050(G12050,G35982,G12054);
  nand GNAME12051(G12051,G12050,G35983);
  nand GNAME12052(G12052,G12054,G35982);
  nand GNAME12053(G12053,G12005,G35981);
  or GNAME12054(G12054,G35981,G12005);
  nand GNAME12055(G12055,G12058,G35978);
  or GNAME12056(G12056,G35978,G12058);
  nand GNAME12057(G12057,G12003,G35977);
  or GNAME12058(G12058,G35977,G12003);
  nand GNAME12059(G12059,G12023,G12062);
  or GNAME12060(G12060,G12023,G36003,G12016);
  nand GNAME12061(G12061,G12016,G36003);
  or GNAME12062(G12062,G36003,G12016);
  nand GNAME12063(G12063,G12015,G36001);
  or GNAME12064(G12064,G36001,G12015);
  nand GNAME12065(G12065,G12068,G35998);
  or GNAME12066(G12066,G35998,G12068);
  nand GNAME12067(G12067,G12013,G35997);
  or GNAME12068(G12068,G35997,G12013);
  nand GNAME12069(G12069,G12072,G35994);
  or GNAME12070(G12070,G35994,G12072);
  nand GNAME12071(G12071,G12011,G35993);
  or GNAME12072(G12072,G35993,G12011);
  or GNAME12073(G12073,G35974,G12030);
  nand GNAME12074(G12074,G12030,G35974);
  nand GNAME12075(G12075,G12078,G35990);
  or GNAME12076(G12076,G35990,G12078);
  nand GNAME12077(G12077,G12009,G35989);
  or GNAME12078(G12078,G35989,G12009);
  nand GNAME12079(G12079,G12082,G35986);
  or GNAME12080(G12080,G35986,G12082);
  nand GNAME12081(G12081,G12007,G35985);
  or GNAME12082(G12082,G35985,G12007);
  and GNAME12083(G12083,G12084,G1244);
  not GNAME12084(G12084,G1242);
  not GNAME12085(G12085,G36209);
  and GNAME12086(G12086,G36207,G12121,G36213);
  not GNAME12087(G12087,G36200);
  not GNAME12088(G12088,G36197);
  not GNAME12089(G12089,G36214);
  nor GNAME12090(G12090,G12088,G12085,G12087);
  not GNAME12091(G12091,G36188);
  and GNAME12092(G12092,G36188,G36214,G12090);
  not GNAME12093(G12093,G36206);
  nand GNAME12094(G12094,G12092,G36206);
  and GNAME12095(G12095,G36196,G12210);
  not GNAME12096(G12096,G36191);
  not GNAME12097(G12097,G36210);
  not GNAME12098(G12098,G36193);
  and GNAME12099(G12099,G36210,G12095,G36191);
  not GNAME12100(G12100,G36203);
  not GNAME12101(G12101,G36186);
  and GNAME12102(G12102,G36203,G36193,G12099);
  not GNAME12103(G12103,G36212);
  not GNAME12104(G12104,G36199);
  and GNAME12105(G12105,G36212,G36186,G12102);
  not GNAME12106(G12106,G36201);
  not GNAME12107(G12107,G36208);
  and GNAME12108(G12108,G36201,G36199,G12105);
  not GNAME12109(G12109,G36189);
  not GNAME12110(G12110,G36204);
  and GNAME12111(G12111,G36189,G36208,G12108);
  not GNAME12112(G12112,G36194);
  not GNAME12113(G12113,G36211);
  and GNAME12114(G12114,G36194,G36204,G12111);
  not GNAME12115(G12115,G36192);
  not GNAME12116(G12116,G36202);
  and GNAME12117(G12117,G36192,G36211,G12114);
  not GNAME12118(G12118,G36198);
  and GNAME12119(G12119,G36198,G36202,G12117);
  not GNAME12120(G12120,G36187);
  and GNAME12121(G12121,G12119,G36187);
  not GNAME12122(G12122,G36213);
  not GNAME12123(G12123,G36207);
  nand GNAME12124(G12124,G12160,G12161);
  nand GNAME12125(G12125,G12162,G12163);
  nand GNAME12126(G12126,G12164,G12165);
  nand GNAME12127(G12127,G12166,G12167);
  nand GNAME12128(G12128,G12168,G12169);
  nand GNAME12129(G12129,G12170,G12171);
  nand GNAME12130(G12130,G12172,G12173);
  nand GNAME12131(G12131,G12174,G12175);
  nand GNAME12132(G12132,G12176,G12177);
  nand GNAME12133(G12133,G12178,G12179);
  nand GNAME12134(G12134,G12180,G12181);
  nand GNAME12135(G12135,G12182,G12183);
  nand GNAME12136(G12136,G12184,G12185);
  nand GNAME12137(G12137,G12186,G12187);
  nand GNAME12138(G12138,G12188,G12189);
  nand GNAME12139(G12139,G12190,G12191);
  nand GNAME12140(G12140,G12192,G12193);
  nand GNAME12141(G12141,G12194,G12195);
  nand GNAME12142(G12142,G12196,G12197);
  nand GNAME12143(G12143,G12198,G12199);
  nand GNAME12144(G12144,G12200,G12201);
  nand GNAME12145(G12145,G12202,G12203);
  nand GNAME12146(G12146,G12204,G12205);
  nand GNAME12147(G12147,G12206,G12207);
  nand GNAME12148(G12148,G12208,G12209);
  and GNAME12149(G12149,G12090,G36188);
  nor GNAME12150(G12150,G12085,G12088);
  and GNAME12151(G12151,G12121,G36213);
  and GNAME12152(G12152,G12117,G36198);
  and GNAME12153(G12153,G12114,G36192);
  and GNAME12154(G12154,G12111,G36194);
  and GNAME12155(G12155,G12108,G36189);
  and GNAME12156(G12156,G12105,G36201);
  and GNAME12157(G12157,G12102,G36212);
  and GNAME12158(G12158,G12099,G36203);
  and GNAME12159(G12159,G12095,G36210);
  nand GNAME12160(G12160,G12094,G36196);
  or GNAME12161(G12161,G36196,G12094);
  or GNAME12162(G12162,G12092,G12093);
  nand GNAME12163(G12163,G12093,G12092);
  or GNAME12164(G12164,G12149,G12089);
  nand GNAME12165(G12165,G12089,G12149);
  or GNAME12166(G12166,G12090,G12091);
  nand GNAME12167(G12167,G12091,G12090);
  or GNAME12168(G12168,G12150,G12087);
  nand GNAME12169(G12169,G12087,G12150);
  or GNAME12170(G12170,G36209,G12088);
  or GNAME12171(G12171,G36197,G12085);
  or GNAME12172(G12172,G12151,G12123);
  nand GNAME12173(G12173,G12123,G12151);
  or GNAME12174(G12174,G12121,G12122);
  nand GNAME12175(G12175,G12122,G12121);
  or GNAME12176(G12176,G12119,G12120);
  nand GNAME12177(G12177,G12120,G12119);
  or GNAME12178(G12178,G12152,G12116);
  nand GNAME12179(G12179,G12116,G12152);
  or GNAME12180(G12180,G12117,G12118);
  nand GNAME12181(G12181,G12118,G12117);
  or GNAME12182(G12182,G12153,G12113);
  nand GNAME12183(G12183,G12113,G12153);
  or GNAME12184(G12184,G12114,G12115);
  nand GNAME12185(G12185,G12115,G12114);
  or GNAME12186(G12186,G12154,G12110);
  nand GNAME12187(G12187,G12110,G12154);
  or GNAME12188(G12188,G12111,G12112);
  nand GNAME12189(G12189,G12112,G12111);
  or GNAME12190(G12190,G12155,G12107);
  nand GNAME12191(G12191,G12107,G12155);
  or GNAME12192(G12192,G12108,G12109);
  nand GNAME12193(G12193,G12109,G12108);
  or GNAME12194(G12194,G12156,G12104);
  nand GNAME12195(G12195,G12104,G12156);
  or GNAME12196(G12196,G12105,G12106);
  nand GNAME12197(G12197,G12106,G12105);
  or GNAME12198(G12198,G12157,G12101);
  nand GNAME12199(G12199,G12101,G12157);
  or GNAME12200(G12200,G12102,G12103);
  nand GNAME12201(G12201,G12103,G12102);
  or GNAME12202(G12202,G12158,G12098);
  nand GNAME12203(G12203,G12098,G12158);
  or GNAME12204(G12204,G12099,G12100);
  nand GNAME12205(G12205,G12100,G12099);
  or GNAME12206(G12206,G12159,G12096);
  nand GNAME12207(G12207,G12096,G12159);
  or GNAME12208(G12208,G12095,G12097);
  nand GNAME12209(G12209,G12097,G12095);
  not GNAME12210(G12210,G12094);
  nand GNAME12211(G12211,G12431,G12429);
  nand GNAME12212(G12212,G12432,G12366);
  not GNAME12213(G12213,G1373);
  nor GNAME12214(G12214,G1405,G12213);
  not GNAME12215(G12215,G1372);
  not GNAME12216(G12216,G1403);
  not GNAME12217(G12217,G1371);
  not GNAME12218(G12218,G1402);
  not GNAME12219(G12219,G1370);
  not GNAME12220(G12220,G1401);
  not GNAME12221(G12221,G1369);
  not GNAME12222(G12222,G1400);
  not GNAME12223(G12223,G1368);
  not GNAME12224(G12224,G1399);
  not GNAME12225(G12225,G1367);
  not GNAME12226(G12226,G1398);
  not GNAME12227(G12227,G1366);
  not GNAME12228(G12228,G1397);
  not GNAME12229(G12229,G1365);
  not GNAME12230(G12230,G1396);
  not GNAME12231(G12231,G1364);
  not GNAME12232(G12232,G1395);
  not GNAME12233(G12233,G1363);
  not GNAME12234(G12234,G1394);
  not GNAME12235(G12235,G1362);
  not GNAME12236(G12236,G1393);
  not GNAME12237(G12237,G1361);
  not GNAME12238(G12238,G1392);
  not GNAME12239(G12239,G1360);
  not GNAME12240(G12240,G1391);
  not GNAME12241(G12241,G1359);
  not GNAME12242(G12242,G1390);
  not GNAME12243(G12243,G1358);
  not GNAME12244(G12244,G1389);
  not GNAME12245(G12245,G1357);
  not GNAME12246(G12246,G1388);
  not GNAME12247(G12247,G1356);
  not GNAME12248(G12248,G1387);
  not GNAME12249(G12249,G1355);
  not GNAME12250(G12250,G1386);
  not GNAME12251(G12251,G1354);
  not GNAME12252(G12252,G1385);
  not GNAME12253(G12253,G1353);
  not GNAME12254(G12254,G1384);
  not GNAME12255(G12255,G1352);
  not GNAME12256(G12256,G1383);
  not GNAME12257(G12257,G1351);
  not GNAME12258(G12258,G1382);
  not GNAME12259(G12259,G1350);
  not GNAME12260(G12260,G1381);
  not GNAME12261(G12261,G1349);
  not GNAME12262(G12262,G1380);
  not GNAME12263(G12263,G1348);
  not GNAME12264(G12264,G1379);
  not GNAME12265(G12265,G1347);
  not GNAME12266(G12266,G1378);
  not GNAME12267(G12267,G1346);
  not GNAME12268(G12268,G1377);
  not GNAME12269(G12269,G1345);
  not GNAME12270(G12270,G1376);
  not GNAME12271(G12271,G1344);
  not GNAME12272(G12272,G1343);
  and GNAME12273(G12273,G12426,G12472);
  not GNAME12274(G12274,G1375);
  nand GNAME12275(G12275,G12513,G12514);
  and GNAME12276(G12276,G12433,G12386);
  and GNAME12277(G12277,G12436,G12437);
  and GNAME12278(G12278,G12440,G12441);
  and GNAME12279(G12279,G12444,G12445);
  and GNAME12280(G12280,G12448,G12449);
  and GNAME12281(G12281,G12452,G12453);
  and GNAME12282(G12282,G12456,G12457);
  and GNAME12283(G12283,G12463,G12464);
  and GNAME12284(G12284,G12467,G12468);
  and GNAME12285(G12285,G12471,G12472);
  and GNAME12286(G12286,G12475,G12476);
  and GNAME12287(G12287,G12479,G12480);
  and GNAME12288(G12288,G12483,G12484);
  and GNAME12289(G12289,G12487,G12488);
  and GNAME12290(G12290,G12491,G12492);
  and GNAME12291(G12291,G12495,G12496);
  and GNAME12292(G12292,G12499,G12500);
  and GNAME12293(G12293,G12503,G12504);
  and GNAME12294(G12294,G12507,G12508);
  and GNAME12295(G12295,G12511,G12512);
  and GNAME12296(G12296,G12515,G12516);
  and GNAME12297(G12297,G12519,G12520);
  and GNAME12298(G12298,G12523,G12524);
  and GNAME12299(G12299,G12527,G12528);
  and GNAME12300(G12300,G12531,G12532);
  and GNAME12301(G12301,G12535,G12536);
  and GNAME12302(G12302,G12539,G12540);
  and GNAME12303(G12303,G12543,G12544);
  and GNAME12304(G12304,G12547,G12548);
  and GNAME12305(G12305,G12551,G12552);
  and GNAME12306(G12306,G12383,G12437);
  and GNAME12307(G12307,G12434,G12435);
  and GNAME12308(G12308,G12381,G12441);
  and GNAME12309(G12309,G12438,G12439);
  and GNAME12310(G12310,G12379,G12445);
  and GNAME12311(G12311,G12442,G12443);
  and GNAME12312(G12312,G12377,G12449);
  and GNAME12313(G12313,G12446,G12447);
  and GNAME12314(G12314,G12375,G12453);
  and GNAME12315(G12315,G12450,G12451);
  and GNAME12316(G12316,G12373,G12457);
  and GNAME12317(G12317,G12454,G12455);
  and GNAME12318(G12318,G12371,G12468);
  and GNAME12319(G12319,G12458,G12459);
  not GNAME12320(G12320,G1374);
  not GNAME12321(G12321,G1342);
  and GNAME12322(G12322,G12465,G12466);
  and GNAME12323(G12323,G12368,G12369);
  and GNAME12324(G12324,G12469,G12470);
  and GNAME12325(G12325,G12424,G12476);
  and GNAME12326(G12326,G12473,G12474);
  and GNAME12327(G12327,G12422,G12480);
  and GNAME12328(G12328,G12477,G12478);
  and GNAME12329(G12329,G12420,G12484);
  and GNAME12330(G12330,G12481,G12482);
  and GNAME12331(G12331,G12418,G12488);
  and GNAME12332(G12332,G12485,G12486);
  and GNAME12333(G12333,G12416,G12492);
  and GNAME12334(G12334,G12489,G12490);
  and GNAME12335(G12335,G12414,G12496);
  and GNAME12336(G12336,G12493,G12494);
  and GNAME12337(G12337,G12412,G12500);
  and GNAME12338(G12338,G12497,G12498);
  and GNAME12339(G12339,G12410,G12504);
  and GNAME12340(G12340,G12501,G12502);
  and GNAME12341(G12341,G12408,G12508);
  and GNAME12342(G12342,G12505,G12506);
  and GNAME12343(G12343,G12406,G12516);
  and GNAME12344(G12344,G12509,G12510);
  not GNAME12345(G12345,G1404);
  and GNAME12346(G12346,G12404,G12520);
  and GNAME12347(G12347,G12517,G12518);
  and GNAME12348(G12348,G12402,G12524);
  and GNAME12349(G12349,G12521,G12522);
  and GNAME12350(G12350,G12400,G12528);
  and GNAME12351(G12351,G12525,G12526);
  and GNAME12352(G12352,G12398,G12532);
  and GNAME12353(G12353,G12529,G12530);
  and GNAME12354(G12354,G12396,G12536);
  and GNAME12355(G12355,G12533,G12534);
  and GNAME12356(G12356,G12394,G12540);
  and GNAME12357(G12357,G12537,G12538);
  and GNAME12358(G12358,G12392,G12544);
  and GNAME12359(G12359,G12541,G12542);
  and GNAME12360(G12360,G12390,G12548);
  and GNAME12361(G12361,G12545,G12546);
  and GNAME12362(G12362,G12388,G12552);
  and GNAME12363(G12363,G12549,G12550);
  and GNAME12364(G12364,G12385,G12386);
  and GNAME12365(G12365,G12553,G12554);
  not GNAME12366(G12366,G12214);
  or GNAME12367(G12367,G12214,G1372);
  nand GNAME12368(G12368,G12345,G12367);
  or GNAME12369(G12369,G12366,G12215);
  nor GNAME12370(G12370,G1371,G12216);
  or GNAME12371(G12371,G12323,G12370);
  nor GNAME12372(G12372,G1370,G12218);
  or GNAME12373(G12373,G12318,G12372);
  nor GNAME12374(G12374,G1369,G12220);
  or GNAME12375(G12375,G12316,G12374);
  nor GNAME12376(G12376,G1368,G12222);
  or GNAME12377(G12377,G12314,G12376);
  nor GNAME12378(G12378,G1367,G12224);
  or GNAME12379(G12379,G12312,G12378);
  nor GNAME12380(G12380,G1366,G12226);
  or GNAME12381(G12381,G12310,G12380);
  nor GNAME12382(G12382,G1365,G12228);
  or GNAME12383(G12383,G12308,G12382);
  nor GNAME12384(G12384,G1364,G12230);
  or GNAME12385(G12385,G12306,G12384);
  or GNAME12386(G12386,G1396,G12231);
  nor GNAME12387(G12387,G1363,G12232);
  or GNAME12388(G12388,G12364,G12387);
  nor GNAME12389(G12389,G1362,G12234);
  or GNAME12390(G12390,G12362,G12389);
  nor GNAME12391(G12391,G1361,G12236);
  or GNAME12392(G12392,G12360,G12391);
  nor GNAME12393(G12393,G1360,G12238);
  or GNAME12394(G12394,G12358,G12393);
  nor GNAME12395(G12395,G1359,G12240);
  or GNAME12396(G12396,G12356,G12395);
  nor GNAME12397(G12397,G1358,G12242);
  or GNAME12398(G12398,G12354,G12397);
  nor GNAME12399(G12399,G1357,G12244);
  or GNAME12400(G12400,G12352,G12399);
  nor GNAME12401(G12401,G1356,G12246);
  or GNAME12402(G12402,G12350,G12401);
  nor GNAME12403(G12403,G1355,G12248);
  or GNAME12404(G12404,G12348,G12403);
  nor GNAME12405(G12405,G1354,G12250);
  or GNAME12406(G12406,G12346,G12405);
  nor GNAME12407(G12407,G1353,G12252);
  or GNAME12408(G12408,G12343,G12407);
  nor GNAME12409(G12409,G1352,G12254);
  or GNAME12410(G12410,G12341,G12409);
  nor GNAME12411(G12411,G1351,G12256);
  or GNAME12412(G12412,G12339,G12411);
  nor GNAME12413(G12413,G1350,G12258);
  or GNAME12414(G12414,G12337,G12413);
  nor GNAME12415(G12415,G1349,G12260);
  or GNAME12416(G12416,G12335,G12415);
  nor GNAME12417(G12417,G1348,G12262);
  or GNAME12418(G12418,G12333,G12417);
  nor GNAME12419(G12419,G1347,G12264);
  or GNAME12420(G12420,G12331,G12419);
  nor GNAME12421(G12421,G1346,G12266);
  or GNAME12422(G12422,G12329,G12421);
  nor GNAME12423(G12423,G1345,G12268);
  or GNAME12424(G12424,G12327,G12423);
  nor GNAME12425(G12425,G1344,G12270);
  or GNAME12426(G12426,G12325,G12425);
  nor GNAME12427(G12427,G1343,G12274);
  or GNAME12428(G12428,G12273,G12427);
  nand GNAME12429(G12429,G12462,G12428,G12464);
  nand GNAME12430(G12430,G12464,G12273);
  nand GNAME12431(G12431,G12460,G12461,G12430,G12463);
  nand GNAME12432(G12432,G12213,G1405);
  or GNAME12433(G12433,G1364,G12230);
  nand GNAME12434(G12434,G12276,G12306);
  or GNAME12435(G12435,G12306,G12276);
  or GNAME12436(G12436,G1365,G12228);
  or GNAME12437(G12437,G1397,G12229);
  nand GNAME12438(G12438,G12277,G12308);
  or GNAME12439(G12439,G12308,G12277);
  or GNAME12440(G12440,G1366,G12226);
  or GNAME12441(G12441,G1398,G12227);
  nand GNAME12442(G12442,G12278,G12310);
  or GNAME12443(G12443,G12310,G12278);
  or GNAME12444(G12444,G1367,G12224);
  or GNAME12445(G12445,G1399,G12225);
  nand GNAME12446(G12446,G12279,G12312);
  or GNAME12447(G12447,G12312,G12279);
  or GNAME12448(G12448,G1368,G12222);
  or GNAME12449(G12449,G1400,G12223);
  nand GNAME12450(G12450,G12280,G12314);
  or GNAME12451(G12451,G12314,G12280);
  or GNAME12452(G12452,G1369,G12220);
  or GNAME12453(G12453,G1401,G12221);
  nand GNAME12454(G12454,G12281,G12316);
  or GNAME12455(G12455,G12316,G12281);
  or GNAME12456(G12456,G1370,G12218);
  or GNAME12457(G12457,G1402,G12219);
  nand GNAME12458(G12458,G12282,G12318);
  or GNAME12459(G12459,G12318,G12282);
  or GNAME12460(G12460,G1342,G12320);
  or GNAME12461(G12461,G1374,G12321);
  nand GNAME12462(G12462,G12460,G12461);
  or GNAME12463(G12463,G1343,G12274);
  or GNAME12464(G12464,G1375,G12272);
  nand GNAME12465(G12465,G12273,G12283);
  or GNAME12466(G12466,G12273,G12283);
  or GNAME12467(G12467,G1371,G12216);
  or GNAME12468(G12468,G1403,G12217);
  nand GNAME12469(G12469,G12284,G12323);
  or GNAME12470(G12470,G12323,G12284);
  or GNAME12471(G12471,G1344,G12270);
  or GNAME12472(G12472,G1376,G12271);
  nand GNAME12473(G12473,G12285,G12325);
  or GNAME12474(G12474,G12325,G12285);
  or GNAME12475(G12475,G1345,G12268);
  or GNAME12476(G12476,G1377,G12269);
  nand GNAME12477(G12477,G12286,G12327);
  or GNAME12478(G12478,G12327,G12286);
  or GNAME12479(G12479,G1346,G12266);
  or GNAME12480(G12480,G1378,G12267);
  nand GNAME12481(G12481,G12287,G12329);
  or GNAME12482(G12482,G12329,G12287);
  or GNAME12483(G12483,G1347,G12264);
  or GNAME12484(G12484,G1379,G12265);
  nand GNAME12485(G12485,G12288,G12331);
  or GNAME12486(G12486,G12331,G12288);
  or GNAME12487(G12487,G1348,G12262);
  or GNAME12488(G12488,G1380,G12263);
  nand GNAME12489(G12489,G12289,G12333);
  or GNAME12490(G12490,G12333,G12289);
  or GNAME12491(G12491,G1349,G12260);
  or GNAME12492(G12492,G1381,G12261);
  nand GNAME12493(G12493,G12290,G12335);
  or GNAME12494(G12494,G12335,G12290);
  or GNAME12495(G12495,G1350,G12258);
  or GNAME12496(G12496,G1382,G12259);
  nand GNAME12497(G12497,G12291,G12337);
  or GNAME12498(G12498,G12337,G12291);
  or GNAME12499(G12499,G1351,G12256);
  or GNAME12500(G12500,G1383,G12257);
  nand GNAME12501(G12501,G12292,G12339);
  or GNAME12502(G12502,G12339,G12292);
  or GNAME12503(G12503,G1352,G12254);
  or GNAME12504(G12504,G1384,G12255);
  nand GNAME12505(G12505,G12293,G12341);
  or GNAME12506(G12506,G12341,G12293);
  or GNAME12507(G12507,G1353,G12252);
  or GNAME12508(G12508,G1385,G12253);
  nand GNAME12509(G12509,G12294,G12343);
  or GNAME12510(G12510,G12343,G12294);
  or GNAME12511(G12511,G1372,G12345);
  or GNAME12512(G12512,G1404,G12215);
  nand GNAME12513(G12513,G12214,G12295);
  or GNAME12514(G12514,G12214,G12295);
  or GNAME12515(G12515,G1354,G12250);
  or GNAME12516(G12516,G1386,G12251);
  nand GNAME12517(G12517,G12296,G12346);
  or GNAME12518(G12518,G12346,G12296);
  or GNAME12519(G12519,G1355,G12248);
  or GNAME12520(G12520,G1387,G12249);
  nand GNAME12521(G12521,G12297,G12348);
  or GNAME12522(G12522,G12348,G12297);
  or GNAME12523(G12523,G1356,G12246);
  or GNAME12524(G12524,G1388,G12247);
  nand GNAME12525(G12525,G12298,G12350);
  or GNAME12526(G12526,G12350,G12298);
  or GNAME12527(G12527,G1357,G12244);
  or GNAME12528(G12528,G1389,G12245);
  nand GNAME12529(G12529,G12299,G12352);
  or GNAME12530(G12530,G12352,G12299);
  or GNAME12531(G12531,G1358,G12242);
  or GNAME12532(G12532,G1390,G12243);
  nand GNAME12533(G12533,G12300,G12354);
  or GNAME12534(G12534,G12354,G12300);
  or GNAME12535(G12535,G1359,G12240);
  or GNAME12536(G12536,G1391,G12241);
  nand GNAME12537(G12537,G12301,G12356);
  or GNAME12538(G12538,G12356,G12301);
  or GNAME12539(G12539,G1360,G12238);
  or GNAME12540(G12540,G1392,G12239);
  nand GNAME12541(G12541,G12302,G12358);
  or GNAME12542(G12542,G12358,G12302);
  or GNAME12543(G12543,G1361,G12236);
  or GNAME12544(G12544,G1393,G12237);
  nand GNAME12545(G12545,G12303,G12360);
  or GNAME12546(G12546,G12360,G12303);
  or GNAME12547(G12547,G1362,G12234);
  or GNAME12548(G12548,G1394,G12235);
  nand GNAME12549(G12549,G12304,G12362);
  or GNAME12550(G12550,G12362,G12304);
  or GNAME12551(G12551,G1363,G12232);
  or GNAME12552(G12552,G1395,G12233);
  nand GNAME12553(G12553,G12305,G12364);
  or GNAME12554(G12554,G12364,G12305);
  and GNAME12555(G12555,G12833,G12834);
  and GNAME12556(G12556,G12829,G12831);
  and GNAME12557(G12557,G12825,G12826);
  and GNAME12558(G12558,G12822,G12823);
  and GNAME12559(G12559,G12818,G12820);
  and GNAME12560(G12560,G12815,G12817);
  and GNAME12561(G12561,G12727,G12729);
  and GNAME12562(G12562,G12721,G12722);
  and GNAME12563(G12563,G12717,G12719);
  not GNAME12564(G12564,G4174);
  not GNAME12565(G12565,G4239);
  not GNAME12566(G12566,G4238);
  not GNAME12567(G12567,G4237);
  not GNAME12568(G12568,G4236);
  not GNAME12569(G12569,G4235);
  not GNAME12570(G12570,G4234);
  not GNAME12571(G12571,G4233);
  not GNAME12572(G12572,G4232);
  not GNAME12573(G12573,G4231);
  not GNAME12574(G12574,G4230);
  and GNAME12575(G12575,G12715,G12690);
  or GNAME12576(G12576,G12687,G12575);
  not GNAME12577(G12577,G4208);
  not GNAME12578(G12578,G4229);
  not GNAME12579(G12579,G4228);
  not GNAME12580(G12580,G4227);
  not GNAME12581(G12581,G4226);
  not GNAME12582(G12582,G4225);
  not GNAME12583(G12583,G4224);
  not GNAME12584(G12584,G4223);
  not GNAME12585(G12585,G4222);
  not GNAME12586(G12586,G4221);
  not GNAME12587(G12587,G4220);
  not GNAME12588(G12588,G4219);
  not GNAME12589(G12589,G4218);
  not GNAME12590(G12590,G4217);
  not GNAME12591(G12591,G4216);
  not GNAME12592(G12592,G4215);
  not GNAME12593(G12593,G4214);
  not GNAME12594(G12594,G4213);
  not GNAME12595(G12595,G4212);
  not GNAME12596(G12596,G4211);
  not GNAME12597(G12597,G4210);
  nor GNAME12598(G12598,G12811,G12599);
  and GNAME12599(G12599,G12810,G12809);
  and GNAME12600(G12600,G12725,G12696);
  or GNAME12601(G12601,G12693,G12600);
  and GNAME12602(G12602,G12751,G12750);
  nor GNAME12603(G12603,G12752,G12602);
  and GNAME12604(G12604,G12827,G12712);
  or GNAME12605(G12605,G12736,G12604);
  and GNAME12606(G12606,G12873,G12874);
  and GNAME12607(G12607,G12878,G12879);
  and GNAME12608(G12608,G12883,G12884);
  nand GNAME12609(G12609,G12995,G12996);
  nand GNAME12610(G12610,G12885,G12886);
  nand GNAME12611(G12611,G12887,G12888);
  nand GNAME12612(G12612,G12889,G12890);
  nand GNAME12613(G12613,G12891,G12892);
  nand GNAME12614(G12614,G12959,G12960);
  nand GNAME12615(G12615,G12961,G12962);
  nand GNAME12616(G12616,G12963,G12964);
  nand GNAME12617(G12617,G12965,G12966);
  nand GNAME12618(G12618,G12967,G12968);
  nand GNAME12619(G12619,G12969,G12970);
  nand GNAME12620(G12620,G12971,G12972);
  nand GNAME12621(G12621,G12973,G12974);
  nand GNAME12622(G12622,G12975,G12976);
  nand GNAME12623(G12623,G12977,G12978);
  nand GNAME12624(G12624,G12979,G12980);
  nand GNAME12625(G12625,G12981,G12982);
  nand GNAME12626(G12626,G12983,G12984);
  nand GNAME12627(G12627,G12985,G12986);
  nand GNAME12628(G12628,G12987,G12988);
  nand GNAME12629(G12629,G12989,G12990);
  nand GNAME12630(G12630,G12991,G12992);
  nand GNAME12631(G12631,G12993,G12994);
  not GNAME12632(G12632,G4196);
  not GNAME12633(G12633,G4198);
  not GNAME12634(G12634,G4199);
  not GNAME12635(G12635,G4200);
  not GNAME12636(G12636,G4202);
  not GNAME12637(G12637,G4203);
  not GNAME12638(G12638,G4204);
  nand GNAME12639(G12639,G12707,G12686);
  nand GNAME12640(G12640,G12713,G12684);
  nand GNAME12641(G12641,G12701,G12692);
  not GNAME12642(G12642,G4176);
  not GNAME12643(G12643,G4175);
  not GNAME12644(G12644,G4190);
  not GNAME12645(G12645,G4191);
  not GNAME12646(G12646,G4194);
  not GNAME12647(G12647,G4195);
  not GNAME12648(G12648,G4193);
  not GNAME12649(G12649,G4192);
  not GNAME12650(G12650,G4189);
  not GNAME12651(G12651,G4188);
  not GNAME12652(G12652,G4187);
  not GNAME12653(G12653,G4186);
  not GNAME12654(G12654,G4185);
  not GNAME12655(G12655,G4184);
  not GNAME12656(G12656,G4183);
  not GNAME12657(G12657,G4182);
  not GNAME12658(G12658,G4181);
  not GNAME12659(G12659,G4180);
  not GNAME12660(G12660,G4179);
  not GNAME12661(G12661,G4178);
  not GNAME12662(G12662,G4177);
  nand GNAME12663(G12663,G12806,G12805);
  nand GNAME12664(G12664,G12802,G12801);
  nand GNAME12665(G12665,G12798,G12797);
  nand GNAME12666(G12666,G12794,G12793);
  nand GNAME12667(G12667,G12790,G12789);
  nand GNAME12668(G12668,G12786,G12785);
  nand GNAME12669(G12669,G12782,G12781);
  nand GNAME12670(G12670,G12778,G12777);
  nand GNAME12671(G12671,G12774,G12773);
  nand GNAME12672(G12672,G12770,G12769);
  nand GNAME12673(G12673,G12723,G12683);
  nand GNAME12674(G12674,G12766,G12765);
  nand GNAME12675(G12675,G12762,G12761);
  nand GNAME12676(G12676,G12758,G12757);
  nand GNAME12677(G12677,G12754,G12732);
  or GNAME12678(G12678,G12603,G12733);
  nand GNAME12679(G12679,G12747,G12746);
  nand GNAME12680(G12680,G12743,G12735);
  nand GNAME12681(G12681,G12697,G12683);
  or GNAME12682(G12682,G12608,G12573);
  or GNAME12683(G12683,G12606,G12565);
  or GNAME12684(G12684,G12607,G12569);
  nand GNAME12685(G12685,G12572,G12861,G12862);
  nand GNAME12686(G12686,G12882,G4232);
  and GNAME12687(G12687,G12571,G12863,G12864);
  nand GNAME12688(G12688,G12881,G4233);
  nand GNAME12689(G12689,G12570,G12865,G12866);
  nand GNAME12690(G12690,G12880,G4234);
  nand GNAME12691(G12691,G12568,G12867,G12868);
  nand GNAME12692(G12692,G12877,G4236);
  and GNAME12693(G12693,G12567,G12869,G12870);
  nand GNAME12694(G12694,G12876,G4237);
  nand GNAME12695(G12695,G12566,G12871,G12872);
  nand GNAME12696(G12696,G12875,G4238);
  nand GNAME12697(G12697,G12565,G12606);
  nand GNAME12698(G12698,G12725,G12696);
  nand GNAME12699(G12699,G12998,G12698);
  nand GNAME12700(G12700,G12699,G12694);
  nand GNAME12701(G12701,G12691,G12700);
  not GNAME12702(G12702,G12641);
  nand GNAME12703(G12703,G12569,G12607);
  nand GNAME12704(G12704,G12715,G12690);
  nand GNAME12705(G12705,G12997,G12704);
  nand GNAME12706(G12706,G12705,G12688);
  nand GNAME12707(G12707,G12685,G12706);
  not GNAME12708(G12708,G12639);
  nand GNAME12709(G12709,G12573,G12608);
  not GNAME12710(G12710,G12739);
  nand GNAME12711(G12711,G12574,G12858,G12859);
  nand GNAME12712(G12712,G12860,G4230);
  nand GNAME12713(G12713,G12641,G12703);
  not GNAME12714(G12714,G12640);
  nand GNAME12715(G12715,G12689,G12640);
  nand GNAME12716(G12716,G12688,G12576);
  nand GNAME12717(G12717,G12716,G12685,G12686);
  nand GNAME12718(G12718,G12685,G12686);
  nand GNAME12719(G12719,G12718,G12688,G12576);
  or GNAME12720(G12720,G12687,G13000);
  nand GNAME12721(G12721,G12720,G12575);
  or GNAME12722(G12722,G13000,G12576);
  nand GNAME12723(G12723,G12697,G4174);
  not GNAME12724(G12724,G12673);
  nand GNAME12725(G12725,G12695,G12673);
  nand GNAME12726(G12726,G12694,G12601);
  nand GNAME12727(G12727,G12726,G12691,G12692);
  nand GNAME12728(G12728,G12691,G12692);
  nand GNAME12729(G12729,G12728,G12694,G12601);
  and GNAME12730(G12730,G12896,G4208);
  nand GNAME12731(G12731,G12583,G12899,G12900);
  nand GNAME12732(G12732,G12916,G4224);
  and GNAME12733(G12733,G12915,G4225);
  nand GNAME12734(G12734,G12579,G12903,G12904);
  nand GNAME12735(G12735,G12908,G4228);
  and GNAME12736(G12736,G12578,G12905,G12906);
  nand GNAME12737(G12737,G12907,G4229);
  nand GNAME12738(G12738,G12639,G12709);
  nand GNAME12739(G12739,G12738,G12682);
  nand GNAME12740(G12740,G12827,G12712);
  nand GNAME12741(G12741,G12999,G12740);
  nand GNAME12742(G12742,G12741,G12737);
  nand GNAME12743(G12743,G12734,G12742);
  not GNAME12744(G12744,G12680);
  nand GNAME12745(G12745,G12580,G12909,G12910);
  nand GNAME12746(G12746,G12911,G4227);
  nand GNAME12747(G12747,G12680,G12745);
  not GNAME12748(G12748,G12679);
  nand GNAME12749(G12749,G12581,G12912,G12913);
  nand GNAME12750(G12750,G12914,G4226);
  nand GNAME12751(G12751,G12679,G12749);
  and GNAME12752(G12752,G12582,G12901,G12902);
  not GNAME12753(G12753,G12678);
  nand GNAME12754(G12754,G12731,G12678);
  not GNAME12755(G12755,G12677);
  nand GNAME12756(G12756,G12584,G12917,G12918);
  nand GNAME12757(G12757,G12919,G4223);
  nand GNAME12758(G12758,G12677,G12756);
  not GNAME12759(G12759,G12676);
  nand GNAME12760(G12760,G12585,G12920,G12921);
  nand GNAME12761(G12761,G12922,G4222);
  nand GNAME12762(G12762,G12676,G12760);
  not GNAME12763(G12763,G12675);
  nand GNAME12764(G12764,G12586,G12923,G12924);
  nand GNAME12765(G12765,G12925,G4221);
  nand GNAME12766(G12766,G12675,G12764);
  not GNAME12767(G12767,G12674);
  nand GNAME12768(G12768,G12587,G12926,G12927);
  nand GNAME12769(G12769,G12928,G4220);
  nand GNAME12770(G12770,G12674,G12768);
  not GNAME12771(G12771,G12672);
  nand GNAME12772(G12772,G12588,G12929,G12930);
  nand GNAME12773(G12773,G12931,G4219);
  nand GNAME12774(G12774,G12672,G12772);
  not GNAME12775(G12775,G12671);
  nand GNAME12776(G12776,G12589,G12932,G12933);
  nand GNAME12777(G12777,G12934,G4218);
  nand GNAME12778(G12778,G12671,G12776);
  not GNAME12779(G12779,G12670);
  nand GNAME12780(G12780,G12590,G12935,G12936);
  nand GNAME12781(G12781,G12937,G4217);
  nand GNAME12782(G12782,G12670,G12780);
  not GNAME12783(G12783,G12669);
  nand GNAME12784(G12784,G12591,G12938,G12939);
  nand GNAME12785(G12785,G12940,G4216);
  nand GNAME12786(G12786,G12669,G12784);
  not GNAME12787(G12787,G12668);
  nand GNAME12788(G12788,G12592,G12941,G12942);
  nand GNAME12789(G12789,G12943,G4215);
  nand GNAME12790(G12790,G12668,G12788);
  not GNAME12791(G12791,G12667);
  nand GNAME12792(G12792,G12593,G12944,G12945);
  nand GNAME12793(G12793,G12946,G4214);
  nand GNAME12794(G12794,G12667,G12792);
  not GNAME12795(G12795,G12666);
  nand GNAME12796(G12796,G12594,G12947,G12948);
  nand GNAME12797(G12797,G12949,G4213);
  nand GNAME12798(G12798,G12666,G12796);
  not GNAME12799(G12799,G12665);
  nand GNAME12800(G12800,G12595,G12950,G12951);
  nand GNAME12801(G12801,G12952,G4212);
  nand GNAME12802(G12802,G12665,G12800);
  not GNAME12803(G12803,G12664);
  nand GNAME12804(G12804,G12596,G12953,G12954);
  nand GNAME12805(G12805,G12955,G4211);
  nand GNAME12806(G12806,G12664,G12804);
  not GNAME12807(G12807,G12663);
  nand GNAME12808(G12808,G12597,G12956,G12957);
  nand GNAME12809(G12809,G12958,G4210);
  nand GNAME12810(G12810,G12663,G12808);
  and GNAME12811(G12811,G12577,G12897,G12898);
  or GNAME12812(G12812,G12730,G12598);
  nand GNAME12813(G12813,G12812,G4206);
  or GNAME12814(G12814,G12598,G4206,G12730);
  nand GNAME12815(G12815,G12895,G12813,G12814);
  nand GNAME12816(G12816,G12813,G12814);
  nand GNAME12817(G12817,G12816,G12893,G12894);
  or GNAME12818(G12818,G12730,G13001);
  or GNAME12819(G12819,G12730,G12811);
  nand GNAME12820(G12820,G12819,G12599);
  or GNAME12821(G12821,G12693,G13002);
  nand GNAME12822(G12822,G12821,G12600);
  or GNAME12823(G12823,G13002,G12601);
  or GNAME12824(G12824,G12733,G12752);
  nand GNAME12825(G12825,G12824,G12602);
  or GNAME12826(G12826,G12733,G13003);
  nand GNAME12827(G12827,G12739,G12711);
  nand GNAME12828(G12828,G12737,G12605);
  nand GNAME12829(G12829,G12828,G12734,G12735);
  nand GNAME12830(G12830,G12734,G12735);
  nand GNAME12831(G12831,G12830,G12737,G12605);
  or GNAME12832(G12832,G12736,G13004);
  nand GNAME12833(G12833,G12832,G12604);
  or GNAME12834(G12834,G13004,G12605);
  not GNAME12835(G12835,G12681);
  nand GNAME12836(G12836,G12711,G12712);
  nand GNAME12837(G12837,G12682,G12709);
  nand GNAME12838(G12838,G12689,G12690);
  nand GNAME12839(G12839,G12684,G12703);
  nand GNAME12840(G12840,G12808,G12809);
  nand GNAME12841(G12841,G12804,G12805);
  nand GNAME12842(G12842,G12800,G12801);
  nand GNAME12843(G12843,G12796,G12797);
  nand GNAME12844(G12844,G12792,G12793);
  nand GNAME12845(G12845,G12788,G12789);
  nand GNAME12846(G12846,G12784,G12785);
  nand GNAME12847(G12847,G12780,G12781);
  nand GNAME12848(G12848,G12776,G12777);
  nand GNAME12849(G12849,G12772,G12773);
  nand GNAME12850(G12850,G12695,G12696);
  nand GNAME12851(G12851,G12768,G12769);
  nand GNAME12852(G12852,G12764,G12765);
  nand GNAME12853(G12853,G12760,G12761);
  nand GNAME12854(G12854,G12756,G12757);
  nand GNAME12855(G12855,G12731,G12732);
  nand GNAME12856(G12856,G12749,G12750);
  nand GNAME12857(G12857,G12745,G12746);
  nand GNAME12858(G12858,G12632,G4174);
  nand GNAME12859(G12859,G12564,G4196);
  nand GNAME12860(G12860,G12858,G12859);
  nand GNAME12861(G12861,G12633,G4174);
  nand GNAME12862(G12862,G12564,G4198);
  nand GNAME12863(G12863,G12634,G4174);
  nand GNAME12864(G12864,G12564,G4199);
  nand GNAME12865(G12865,G12635,G4174);
  nand GNAME12866(G12866,G12564,G4200);
  nand GNAME12867(G12867,G12636,G4174);
  nand GNAME12868(G12868,G12564,G4202);
  nand GNAME12869(G12869,G12637,G4174);
  nand GNAME12870(G12870,G12564,G4203);
  nand GNAME12871(G12871,G12638,G4174);
  nand GNAME12872(G12872,G12564,G4204);
  or GNAME12873(G12873,G4205,G12564);
  nand GNAME12874(G12874,G12564,G4205);
  nand GNAME12875(G12875,G12871,G12872);
  nand GNAME12876(G12876,G12869,G12870);
  nand GNAME12877(G12877,G12867,G12868);
  or GNAME12878(G12878,G4201,G12564);
  nand GNAME12879(G12879,G12564,G4201);
  nand GNAME12880(G12880,G12865,G12866);
  nand GNAME12881(G12881,G12863,G12864);
  nand GNAME12882(G12882,G12861,G12862);
  or GNAME12883(G12883,G4197,G12564);
  nand GNAME12884(G12884,G12564,G4197);
  nand GNAME12885(G12885,G12739,G12836);
  nand GNAME12886(G12886,G12710,G12711,G12712);
  nand GNAME12887(G12887,G12639,G12837);
  nand GNAME12888(G12888,G12708,G12682,G12709);
  nand GNAME12889(G12889,G12640,G12838);
  nand GNAME12890(G12890,G12714,G12689,G12690);
  nand GNAME12891(G12891,G12641,G12839);
  nand GNAME12892(G12892,G12702,G12684,G12703);
  nand GNAME12893(G12893,G12642,G4174);
  nand GNAME12894(G12894,G12564,G4176);
  nand GNAME12895(G12895,G12893,G12894);
  nand GNAME12896(G12896,G12897,G12898);
  nand GNAME12897(G12897,G12643,G4174);
  nand GNAME12898(G12898,G12564,G4175);
  nand GNAME12899(G12899,G12644,G4174);
  nand GNAME12900(G12900,G12564,G4190);
  nand GNAME12901(G12901,G12645,G4174);
  nand GNAME12902(G12902,G12564,G4191);
  nand GNAME12903(G12903,G12646,G4174);
  nand GNAME12904(G12904,G12564,G4194);
  nand GNAME12905(G12905,G12647,G4174);
  nand GNAME12906(G12906,G12564,G4195);
  nand GNAME12907(G12907,G12905,G12906);
  nand GNAME12908(G12908,G12903,G12904);
  nand GNAME12909(G12909,G12648,G4174);
  nand GNAME12910(G12910,G12564,G4193);
  nand GNAME12911(G12911,G12909,G12910);
  nand GNAME12912(G12912,G12649,G4174);
  nand GNAME12913(G12913,G12564,G4192);
  nand GNAME12914(G12914,G12912,G12913);
  nand GNAME12915(G12915,G12901,G12902);
  nand GNAME12916(G12916,G12899,G12900);
  nand GNAME12917(G12917,G12650,G4174);
  nand GNAME12918(G12918,G12564,G4189);
  nand GNAME12919(G12919,G12917,G12918);
  nand GNAME12920(G12920,G12651,G4174);
  nand GNAME12921(G12921,G12564,G4188);
  nand GNAME12922(G12922,G12920,G12921);
  nand GNAME12923(G12923,G12652,G4174);
  nand GNAME12924(G12924,G12564,G4187);
  nand GNAME12925(G12925,G12923,G12924);
  nand GNAME12926(G12926,G12653,G4174);
  nand GNAME12927(G12927,G12564,G4186);
  nand GNAME12928(G12928,G12926,G12927);
  nand GNAME12929(G12929,G12654,G4174);
  nand GNAME12930(G12930,G12564,G4185);
  nand GNAME12931(G12931,G12929,G12930);
  nand GNAME12932(G12932,G12655,G4174);
  nand GNAME12933(G12933,G12564,G4184);
  nand GNAME12934(G12934,G12932,G12933);
  nand GNAME12935(G12935,G12656,G4174);
  nand GNAME12936(G12936,G12564,G4183);
  nand GNAME12937(G12937,G12935,G12936);
  nand GNAME12938(G12938,G12657,G4174);
  nand GNAME12939(G12939,G12564,G4182);
  nand GNAME12940(G12940,G12938,G12939);
  nand GNAME12941(G12941,G12658,G4174);
  nand GNAME12942(G12942,G12564,G4181);
  nand GNAME12943(G12943,G12941,G12942);
  nand GNAME12944(G12944,G12659,G4174);
  nand GNAME12945(G12945,G12564,G4180);
  nand GNAME12946(G12946,G12944,G12945);
  nand GNAME12947(G12947,G12660,G4174);
  nand GNAME12948(G12948,G12564,G4179);
  nand GNAME12949(G12949,G12947,G12948);
  nand GNAME12950(G12950,G12661,G4174);
  nand GNAME12951(G12951,G12564,G4178);
  nand GNAME12952(G12952,G12950,G12951);
  nand GNAME12953(G12953,G12662,G4174);
  nand GNAME12954(G12954,G12564,G4177);
  nand GNAME12955(G12955,G12953,G12954);
  nand GNAME12956(G12956,G12642,G4174);
  nand GNAME12957(G12957,G12564,G4176);
  nand GNAME12958(G12958,G12956,G12957);
  nand GNAME12959(G12959,G12663,G12840);
  nand GNAME12960(G12960,G12807,G12808,G12809);
  nand GNAME12961(G12961,G12664,G12841);
  nand GNAME12962(G12962,G12803,G12804,G12805);
  nand GNAME12963(G12963,G12665,G12842);
  nand GNAME12964(G12964,G12799,G12800,G12801);
  nand GNAME12965(G12965,G12666,G12843);
  nand GNAME12966(G12966,G12795,G12796,G12797);
  nand GNAME12967(G12967,G12667,G12844);
  nand GNAME12968(G12968,G12791,G12792,G12793);
  nand GNAME12969(G12969,G12668,G12845);
  nand GNAME12970(G12970,G12787,G12788,G12789);
  nand GNAME12971(G12971,G12669,G12846);
  nand GNAME12972(G12972,G12783,G12784,G12785);
  nand GNAME12973(G12973,G12670,G12847);
  nand GNAME12974(G12974,G12779,G12780,G12781);
  nand GNAME12975(G12975,G12671,G12848);
  nand GNAME12976(G12976,G12775,G12776,G12777);
  nand GNAME12977(G12977,G12672,G12849);
  nand GNAME12978(G12978,G12771,G12772,G12773);
  nand GNAME12979(G12979,G12673,G12850);
  nand GNAME12980(G12980,G12724,G12695,G12696);
  nand GNAME12981(G12981,G12674,G12851);
  nand GNAME12982(G12982,G12767,G12768,G12769);
  nand GNAME12983(G12983,G12675,G12852);
  nand GNAME12984(G12984,G12763,G12764,G12765);
  nand GNAME12985(G12985,G12676,G12853);
  nand GNAME12986(G12986,G12759,G12760,G12761);
  nand GNAME12987(G12987,G12677,G12854);
  nand GNAME12988(G12988,G12755,G12756,G12757);
  nand GNAME12989(G12989,G12678,G12855);
  nand GNAME12990(G12990,G12753,G12731,G12732);
  nand GNAME12991(G12991,G12679,G12856);
  nand GNAME12992(G12992,G12748,G12749,G12750);
  nand GNAME12993(G12993,G12680,G12857);
  nand GNAME12994(G12994,G12744,G12745,G12746);
  nand GNAME12995(G12995,G12681,G4174);
  nand GNAME12996(G12996,G12564,G12835);
  not GNAME12997(G12997,G12687);
  not GNAME12998(G12998,G12693);
  not GNAME12999(G12999,G12736);
  not GNAME13000(G13000,G12688);
  not GNAME13001(G13001,G12598);
  not GNAME13002(G13002,G12694);
  not GNAME13003(G13003,G12603);
  not GNAME13004(G13004,G12737);
  nand GNAME13005(G13005,G13132,G13133);
  and GNAME13006(G13006,G13007,G4273);
  not GNAME13007(G13007,G4305);
  not GNAME13008(G13008,G4272);
  not GNAME13009(G13009,G4303);
  not GNAME13010(G13010,G4270);
  not GNAME13011(G13011,G4301);
  not GNAME13012(G13012,G4268);
  not GNAME13013(G13013,G4299);
  not GNAME13014(G13014,G4266);
  not GNAME13015(G13015,G4297);
  not GNAME13016(G13016,G4264);
  not GNAME13017(G13017,G4295);
  not GNAME13018(G13018,G4262);
  not GNAME13019(G13019,G4293);
  not GNAME13020(G13020,G4260);
  not GNAME13021(G13021,G4291);
  not GNAME13022(G13022,G4258);
  not GNAME13023(G13023,G4289);
  not GNAME13024(G13024,G4256);
  not GNAME13025(G13025,G4287);
  not GNAME13026(G13026,G4254);
  not GNAME13027(G13027,G4285);
  not GNAME13028(G13028,G4252);
  not GNAME13029(G13029,G4283);
  not GNAME13030(G13030,G4250);
  not GNAME13031(G13031,G4281);
  not GNAME13032(G13032,G4248);
  not GNAME13033(G13033,G4279);
  not GNAME13034(G13034,G4246);
  not GNAME13035(G13035,G4277);
  not GNAME13036(G13036,G4244);
  not GNAME13037(G13037,G4275);
  not GNAME13038(G13038,G4242);
  not GNAME13039(G13039,G4274);
  or GNAME13040(G13040,G13006,G4241);
  or GNAME13041(G13041,G4273,G13007);
  nand GNAME13042(G13042,G13008,G4304);
  nand GNAME13043(G13043,G13042,G13040,G13041);
  or GNAME13044(G13044,G4304,G13008);
  nand GNAME13045(G13045,G13009,G4271);
  nand GNAME13046(G13046,G13045,G13043,G13044);
  or GNAME13047(G13047,G4271,G13009);
  nand GNAME13048(G13048,G13010,G4302);
  nand GNAME13049(G13049,G13048,G13046,G13047);
  or GNAME13050(G13050,G4302,G13010);
  nand GNAME13051(G13051,G13011,G4269);
  nand GNAME13052(G13052,G13051,G13049,G13050);
  or GNAME13053(G13053,G4269,G13011);
  nand GNAME13054(G13054,G13012,G4300);
  nand GNAME13055(G13055,G13054,G13052,G13053);
  or GNAME13056(G13056,G4300,G13012);
  nand GNAME13057(G13057,G13013,G4267);
  nand GNAME13058(G13058,G13057,G13055,G13056);
  or GNAME13059(G13059,G4267,G13013);
  nand GNAME13060(G13060,G13014,G4298);
  nand GNAME13061(G13061,G13060,G13058,G13059);
  or GNAME13062(G13062,G4298,G13014);
  nand GNAME13063(G13063,G13015,G4265);
  nand GNAME13064(G13064,G13063,G13061,G13062);
  or GNAME13065(G13065,G4265,G13015);
  nand GNAME13066(G13066,G13016,G4296);
  nand GNAME13067(G13067,G13066,G13064,G13065);
  or GNAME13068(G13068,G4296,G13016);
  nand GNAME13069(G13069,G13017,G4263);
  nand GNAME13070(G13070,G13069,G13067,G13068);
  or GNAME13071(G13071,G4263,G13017);
  nand GNAME13072(G13072,G13018,G4294);
  nand GNAME13073(G13073,G13072,G13070,G13071);
  or GNAME13074(G13074,G4294,G13018);
  nand GNAME13075(G13075,G13019,G4261);
  nand GNAME13076(G13076,G13075,G13073,G13074);
  or GNAME13077(G13077,G4261,G13019);
  nand GNAME13078(G13078,G13020,G4292);
  nand GNAME13079(G13079,G13078,G13076,G13077);
  or GNAME13080(G13080,G4292,G13020);
  nand GNAME13081(G13081,G13021,G4259);
  nand GNAME13082(G13082,G13081,G13079,G13080);
  or GNAME13083(G13083,G4259,G13021);
  nand GNAME13084(G13084,G13022,G4290);
  nand GNAME13085(G13085,G13084,G13082,G13083);
  or GNAME13086(G13086,G4290,G13022);
  nand GNAME13087(G13087,G13023,G4257);
  nand GNAME13088(G13088,G13087,G13085,G13086);
  or GNAME13089(G13089,G4257,G13023);
  nand GNAME13090(G13090,G13024,G4288);
  nand GNAME13091(G13091,G13090,G13088,G13089);
  or GNAME13092(G13092,G4288,G13024);
  nand GNAME13093(G13093,G13025,G4255);
  nand GNAME13094(G13094,G13093,G13091,G13092);
  or GNAME13095(G13095,G4255,G13025);
  nand GNAME13096(G13096,G13026,G4286);
  nand GNAME13097(G13097,G13096,G13094,G13095);
  or GNAME13098(G13098,G4286,G13026);
  nand GNAME13099(G13099,G13027,G4253);
  nand GNAME13100(G13100,G13099,G13097,G13098);
  or GNAME13101(G13101,G4253,G13027);
  nand GNAME13102(G13102,G13028,G4284);
  nand GNAME13103(G13103,G13102,G13100,G13101);
  or GNAME13104(G13104,G4284,G13028);
  nand GNAME13105(G13105,G13029,G4251);
  nand GNAME13106(G13106,G13105,G13103,G13104);
  or GNAME13107(G13107,G4251,G13029);
  nand GNAME13108(G13108,G13030,G4282);
  nand GNAME13109(G13109,G13108,G13106,G13107);
  or GNAME13110(G13110,G4282,G13030);
  nand GNAME13111(G13111,G13031,G4249);
  nand GNAME13112(G13112,G13111,G13109,G13110);
  or GNAME13113(G13113,G4249,G13031);
  nand GNAME13114(G13114,G13032,G4280);
  nand GNAME13115(G13115,G13114,G13112,G13113);
  or GNAME13116(G13116,G4280,G13032);
  nand GNAME13117(G13117,G13033,G4247);
  nand GNAME13118(G13118,G13117,G13115,G13116);
  or GNAME13119(G13119,G4247,G13033);
  nand GNAME13120(G13120,G13034,G4278);
  nand GNAME13121(G13121,G13120,G13118,G13119);
  or GNAME13122(G13122,G4278,G13034);
  nand GNAME13123(G13123,G13035,G4245);
  nand GNAME13124(G13124,G13123,G13121,G13122);
  or GNAME13125(G13125,G4245,G13035);
  nand GNAME13126(G13126,G13036,G4276);
  nand GNAME13127(G13127,G13126,G13124,G13125);
  or GNAME13128(G13128,G4276,G13036);
  nand GNAME13129(G13129,G13037,G4243);
  nand GNAME13130(G13130,G13129,G13127,G13128);
  or GNAME13131(G13131,G4243,G13037);
  nand GNAME13132(G13132,G13135,G13136,G13130,G13131);
  nand GNAME13133(G13133,G13134,G13137,G13138);
  or GNAME13134(G13134,G13038,G13039);
  or GNAME13135(G13135,G4274,G13038);
  or GNAME13136(G13136,G4242,G13039);
  or GNAME13137(G13137,G4240,G4242);
  nand GNAME13138(G13138,G13039,G4240);
  and GNAME13139(G13139,G13276,G13277);
  and GNAME13140(G13140,G13272,G13274);
  and GNAME13141(G13141,G13269,G13271);
  and GNAME13142(G13142,G13267,G13268);
  and GNAME13143(G13143,G13262,G13264);
  nand GNAME13144(G13144,G13281,G13316,G13317);
  not GNAME13145(G13145,G4699);
  nand GNAME13146(G13146,G4325,G4699);
  not GNAME13147(G13147,G4324);
  not GNAME13148(G13148,G4708);
  not GNAME13149(G13149,G4323);
  not GNAME13150(G13150,G4711);
  not GNAME13151(G13151,G4322);
  not GNAME13152(G13152,G4723);
  not GNAME13153(G13153,G4318);
  not GNAME13154(G13154,G4726);
  not GNAME13155(G13155,G4317);
  not GNAME13156(G13156,G4316);
  not GNAME13157(G13157,G4729);
  not GNAME13158(G13158,G4314);
  not GNAME13159(G13159,G4738);
  not GNAME13160(G13160,G4313);
  not GNAME13161(G13161,G4741);
  not GNAME13162(G13162,G4312);
  not GNAME13163(G13163,G4309);
  not GNAME13164(G13164,G4750);
  nor GNAME13165(G13165,G13350,G13171);
  not GNAME13166(G13166,G4308);
  not GNAME13167(G13167,G4753);
  and GNAME13168(G13168,G13256,G13257);
  not GNAME13169(G13169,G4307);
  not GNAME13170(G13170,G4756);
  and GNAME13171(G13171,G13250,G13265);
  or GNAME13172(G13172,G13249,G13173);
  and GNAME13173(G13173,G13247,G13248);
  and GNAME13174(G13174,G13240,G13241);
  and GNAME13175(G13175,G13237,G13238);
  or GNAME13176(G13176,G13239,G13175);
  nand GNAME13177(G13177,G13348,G13349);
  nand GNAME13178(G13178,G13285,G13286);
  nand GNAME13179(G13179,G13290,G13291);
  nand GNAME13180(G13180,G13295,G13296);
  nand GNAME13181(G13181,G13297,G13298);
  nand GNAME13182(G13182,G13299,G13300);
  nand GNAME13183(G13183,G13301,G13302);
  nand GNAME13184(G13184,G13306,G13307);
  nand GNAME13185(G13185,G13311,G13312);
  nand GNAME13186(G13186,G13324,G13325);
  nand GNAME13187(G13187,G13329,G13330);
  nand GNAME13188(G13188,G13334,G13335);
  nand GNAME13189(G13189,G13339,G13340);
  nand GNAME13190(G13190,G13344,G13345);
  nand GNAME13191(G13191,G13229,G13230);
  nand GNAME13192(G13192,G13226,G13227);
  nand GNAME13193(G13193,G13231,G13224);
  and GNAME13194(G13194,G13221,G13219);
  and GNAME13195(G13195,G13232,G13217);
  and GNAME13196(G13196,G13213,G13214);
  nand GNAME13197(G13197,G13210,G13211);
  or GNAME13198(G13198,G13208,G13199);
  nor GNAME13199(G13199,G13146,G13147);
  not GNAME13200(G13200,G4306);
  not GNAME13201(G13201,G4697);
  and GNAME13202(G13202,G13252,G13253);
  nand GNAME13203(G13203,G13244,G13245);
  or GNAME13204(G13204,G13242,G13174);
  not GNAME13205(G13205,G13165);
  not GNAME13206(G13206,G13146);
  or GNAME13207(G13207,G13206,G4324);
  and GNAME13208(G13208,G13207,G4705);
  nand GNAME13209(G13209,G13149,G13148);
  nand GNAME13210(G13210,G13198,G13209);
  or GNAME13211(G13211,G13148,G13149);
  nand GNAME13212(G13212,G13151,G13150);
  nand GNAME13213(G13213,G13197,G13212);
  or GNAME13214(G13214,G13150,G13151);
  not GNAME13215(G13215,G13196);
  or GNAME13216(G13216,G4714,G4321);
  nand GNAME13217(G13217,G13215,G13216);
  not GNAME13218(G13218,G13195);
  nand GNAME13219(G13219,G4717,G4320);
  or GNAME13220(G13220,G4320,G4717);
  nand GNAME13221(G13221,G13218,G13220);
  not GNAME13222(G13222,G13194);
  or GNAME13223(G13223,G4319,G4720);
  nand GNAME13224(G13224,G13222,G13223);
  nand GNAME13225(G13225,G13153,G13152);
  nand GNAME13226(G13226,G13193,G13225);
  or GNAME13227(G13227,G13152,G13153);
  nand GNAME13228(G13228,G13155,G13154);
  nand GNAME13229(G13229,G13192,G13228);
  or GNAME13230(G13230,G13154,G13155);
  nand GNAME13231(G13231,G4720,G4319);
  nand GNAME13232(G13232,G4321,G4714);
  nand GNAME13233(G13233,G4747,G4310);
  and GNAME13234(G13234,G4744,G4311);
  and GNAME13235(G13235,G4732,G4315);
  nand GNAME13236(G13236,G13156,G13157);
  nand GNAME13237(G13237,G13191,G13236);
  or GNAME13238(G13238,G13156,G13157);
  nor GNAME13239(G13239,G4315,G4732);
  nand GNAME13240(G13240,G13352,G13176);
  or GNAME13241(G13241,G4735,G4314);
  and GNAME13242(G13242,G4735,G4314);
  nand GNAME13243(G13243,G13160,G13159);
  nand GNAME13244(G13244,G13204,G13243);
  or GNAME13245(G13245,G13159,G13160);
  nand GNAME13246(G13246,G13162,G13161);
  nand GNAME13247(G13247,G13203,G13246);
  or GNAME13248(G13248,G13161,G13162);
  nor GNAME13249(G13249,G4311,G4744);
  nand GNAME13250(G13250,G13351,G13172);
  or GNAME13251(G13251,G13163,G13164);
  nand GNAME13252(G13252,G13251,G13165);
  nand GNAME13253(G13253,G13163,G13164);
  not GNAME13254(G13254,G13202);
  or GNAME13255(G13255,G13166,G13167);
  nand GNAME13256(G13256,G13254,G13255);
  nand GNAME13257(G13257,G13166,G13167);
  not GNAME13258(G13258,G13168);
  nand GNAME13259(G13259,G13170,G13169);
  nand GNAME13260(G13260,G13259,G13168);
  or GNAME13261(G13261,G13169,G13170);
  nand GNAME13262(G13262,G13318,G13319,G13260,G13261);
  nand GNAME13263(G13263,G13258,G13261);
  nand GNAME13264(G13264,G13320,G13263,G13259);
  or GNAME13265(G13265,G4310,G4747);
  nand GNAME13266(G13266,G13233,G13265);
  nand GNAME13267(G13267,G13266,G13351,G13172);
  nand GNAME13268(G13268,G13233,G13171);
  or GNAME13269(G13269,G13234,G13172);
  or GNAME13270(G13270,G13234,G13249);
  nand GNAME13271(G13271,G13270,G13173);
  nand GNAME13272(G13272,G13346,G13347,G13352,G13176);
  nand GNAME13273(G13273,G4735,G4314);
  nand GNAME13274(G13274,G13273,G13174);
  or GNAME13275(G13275,G13235,G13239);
  nand GNAME13276(G13276,G13275,G13175);
  or GNAME13277(G13277,G13235,G13176);
  nand GNAME13278(G13278,G13223,G13231);
  nand GNAME13279(G13279,G13219,G13220);
  nand GNAME13280(G13280,G13216,G13232);
  nand GNAME13281(G13281,G13147,G13315);
  or GNAME13282(G13282,G4729,G13156);
  or GNAME13283(G13283,G4316,G13157);
  and GNAME13284(G13284,G13282,G13283);
  nand GNAME13285(G13285,G13191,G13282,G13283);
  or GNAME13286(G13286,G13284,G13191);
  or GNAME13287(G13287,G4726,G13155);
  or GNAME13288(G13288,G4317,G13154);
  and GNAME13289(G13289,G13287,G13288);
  nand GNAME13290(G13290,G13192,G13287,G13288);
  or GNAME13291(G13291,G13289,G13192);
  or GNAME13292(G13292,G4723,G13153);
  or GNAME13293(G13293,G4318,G13152);
  and GNAME13294(G13294,G13292,G13293);
  nand GNAME13295(G13295,G13193,G13292,G13293);
  or GNAME13296(G13296,G13294,G13193);
  nand GNAME13297(G13297,G13222,G13278);
  nand GNAME13298(G13298,G13194,G13223,G13231);
  nand GNAME13299(G13299,G13218,G13279);
  nand GNAME13300(G13300,G13195,G13219,G13220);
  nand GNAME13301(G13301,G13215,G13280);
  nand GNAME13302(G13302,G13196,G13216,G13232);
  or GNAME13303(G13303,G4711,G13151);
  or GNAME13304(G13304,G4322,G13150);
  and GNAME13305(G13305,G13303,G13304);
  nand GNAME13306(G13306,G13197,G13303,G13304);
  or GNAME13307(G13307,G13305,G13197);
  or GNAME13308(G13308,G4708,G13149);
  or GNAME13309(G13309,G4323,G13148);
  and GNAME13310(G13310,G13308,G13309);
  nand GNAME13311(G13311,G13198,G13308,G13309);
  or GNAME13312(G13312,G13310,G13198);
  nand GNAME13313(G13313,G13146,G4705);
  or GNAME13314(G13314,G4705,G13146);
  nand GNAME13315(G13315,G13313,G13314);
  or GNAME13316(G13316,G4705,G13206,G13147);
  nand GNAME13317(G13317,G4705,G13199);
  or GNAME13318(G13318,G4697,G13200);
  or GNAME13319(G13319,G4306,G13201);
  nand GNAME13320(G13320,G13318,G13319);
  or GNAME13321(G13321,G4307,G13170);
  or GNAME13322(G13322,G4756,G13169);
  nand GNAME13323(G13323,G13321,G13322);
  nand GNAME13324(G13324,G13258,G13323);
  nand GNAME13325(G13325,G13168,G13321,G13322);
  or GNAME13326(G13326,G4308,G13167);
  or GNAME13327(G13327,G4753,G13166);
  nand GNAME13328(G13328,G13326,G13327);
  nand GNAME13329(G13329,G13254,G13328);
  nand GNAME13330(G13330,G13202,G13326,G13327);
  or GNAME13331(G13331,G4309,G13164);
  or GNAME13332(G13332,G4750,G13163);
  nand GNAME13333(G13333,G13331,G13332);
  nand GNAME13334(G13334,G13205,G13331,G13332);
  nand GNAME13335(G13335,G13165,G13333);
  or GNAME13336(G13336,G4741,G13162);
  or GNAME13337(G13337,G4312,G13161);
  and GNAME13338(G13338,G13336,G13337);
  nand GNAME13339(G13339,G13203,G13336,G13337);
  or GNAME13340(G13340,G13338,G13203);
  or GNAME13341(G13341,G4738,G13160);
  or GNAME13342(G13342,G4313,G13159);
  and GNAME13343(G13343,G13341,G13342);
  nand GNAME13344(G13344,G13204,G13341,G13342);
  or GNAME13345(G13345,G13343,G13204);
  or GNAME13346(G13346,G4735,G13158);
  nand GNAME13347(G13347,G13158,G4735);
  or GNAME13348(G13348,G4325,G13145);
  nand GNAME13349(G13349,G13145,G4325);
  not GNAME13350(G13350,G13233);
  not GNAME13351(G13351,G13234);
  not GNAME13352(G13352,G13235);
  and GNAME13353(G13353,G13631,G13632);
  and GNAME13354(G13354,G13627,G13629);
  and GNAME13355(G13355,G13623,G13624);
  and GNAME13356(G13356,G13620,G13621);
  and GNAME13357(G13357,G13616,G13618);
  and GNAME13358(G13358,G13613,G13615);
  and GNAME13359(G13359,G13525,G13527);
  and GNAME13360(G13360,G13519,G13520);
  and GNAME13361(G13361,G13515,G13517);
  not GNAME13362(G13362,G4554);
  not GNAME13363(G13363,G4387);
  not GNAME13364(G13364,G4386);
  not GNAME13365(G13365,G4385);
  not GNAME13366(G13366,G4384);
  not GNAME13367(G13367,G4383);
  not GNAME13368(G13368,G4382);
  not GNAME13369(G13369,G4381);
  not GNAME13370(G13370,G4380);
  not GNAME13371(G13371,G4379);
  not GNAME13372(G13372,G4378);
  and GNAME13373(G13373,G13513,G13488);
  or GNAME13374(G13374,G13485,G13373);
  not GNAME13375(G13375,G4358);
  not GNAME13376(G13376,G4377);
  not GNAME13377(G13377,G4376);
  not GNAME13378(G13378,G4375);
  not GNAME13379(G13379,G4374);
  not GNAME13380(G13380,G4373);
  not GNAME13381(G13381,G4372);
  not GNAME13382(G13382,G4371);
  not GNAME13383(G13383,G4370);
  not GNAME13384(G13384,G4369);
  not GNAME13385(G13385,G4368);
  not GNAME13386(G13386,G4367);
  not GNAME13387(G13387,G4366);
  not GNAME13388(G13388,G4365);
  not GNAME13389(G13389,G4364);
  not GNAME13390(G13390,G4363);
  not GNAME13391(G13391,G4362);
  not GNAME13392(G13392,G4361);
  not GNAME13393(G13393,G4360);
  not GNAME13394(G13394,G4359);
  nor GNAME13395(G13395,G13609,G13396);
  and GNAME13396(G13396,G13608,G13607);
  and GNAME13397(G13397,G13523,G13494);
  or GNAME13398(G13398,G13491,G13397);
  and GNAME13399(G13399,G13549,G13548);
  nor GNAME13400(G13400,G13550,G13399);
  and GNAME13401(G13401,G13625,G13510);
  or GNAME13402(G13402,G13534,G13401);
  and GNAME13403(G13403,G13671,G13672);
  and GNAME13404(G13404,G13676,G13677);
  and GNAME13405(G13405,G13681,G13682);
  nand GNAME13406(G13406,G13793,G13794);
  nand GNAME13407(G13407,G13683,G13684);
  nand GNAME13408(G13408,G13685,G13686);
  nand GNAME13409(G13409,G13687,G13688);
  nand GNAME13410(G13410,G13689,G13690);
  nand GNAME13411(G13411,G13757,G13758);
  nand GNAME13412(G13412,G13759,G13760);
  nand GNAME13413(G13413,G13761,G13762);
  nand GNAME13414(G13414,G13763,G13764);
  nand GNAME13415(G13415,G13765,G13766);
  nand GNAME13416(G13416,G13767,G13768);
  nand GNAME13417(G13417,G13769,G13770);
  nand GNAME13418(G13418,G13771,G13772);
  nand GNAME13419(G13419,G13773,G13774);
  nand GNAME13420(G13420,G13775,G13776);
  nand GNAME13421(G13421,G13777,G13778);
  nand GNAME13422(G13422,G13779,G13780);
  nand GNAME13423(G13423,G13781,G13782);
  nand GNAME13424(G13424,G13783,G13784);
  nand GNAME13425(G13425,G13785,G13786);
  nand GNAME13426(G13426,G13787,G13788);
  nand GNAME13427(G13427,G13789,G13790);
  nand GNAME13428(G13428,G13791,G13792);
  not GNAME13429(G13429,G4348);
  not GNAME13430(G13430,G4350);
  not GNAME13431(G13431,G4351);
  not GNAME13432(G13432,G4352);
  not GNAME13433(G13433,G4354);
  not GNAME13434(G13434,G4355);
  not GNAME13435(G13435,G4356);
  nand GNAME13436(G13436,G13505,G13484);
  nand GNAME13437(G13437,G13511,G13482);
  nand GNAME13438(G13438,G13499,G13490);
  not GNAME13439(G13439,G4326);
  not GNAME13440(G13440,G4327);
  not GNAME13441(G13441,G4342);
  not GNAME13442(G13442,G4343);
  not GNAME13443(G13443,G4346);
  not GNAME13444(G13444,G4347);
  not GNAME13445(G13445,G4345);
  not GNAME13446(G13446,G4344);
  not GNAME13447(G13447,G4341);
  not GNAME13448(G13448,G4340);
  not GNAME13449(G13449,G4339);
  not GNAME13450(G13450,G4338);
  not GNAME13451(G13451,G4337);
  not GNAME13452(G13452,G4336);
  not GNAME13453(G13453,G4335);
  not GNAME13454(G13454,G4334);
  not GNAME13455(G13455,G4333);
  not GNAME13456(G13456,G4332);
  not GNAME13457(G13457,G4331);
  not GNAME13458(G13458,G4330);
  not GNAME13459(G13459,G4329);
  not GNAME13460(G13460,G4328);
  nand GNAME13461(G13461,G13604,G13603);
  nand GNAME13462(G13462,G13600,G13599);
  nand GNAME13463(G13463,G13596,G13595);
  nand GNAME13464(G13464,G13592,G13591);
  nand GNAME13465(G13465,G13588,G13587);
  nand GNAME13466(G13466,G13584,G13583);
  nand GNAME13467(G13467,G13580,G13579);
  nand GNAME13468(G13468,G13576,G13575);
  nand GNAME13469(G13469,G13572,G13571);
  nand GNAME13470(G13470,G13568,G13567);
  nand GNAME13471(G13471,G13521,G13481);
  nand GNAME13472(G13472,G13564,G13563);
  nand GNAME13473(G13473,G13560,G13559);
  nand GNAME13474(G13474,G13556,G13555);
  nand GNAME13475(G13475,G13552,G13530);
  or GNAME13476(G13476,G13400,G13531);
  nand GNAME13477(G13477,G13545,G13544);
  nand GNAME13478(G13478,G13541,G13533);
  nand GNAME13479(G13479,G13495,G13481);
  or GNAME13480(G13480,G13405,G13371);
  or GNAME13481(G13481,G13403,G13363);
  or GNAME13482(G13482,G13404,G13367);
  nand GNAME13483(G13483,G13370,G13659,G13660);
  nand GNAME13484(G13484,G13680,G4380);
  and GNAME13485(G13485,G13369,G13661,G13662);
  nand GNAME13486(G13486,G13679,G4381);
  nand GNAME13487(G13487,G13368,G13663,G13664);
  nand GNAME13488(G13488,G13678,G4382);
  nand GNAME13489(G13489,G13366,G13665,G13666);
  nand GNAME13490(G13490,G13675,G4384);
  and GNAME13491(G13491,G13365,G13667,G13668);
  nand GNAME13492(G13492,G13674,G4385);
  nand GNAME13493(G13493,G13364,G13669,G13670);
  nand GNAME13494(G13494,G13673,G4386);
  nand GNAME13495(G13495,G13363,G13403);
  nand GNAME13496(G13496,G13523,G13494);
  nand GNAME13497(G13497,G13796,G13496);
  nand GNAME13498(G13498,G13497,G13492);
  nand GNAME13499(G13499,G13489,G13498);
  not GNAME13500(G13500,G13438);
  nand GNAME13501(G13501,G13367,G13404);
  nand GNAME13502(G13502,G13513,G13488);
  nand GNAME13503(G13503,G13795,G13502);
  nand GNAME13504(G13504,G13503,G13486);
  nand GNAME13505(G13505,G13483,G13504);
  not GNAME13506(G13506,G13436);
  nand GNAME13507(G13507,G13371,G13405);
  not GNAME13508(G13508,G13537);
  nand GNAME13509(G13509,G13372,G13656,G13657);
  nand GNAME13510(G13510,G13658,G4378);
  nand GNAME13511(G13511,G13438,G13501);
  not GNAME13512(G13512,G13437);
  nand GNAME13513(G13513,G13487,G13437);
  nand GNAME13514(G13514,G13486,G13374);
  nand GNAME13515(G13515,G13514,G13483,G13484);
  nand GNAME13516(G13516,G13483,G13484);
  nand GNAME13517(G13517,G13516,G13486,G13374);
  or GNAME13518(G13518,G13485,G13798);
  nand GNAME13519(G13519,G13518,G13373);
  or GNAME13520(G13520,G13798,G13374);
  nand GNAME13521(G13521,G13495,G4554);
  not GNAME13522(G13522,G13471);
  nand GNAME13523(G13523,G13493,G13471);
  nand GNAME13524(G13524,G13492,G13398);
  nand GNAME13525(G13525,G13524,G13489,G13490);
  nand GNAME13526(G13526,G13489,G13490);
  nand GNAME13527(G13527,G13526,G13492,G13398);
  and GNAME13528(G13528,G13694,G4358);
  nand GNAME13529(G13529,G13381,G13697,G13698);
  nand GNAME13530(G13530,G13714,G4372);
  and GNAME13531(G13531,G13713,G4373);
  nand GNAME13532(G13532,G13377,G13701,G13702);
  nand GNAME13533(G13533,G13706,G4376);
  and GNAME13534(G13534,G13376,G13703,G13704);
  nand GNAME13535(G13535,G13705,G4377);
  nand GNAME13536(G13536,G13436,G13507);
  nand GNAME13537(G13537,G13536,G13480);
  nand GNAME13538(G13538,G13625,G13510);
  nand GNAME13539(G13539,G13797,G13538);
  nand GNAME13540(G13540,G13539,G13535);
  nand GNAME13541(G13541,G13532,G13540);
  not GNAME13542(G13542,G13478);
  nand GNAME13543(G13543,G13378,G13707,G13708);
  nand GNAME13544(G13544,G13709,G4375);
  nand GNAME13545(G13545,G13478,G13543);
  not GNAME13546(G13546,G13477);
  nand GNAME13547(G13547,G13379,G13710,G13711);
  nand GNAME13548(G13548,G13712,G4374);
  nand GNAME13549(G13549,G13477,G13547);
  and GNAME13550(G13550,G13380,G13699,G13700);
  not GNAME13551(G13551,G13476);
  nand GNAME13552(G13552,G13529,G13476);
  not GNAME13553(G13553,G13475);
  nand GNAME13554(G13554,G13382,G13715,G13716);
  nand GNAME13555(G13555,G13717,G4371);
  nand GNAME13556(G13556,G13475,G13554);
  not GNAME13557(G13557,G13474);
  nand GNAME13558(G13558,G13383,G13718,G13719);
  nand GNAME13559(G13559,G13720,G4370);
  nand GNAME13560(G13560,G13474,G13558);
  not GNAME13561(G13561,G13473);
  nand GNAME13562(G13562,G13384,G13721,G13722);
  nand GNAME13563(G13563,G13723,G4369);
  nand GNAME13564(G13564,G13473,G13562);
  not GNAME13565(G13565,G13472);
  nand GNAME13566(G13566,G13385,G13724,G13725);
  nand GNAME13567(G13567,G13726,G4368);
  nand GNAME13568(G13568,G13472,G13566);
  not GNAME13569(G13569,G13470);
  nand GNAME13570(G13570,G13386,G13727,G13728);
  nand GNAME13571(G13571,G13729,G4367);
  nand GNAME13572(G13572,G13470,G13570);
  not GNAME13573(G13573,G13469);
  nand GNAME13574(G13574,G13387,G13730,G13731);
  nand GNAME13575(G13575,G13732,G4366);
  nand GNAME13576(G13576,G13469,G13574);
  not GNAME13577(G13577,G13468);
  nand GNAME13578(G13578,G13388,G13733,G13734);
  nand GNAME13579(G13579,G13735,G4365);
  nand GNAME13580(G13580,G13468,G13578);
  not GNAME13581(G13581,G13467);
  nand GNAME13582(G13582,G13389,G13736,G13737);
  nand GNAME13583(G13583,G13738,G4364);
  nand GNAME13584(G13584,G13467,G13582);
  not GNAME13585(G13585,G13466);
  nand GNAME13586(G13586,G13390,G13739,G13740);
  nand GNAME13587(G13587,G13741,G4363);
  nand GNAME13588(G13588,G13466,G13586);
  not GNAME13589(G13589,G13465);
  nand GNAME13590(G13590,G13391,G13742,G13743);
  nand GNAME13591(G13591,G13744,G4362);
  nand GNAME13592(G13592,G13465,G13590);
  not GNAME13593(G13593,G13464);
  nand GNAME13594(G13594,G13392,G13745,G13746);
  nand GNAME13595(G13595,G13747,G4361);
  nand GNAME13596(G13596,G13464,G13594);
  not GNAME13597(G13597,G13463);
  nand GNAME13598(G13598,G13393,G13748,G13749);
  nand GNAME13599(G13599,G13750,G4360);
  nand GNAME13600(G13600,G13463,G13598);
  not GNAME13601(G13601,G13462);
  nand GNAME13602(G13602,G13394,G13751,G13752);
  nand GNAME13603(G13603,G13753,G4359);
  nand GNAME13604(G13604,G13462,G13602);
  not GNAME13605(G13605,G13461);
  nand GNAME13606(G13606,G13375,G13754,G13755);
  nand GNAME13607(G13607,G13756,G4358);
  nand GNAME13608(G13608,G13461,G13606);
  and GNAME13609(G13609,G13375,G13695,G13696);
  or GNAME13610(G13610,G13528,G13395);
  nand GNAME13611(G13611,G13610,G4358);
  or GNAME13612(G13612,G13395,G4358,G13528);
  nand GNAME13613(G13613,G13693,G13611,G13612);
  nand GNAME13614(G13614,G13611,G13612);
  nand GNAME13615(G13615,G13614,G13691,G13692);
  or GNAME13616(G13616,G13528,G13799);
  or GNAME13617(G13617,G13528,G13609);
  nand GNAME13618(G13618,G13617,G13396);
  or GNAME13619(G13619,G13491,G13800);
  nand GNAME13620(G13620,G13619,G13397);
  or GNAME13621(G13621,G13800,G13398);
  or GNAME13622(G13622,G13531,G13550);
  nand GNAME13623(G13623,G13622,G13399);
  or GNAME13624(G13624,G13531,G13801);
  nand GNAME13625(G13625,G13537,G13509);
  nand GNAME13626(G13626,G13535,G13402);
  nand GNAME13627(G13627,G13626,G13532,G13533);
  nand GNAME13628(G13628,G13532,G13533);
  nand GNAME13629(G13629,G13628,G13535,G13402);
  or GNAME13630(G13630,G13534,G13802);
  nand GNAME13631(G13631,G13630,G13401);
  or GNAME13632(G13632,G13802,G13402);
  not GNAME13633(G13633,G13479);
  nand GNAME13634(G13634,G13509,G13510);
  nand GNAME13635(G13635,G13480,G13507);
  nand GNAME13636(G13636,G13487,G13488);
  nand GNAME13637(G13637,G13482,G13501);
  nand GNAME13638(G13638,G13606,G13607);
  nand GNAME13639(G13639,G13602,G13603);
  nand GNAME13640(G13640,G13598,G13599);
  nand GNAME13641(G13641,G13594,G13595);
  nand GNAME13642(G13642,G13590,G13591);
  nand GNAME13643(G13643,G13586,G13587);
  nand GNAME13644(G13644,G13582,G13583);
  nand GNAME13645(G13645,G13578,G13579);
  nand GNAME13646(G13646,G13574,G13575);
  nand GNAME13647(G13647,G13570,G13571);
  nand GNAME13648(G13648,G13493,G13494);
  nand GNAME13649(G13649,G13566,G13567);
  nand GNAME13650(G13650,G13562,G13563);
  nand GNAME13651(G13651,G13558,G13559);
  nand GNAME13652(G13652,G13554,G13555);
  nand GNAME13653(G13653,G13529,G13530);
  nand GNAME13654(G13654,G13547,G13548);
  nand GNAME13655(G13655,G13543,G13544);
  nand GNAME13656(G13656,G13429,G4554);
  nand GNAME13657(G13657,G13362,G4348);
  nand GNAME13658(G13658,G13656,G13657);
  nand GNAME13659(G13659,G13430,G4554);
  nand GNAME13660(G13660,G13362,G4350);
  nand GNAME13661(G13661,G13431,G4554);
  nand GNAME13662(G13662,G13362,G4351);
  nand GNAME13663(G13663,G13432,G4554);
  nand GNAME13664(G13664,G13362,G4352);
  nand GNAME13665(G13665,G13433,G4554);
  nand GNAME13666(G13666,G13362,G4354);
  nand GNAME13667(G13667,G13434,G4554);
  nand GNAME13668(G13668,G13362,G4355);
  nand GNAME13669(G13669,G13435,G4554);
  nand GNAME13670(G13670,G13362,G4356);
  or GNAME13671(G13671,G4357,G13362);
  nand GNAME13672(G13672,G13362,G4357);
  nand GNAME13673(G13673,G13669,G13670);
  nand GNAME13674(G13674,G13667,G13668);
  nand GNAME13675(G13675,G13665,G13666);
  or GNAME13676(G13676,G4353,G13362);
  nand GNAME13677(G13677,G13362,G4353);
  nand GNAME13678(G13678,G13663,G13664);
  nand GNAME13679(G13679,G13661,G13662);
  nand GNAME13680(G13680,G13659,G13660);
  or GNAME13681(G13681,G4349,G13362);
  nand GNAME13682(G13682,G13362,G4349);
  nand GNAME13683(G13683,G13537,G13634);
  nand GNAME13684(G13684,G13508,G13509,G13510);
  nand GNAME13685(G13685,G13436,G13635);
  nand GNAME13686(G13686,G13506,G13480,G13507);
  nand GNAME13687(G13687,G13437,G13636);
  nand GNAME13688(G13688,G13512,G13487,G13488);
  nand GNAME13689(G13689,G13438,G13637);
  nand GNAME13690(G13690,G13500,G13482,G13501);
  nand GNAME13691(G13691,G13439,G4554);
  nand GNAME13692(G13692,G13362,G4326);
  nand GNAME13693(G13693,G13691,G13692);
  nand GNAME13694(G13694,G13695,G13696);
  nand GNAME13695(G13695,G13440,G4554);
  nand GNAME13696(G13696,G13362,G4327);
  nand GNAME13697(G13697,G13441,G4554);
  nand GNAME13698(G13698,G13362,G4342);
  nand GNAME13699(G13699,G13442,G4554);
  nand GNAME13700(G13700,G13362,G4343);
  nand GNAME13701(G13701,G13443,G4554);
  nand GNAME13702(G13702,G13362,G4346);
  nand GNAME13703(G13703,G13444,G4554);
  nand GNAME13704(G13704,G13362,G4347);
  nand GNAME13705(G13705,G13703,G13704);
  nand GNAME13706(G13706,G13701,G13702);
  nand GNAME13707(G13707,G13445,G4554);
  nand GNAME13708(G13708,G13362,G4345);
  nand GNAME13709(G13709,G13707,G13708);
  nand GNAME13710(G13710,G13446,G4554);
  nand GNAME13711(G13711,G13362,G4344);
  nand GNAME13712(G13712,G13710,G13711);
  nand GNAME13713(G13713,G13699,G13700);
  nand GNAME13714(G13714,G13697,G13698);
  nand GNAME13715(G13715,G13447,G4554);
  nand GNAME13716(G13716,G13362,G4341);
  nand GNAME13717(G13717,G13715,G13716);
  nand GNAME13718(G13718,G13448,G4554);
  nand GNAME13719(G13719,G13362,G4340);
  nand GNAME13720(G13720,G13718,G13719);
  nand GNAME13721(G13721,G13449,G4554);
  nand GNAME13722(G13722,G13362,G4339);
  nand GNAME13723(G13723,G13721,G13722);
  nand GNAME13724(G13724,G13450,G4554);
  nand GNAME13725(G13725,G13362,G4338);
  nand GNAME13726(G13726,G13724,G13725);
  nand GNAME13727(G13727,G13451,G4554);
  nand GNAME13728(G13728,G13362,G4337);
  nand GNAME13729(G13729,G13727,G13728);
  nand GNAME13730(G13730,G13452,G4554);
  nand GNAME13731(G13731,G13362,G4336);
  nand GNAME13732(G13732,G13730,G13731);
  nand GNAME13733(G13733,G13453,G4554);
  nand GNAME13734(G13734,G13362,G4335);
  nand GNAME13735(G13735,G13733,G13734);
  nand GNAME13736(G13736,G13454,G4554);
  nand GNAME13737(G13737,G13362,G4334);
  nand GNAME13738(G13738,G13736,G13737);
  nand GNAME13739(G13739,G13455,G4554);
  nand GNAME13740(G13740,G13362,G4333);
  nand GNAME13741(G13741,G13739,G13740);
  nand GNAME13742(G13742,G13456,G4554);
  nand GNAME13743(G13743,G13362,G4332);
  nand GNAME13744(G13744,G13742,G13743);
  nand GNAME13745(G13745,G13457,G4554);
  nand GNAME13746(G13746,G13362,G4331);
  nand GNAME13747(G13747,G13745,G13746);
  nand GNAME13748(G13748,G13458,G4554);
  nand GNAME13749(G13749,G13362,G4330);
  nand GNAME13750(G13750,G13748,G13749);
  nand GNAME13751(G13751,G13459,G4554);
  nand GNAME13752(G13752,G13362,G4329);
  nand GNAME13753(G13753,G13751,G13752);
  nand GNAME13754(G13754,G13460,G4554);
  nand GNAME13755(G13755,G13362,G4328);
  nand GNAME13756(G13756,G13754,G13755);
  nand GNAME13757(G13757,G13461,G13638);
  nand GNAME13758(G13758,G13605,G13606,G13607);
  nand GNAME13759(G13759,G13462,G13639);
  nand GNAME13760(G13760,G13601,G13602,G13603);
  nand GNAME13761(G13761,G13463,G13640);
  nand GNAME13762(G13762,G13597,G13598,G13599);
  nand GNAME13763(G13763,G13464,G13641);
  nand GNAME13764(G13764,G13593,G13594,G13595);
  nand GNAME13765(G13765,G13465,G13642);
  nand GNAME13766(G13766,G13589,G13590,G13591);
  nand GNAME13767(G13767,G13466,G13643);
  nand GNAME13768(G13768,G13585,G13586,G13587);
  nand GNAME13769(G13769,G13467,G13644);
  nand GNAME13770(G13770,G13581,G13582,G13583);
  nand GNAME13771(G13771,G13468,G13645);
  nand GNAME13772(G13772,G13577,G13578,G13579);
  nand GNAME13773(G13773,G13469,G13646);
  nand GNAME13774(G13774,G13573,G13574,G13575);
  nand GNAME13775(G13775,G13470,G13647);
  nand GNAME13776(G13776,G13569,G13570,G13571);
  nand GNAME13777(G13777,G13471,G13648);
  nand GNAME13778(G13778,G13522,G13493,G13494);
  nand GNAME13779(G13779,G13472,G13649);
  nand GNAME13780(G13780,G13565,G13566,G13567);
  nand GNAME13781(G13781,G13473,G13650);
  nand GNAME13782(G13782,G13561,G13562,G13563);
  nand GNAME13783(G13783,G13474,G13651);
  nand GNAME13784(G13784,G13557,G13558,G13559);
  nand GNAME13785(G13785,G13475,G13652);
  nand GNAME13786(G13786,G13553,G13554,G13555);
  nand GNAME13787(G13787,G13476,G13653);
  nand GNAME13788(G13788,G13551,G13529,G13530);
  nand GNAME13789(G13789,G13477,G13654);
  nand GNAME13790(G13790,G13546,G13547,G13548);
  nand GNAME13791(G13791,G13478,G13655);
  nand GNAME13792(G13792,G13542,G13543,G13544);
  nand GNAME13793(G13793,G13479,G4554);
  nand GNAME13794(G13794,G13362,G13633);
  not GNAME13795(G13795,G13485);
  not GNAME13796(G13796,G13491);
  not GNAME13797(G13797,G13534);
  not GNAME13798(G13798,G13486);
  not GNAME13799(G13799,G13395);
  not GNAME13800(G13800,G13492);
  not GNAME13801(G13801,G13400);
  not GNAME13802(G13802,G13535);
  and GNAME13803(G13803,G13822,G13867);
  and GNAME13804(G13804,G13823,G13865);
  and GNAME13805(G13805,G13824,G13864);
  and GNAME13806(G13806,G13825,G13863);
  and GNAME13807(G13807,G13826,G13862);
  and GNAME13808(G13808,G13827,G13861);
  and GNAME13809(G13809,G13828,G13860);
  and GNAME13810(G13810,G13829,G13859);
  and GNAME13811(G13811,G13830,G13858);
  and GNAME13812(G13812,G13831,G13857);
  and GNAME13813(G13813,G13832,G13856);
  and GNAME13814(G13814,G13818,G13855);
  and GNAME13815(G13815,G13819,G13853);
  and GNAME13816(G13816,G13820,G13852);
  and GNAME13817(G13817,G13821,G13851);
  or GNAME13818(G13818,G36219,G36220,G36218);
  or GNAME13819(G13819,G36221,G13818);
  or GNAME13820(G13820,G13874,G36223,G36224);
  or GNAME13821(G13821,G36225,G13820);
  or GNAME13822(G13822,G13870,G36228,G36227);
  or GNAME13823(G13823,G36229,G13822);
  or GNAME13824(G13824,G13898,G36231,G36232);
  or GNAME13825(G13825,G36233,G13824);
  or GNAME13826(G13826,G13894,G36235,G36236);
  or GNAME13827(G13827,G36237,G13826);
  or GNAME13828(G13828,G13888,G36239,G36240);
  or GNAME13829(G13829,G36241,G13828);
  or GNAME13830(G13830,G13884,G36243,G36244);
  or GNAME13831(G13831,G36245,G13830);
  or GNAME13832(G13832,G13831,G36246,G36247);
  nand GNAME13833(G13833,G13889,G13890);
  nand GNAME13834(G13834,G13875,G13876);
  and GNAME13835(G13835,G13866,G13868);
  and GNAME13836(G13836,G13869,G13870);
  and GNAME13837(G13837,G13871,G13872);
  and GNAME13838(G13838,G13873,G13874);
  not GNAME13839(G13839,G36249);
  and GNAME13840(G13840,G13877,G13878);
  and GNAME13841(G13841,G13879,G13880);
  and GNAME13842(G13842,G13881,G13882);
  and GNAME13843(G13843,G13883,G13884);
  and GNAME13844(G13844,G13885,G13886);
  and GNAME13845(G13845,G13887,G13888);
  not GNAME13846(G13846,G36218);
  and GNAME13847(G13847,G13891,G13892);
  and GNAME13848(G13848,G13893,G13894);
  and GNAME13849(G13849,G13895,G13896);
  and GNAME13850(G13850,G13897,G13898);
  nand GNAME13851(G13851,G13820,G36225);
  nand GNAME13852(G13852,G13872,G36224);
  nand GNAME13853(G13853,G13818,G36221);
  or GNAME13854(G13854,G36219,G36218);
  nand GNAME13855(G13855,G13854,G36220);
  nand GNAME13856(G13856,G13880,G36247);
  nand GNAME13857(G13857,G13830,G36245);
  nand GNAME13858(G13858,G13882,G36244);
  nand GNAME13859(G13859,G13828,G36241);
  nand GNAME13860(G13860,G13886,G36240);
  nand GNAME13861(G13861,G13826,G36237);
  nand GNAME13862(G13862,G13892,G36236);
  nand GNAME13863(G13863,G13824,G36233);
  nand GNAME13864(G13864,G13896,G36232);
  nand GNAME13865(G13865,G13822,G36229);
  or GNAME13866(G13866,G36227,G13870);
  nand GNAME13867(G13867,G13866,G36228);
  nand GNAME13868(G13868,G13870,G36227);
  nand GNAME13869(G13869,G13821,G36226);
  or GNAME13870(G13870,G36226,G13821);
  nand GNAME13871(G13871,G13874,G36223);
  or GNAME13872(G13872,G36223,G13874);
  nand GNAME13873(G13873,G13819,G36222);
  or GNAME13874(G13874,G36222,G13819);
  nand GNAME13875(G13875,G13839,G13878);
  or GNAME13876(G13876,G13839,G36248,G13832);
  nand GNAME13877(G13877,G13832,G36248);
  or GNAME13878(G13878,G36248,G13832);
  nand GNAME13879(G13879,G13831,G36246);
  or GNAME13880(G13880,G36246,G13831);
  nand GNAME13881(G13881,G13884,G36243);
  or GNAME13882(G13882,G36243,G13884);
  nand GNAME13883(G13883,G13829,G36242);
  or GNAME13884(G13884,G36242,G13829);
  nand GNAME13885(G13885,G13888,G36239);
  or GNAME13886(G13886,G36239,G13888);
  nand GNAME13887(G13887,G13827,G36238);
  or GNAME13888(G13888,G36238,G13827);
  or GNAME13889(G13889,G36219,G13846);
  nand GNAME13890(G13890,G13846,G36219);
  nand GNAME13891(G13891,G13894,G36235);
  or GNAME13892(G13892,G36235,G13894);
  nand GNAME13893(G13893,G13825,G36234);
  or GNAME13894(G13894,G36234,G13825);
  nand GNAME13895(G13895,G13898,G36231);
  or GNAME13896(G13896,G36231,G13898);
  nand GNAME13897(G13897,G13823,G36230);
  or GNAME13898(G13898,G36230,G13823);
  and GNAME13899(G13899,G13900,G4209);
  not GNAME13900(G13900,G4207);
  not GNAME13901(G13901,G36454);
  and GNAME13902(G13902,G36452,G13937,G36458);
  not GNAME13903(G13903,G36445);
  not GNAME13904(G13904,G36442);
  not GNAME13905(G13905,G36459);
  nor GNAME13906(G13906,G13904,G13901,G13903);
  not GNAME13907(G13907,G36433);
  and GNAME13908(G13908,G36433,G36459,G13906);
  not GNAME13909(G13909,G36451);
  nand GNAME13910(G13910,G13908,G36451);
  and GNAME13911(G13911,G36441,G14026);
  not GNAME13912(G13912,G36436);
  not GNAME13913(G13913,G36455);
  not GNAME13914(G13914,G36438);
  and GNAME13915(G13915,G36455,G13911,G36436);
  not GNAME13916(G13916,G36448);
  not GNAME13917(G13917,G36431);
  and GNAME13918(G13918,G36448,G36438,G13915);
  not GNAME13919(G13919,G36457);
  not GNAME13920(G13920,G36444);
  and GNAME13921(G13921,G36457,G36431,G13918);
  not GNAME13922(G13922,G36446);
  not GNAME13923(G13923,G36453);
  and GNAME13924(G13924,G36446,G36444,G13921);
  not GNAME13925(G13925,G36434);
  not GNAME13926(G13926,G36449);
  and GNAME13927(G13927,G36434,G36453,G13924);
  not GNAME13928(G13928,G36439);
  not GNAME13929(G13929,G36456);
  and GNAME13930(G13930,G36439,G36449,G13927);
  not GNAME13931(G13931,G36437);
  not GNAME13932(G13932,G36447);
  and GNAME13933(G13933,G36437,G36456,G13930);
  not GNAME13934(G13934,G36443);
  and GNAME13935(G13935,G36443,G36447,G13933);
  not GNAME13936(G13936,G36432);
  and GNAME13937(G13937,G13935,G36432);
  not GNAME13938(G13938,G36458);
  not GNAME13939(G13939,G36452);
  nand GNAME13940(G13940,G13976,G13977);
  nand GNAME13941(G13941,G13978,G13979);
  nand GNAME13942(G13942,G13980,G13981);
  nand GNAME13943(G13943,G13982,G13983);
  nand GNAME13944(G13944,G13984,G13985);
  nand GNAME13945(G13945,G13986,G13987);
  nand GNAME13946(G13946,G13988,G13989);
  nand GNAME13947(G13947,G13990,G13991);
  nand GNAME13948(G13948,G13992,G13993);
  nand GNAME13949(G13949,G13994,G13995);
  nand GNAME13950(G13950,G13996,G13997);
  nand GNAME13951(G13951,G13998,G13999);
  nand GNAME13952(G13952,G14000,G14001);
  nand GNAME13953(G13953,G14002,G14003);
  nand GNAME13954(G13954,G14004,G14005);
  nand GNAME13955(G13955,G14006,G14007);
  nand GNAME13956(G13956,G14008,G14009);
  nand GNAME13957(G13957,G14010,G14011);
  nand GNAME13958(G13958,G14012,G14013);
  nand GNAME13959(G13959,G14014,G14015);
  nand GNAME13960(G13960,G14016,G14017);
  nand GNAME13961(G13961,G14018,G14019);
  nand GNAME13962(G13962,G14020,G14021);
  nand GNAME13963(G13963,G14022,G14023);
  nand GNAME13964(G13964,G14024,G14025);
  and GNAME13965(G13965,G13906,G36433);
  nor GNAME13966(G13966,G13901,G13904);
  and GNAME13967(G13967,G13937,G36458);
  and GNAME13968(G13968,G13933,G36443);
  and GNAME13969(G13969,G13930,G36437);
  and GNAME13970(G13970,G13927,G36439);
  and GNAME13971(G13971,G13924,G36434);
  and GNAME13972(G13972,G13921,G36446);
  and GNAME13973(G13973,G13918,G36457);
  and GNAME13974(G13974,G13915,G36448);
  and GNAME13975(G13975,G13911,G36455);
  nand GNAME13976(G13976,G13910,G36441);
  or GNAME13977(G13977,G36441,G13910);
  or GNAME13978(G13978,G13908,G13909);
  nand GNAME13979(G13979,G13909,G13908);
  or GNAME13980(G13980,G13965,G13905);
  nand GNAME13981(G13981,G13905,G13965);
  or GNAME13982(G13982,G13906,G13907);
  nand GNAME13983(G13983,G13907,G13906);
  or GNAME13984(G13984,G13966,G13903);
  nand GNAME13985(G13985,G13903,G13966);
  or GNAME13986(G13986,G36454,G13904);
  or GNAME13987(G13987,G36442,G13901);
  or GNAME13988(G13988,G13967,G13939);
  nand GNAME13989(G13989,G13939,G13967);
  or GNAME13990(G13990,G13937,G13938);
  nand GNAME13991(G13991,G13938,G13937);
  or GNAME13992(G13992,G13935,G13936);
  nand GNAME13993(G13993,G13936,G13935);
  or GNAME13994(G13994,G13968,G13932);
  nand GNAME13995(G13995,G13932,G13968);
  or GNAME13996(G13996,G13933,G13934);
  nand GNAME13997(G13997,G13934,G13933);
  or GNAME13998(G13998,G13969,G13929);
  nand GNAME13999(G13999,G13929,G13969);
  or GNAME14000(G14000,G13930,G13931);
  nand GNAME14001(G14001,G13931,G13930);
  or GNAME14002(G14002,G13970,G13926);
  nand GNAME14003(G14003,G13926,G13970);
  or GNAME14004(G14004,G13927,G13928);
  nand GNAME14005(G14005,G13928,G13927);
  or GNAME14006(G14006,G13971,G13923);
  nand GNAME14007(G14007,G13923,G13971);
  or GNAME14008(G14008,G13924,G13925);
  nand GNAME14009(G14009,G13925,G13924);
  or GNAME14010(G14010,G13972,G13920);
  nand GNAME14011(G14011,G13920,G13972);
  or GNAME14012(G14012,G13921,G13922);
  nand GNAME14013(G14013,G13922,G13921);
  or GNAME14014(G14014,G13973,G13917);
  nand GNAME14015(G14015,G13917,G13973);
  or GNAME14016(G14016,G13918,G13919);
  nand GNAME14017(G14017,G13919,G13918);
  or GNAME14018(G14018,G13974,G13914);
  nand GNAME14019(G14019,G13914,G13974);
  or GNAME14020(G14020,G13915,G13916);
  nand GNAME14021(G14021,G13916,G13915);
  or GNAME14022(G14022,G13975,G13912);
  nand GNAME14023(G14023,G13912,G13975);
  or GNAME14024(G14024,G13911,G13913);
  nand GNAME14025(G14025,G13913,G13911);
  not GNAME14026(G14026,G13910);
  nand GNAME14027(G14027,G14163,G14161);
  nand GNAME14028(G14028,G14164,G14122);
  not GNAME14029(G14029,G7154);
  nor GNAME14030(G14030,G7669,G14029);
  not GNAME14031(G14031,G7153);
  not GNAME14032(G14032,G7672);
  not GNAME14033(G14033,G7152);
  not GNAME14034(G14034,G7673);
  not GNAME14035(G14035,G7151);
  not GNAME14036(G14036,G7674);
  not GNAME14037(G14037,G7150);
  not GNAME14038(G14038,G7675);
  not GNAME14039(G14039,G7149);
  not GNAME14040(G14040,G7676);
  not GNAME14041(G14041,G7148);
  not GNAME14042(G14042,G7677);
  not GNAME14043(G14043,G7147);
  not GNAME14044(G14044,G7678);
  not GNAME14045(G14045,G7146);
  not GNAME14046(G14046,G7679);
  not GNAME14047(G14047,G7145);
  not GNAME14048(G14048,G7680);
  not GNAME14049(G14049,G7144);
  not GNAME14050(G14050,G7681);
  not GNAME14051(G14051,G7143);
  not GNAME14052(G14052,G7682);
  not GNAME14053(G14053,G7142);
  not GNAME14054(G14054,G7683);
  not GNAME14055(G14055,G7141);
  not GNAME14056(G14056,G7684);
  not GNAME14057(G14057,G7140);
  not GNAME14058(G14058,G7685);
  not GNAME14059(G14059,G7139);
  not GNAME14060(G14060,G7686);
  not GNAME14061(G14061,G7138);
  not GNAME14062(G14062,G7687);
  not GNAME14063(G14063,G7137);
  not GNAME14064(G14064,G7136);
  and GNAME14065(G14065,G14158,G14208);
  not GNAME14066(G14066,G7688);
  nand GNAME14067(G14067,G14198,G14199);
  and GNAME14068(G14068,G14165,G14142);
  and GNAME14069(G14069,G14168,G14169);
  and GNAME14070(G14070,G14172,G14173);
  and GNAME14071(G14071,G14176,G14177);
  and GNAME14072(G14072,G14180,G14181);
  and GNAME14073(G14073,G14184,G14185);
  and GNAME14074(G14074,G14188,G14189);
  and GNAME14075(G14075,G14192,G14193);
  and GNAME14076(G14076,G14196,G14197);
  and GNAME14077(G14077,G14203,G14204);
  and GNAME14078(G14078,G14207,G14208);
  and GNAME14079(G14079,G14211,G14212);
  and GNAME14080(G14080,G14215,G14216);
  and GNAME14081(G14081,G14219,G14220);
  and GNAME14082(G14082,G14223,G14224);
  and GNAME14083(G14083,G14227,G14228);
  and GNAME14084(G14084,G14231,G14232);
  and GNAME14085(G14085,G14235,G14236);
  and GNAME14086(G14086,G14139,G14169);
  and GNAME14087(G14087,G14166,G14167);
  and GNAME14088(G14088,G14137,G14173);
  and GNAME14089(G14089,G14170,G14171);
  and GNAME14090(G14090,G14135,G14177);
  and GNAME14091(G14091,G14174,G14175);
  and GNAME14092(G14092,G14133,G14181);
  and GNAME14093(G14093,G14178,G14179);
  and GNAME14094(G14094,G14131,G14185);
  and GNAME14095(G14095,G14182,G14183);
  and GNAME14096(G14096,G14129,G14189);
  and GNAME14097(G14097,G14186,G14187);
  and GNAME14098(G14098,G14127,G14193);
  and GNAME14099(G14099,G14190,G14191);
  and GNAME14100(G14100,G14124,G14125);
  and GNAME14101(G14101,G14194,G14195);
  not GNAME14102(G14102,G7671);
  not GNAME14103(G14103,G7665);
  not GNAME14104(G14104,G7135);
  and GNAME14105(G14105,G14205,G14206);
  and GNAME14106(G14106,G14156,G14212);
  and GNAME14107(G14107,G14209,G14210);
  and GNAME14108(G14108,G14154,G14216);
  and GNAME14109(G14109,G14213,G14214);
  and GNAME14110(G14110,G14152,G14220);
  and GNAME14111(G14111,G14217,G14218);
  and GNAME14112(G14112,G14150,G14224);
  and GNAME14113(G14113,G14221,G14222);
  and GNAME14114(G14114,G14148,G14228);
  and GNAME14115(G14115,G14225,G14226);
  and GNAME14116(G14116,G14146,G14232);
  and GNAME14117(G14117,G14229,G14230);
  and GNAME14118(G14118,G14144,G14236);
  and GNAME14119(G14119,G14233,G14234);
  and GNAME14120(G14120,G14141,G14142);
  and GNAME14121(G14121,G14237,G14238);
  not GNAME14122(G14122,G14030);
  or GNAME14123(G14123,G14030,G7153);
  nand GNAME14124(G14124,G14102,G14123);
  or GNAME14125(G14125,G14122,G14031);
  nor GNAME14126(G14126,G7152,G14032);
  or GNAME14127(G14127,G14100,G14126);
  nor GNAME14128(G14128,G7151,G14034);
  or GNAME14129(G14129,G14098,G14128);
  nor GNAME14130(G14130,G7150,G14036);
  or GNAME14131(G14131,G14096,G14130);
  nor GNAME14132(G14132,G7149,G14038);
  or GNAME14133(G14133,G14094,G14132);
  nor GNAME14134(G14134,G7148,G14040);
  or GNAME14135(G14135,G14092,G14134);
  nor GNAME14136(G14136,G7147,G14042);
  or GNAME14137(G14137,G14090,G14136);
  nor GNAME14138(G14138,G7146,G14044);
  or GNAME14139(G14139,G14088,G14138);
  nor GNAME14140(G14140,G7145,G14046);
  or GNAME14141(G14141,G14086,G14140);
  or GNAME14142(G14142,G7679,G14047);
  nor GNAME14143(G14143,G7144,G14048);
  or GNAME14144(G14144,G14120,G14143);
  nor GNAME14145(G14145,G7143,G14050);
  or GNAME14146(G14146,G14118,G14145);
  nor GNAME14147(G14147,G7142,G14052);
  or GNAME14148(G14148,G14116,G14147);
  nor GNAME14149(G14149,G7141,G14054);
  or GNAME14150(G14150,G14114,G14149);
  nor GNAME14151(G14151,G7140,G14056);
  or GNAME14152(G14152,G14112,G14151);
  nor GNAME14153(G14153,G7139,G14058);
  or GNAME14154(G14154,G14110,G14153);
  nor GNAME14155(G14155,G7138,G14060);
  or GNAME14156(G14156,G14108,G14155);
  nor GNAME14157(G14157,G7137,G14062);
  or GNAME14158(G14158,G14106,G14157);
  nor GNAME14159(G14159,G7136,G14066);
  or GNAME14160(G14160,G14065,G14159);
  nand GNAME14161(G14161,G14202,G14160,G14204);
  nand GNAME14162(G14162,G14204,G14065);
  nand GNAME14163(G14163,G14200,G14201,G14162,G14203);
  nand GNAME14164(G14164,G14029,G7669);
  or GNAME14165(G14165,G7145,G14046);
  nand GNAME14166(G14166,G14068,G14086);
  or GNAME14167(G14167,G14086,G14068);
  or GNAME14168(G14168,G7146,G14044);
  or GNAME14169(G14169,G7678,G14045);
  nand GNAME14170(G14170,G14069,G14088);
  or GNAME14171(G14171,G14088,G14069);
  or GNAME14172(G14172,G7147,G14042);
  or GNAME14173(G14173,G7677,G14043);
  nand GNAME14174(G14174,G14070,G14090);
  or GNAME14175(G14175,G14090,G14070);
  or GNAME14176(G14176,G7148,G14040);
  or GNAME14177(G14177,G7676,G14041);
  nand GNAME14178(G14178,G14071,G14092);
  or GNAME14179(G14179,G14092,G14071);
  or GNAME14180(G14180,G7149,G14038);
  or GNAME14181(G14181,G7675,G14039);
  nand GNAME14182(G14182,G14072,G14094);
  or GNAME14183(G14183,G14094,G14072);
  or GNAME14184(G14184,G7150,G14036);
  or GNAME14185(G14185,G7674,G14037);
  nand GNAME14186(G14186,G14073,G14096);
  or GNAME14187(G14187,G14096,G14073);
  or GNAME14188(G14188,G7151,G14034);
  or GNAME14189(G14189,G7673,G14035);
  nand GNAME14190(G14190,G14074,G14098);
  or GNAME14191(G14191,G14098,G14074);
  or GNAME14192(G14192,G7152,G14032);
  or GNAME14193(G14193,G7672,G14033);
  nand GNAME14194(G14194,G14075,G14100);
  or GNAME14195(G14195,G14100,G14075);
  or GNAME14196(G14196,G7153,G14102);
  or GNAME14197(G14197,G7671,G14031);
  nand GNAME14198(G14198,G14030,G14076);
  or GNAME14199(G14199,G14030,G14076);
  or GNAME14200(G14200,G7135,G14103);
  or GNAME14201(G14201,G7665,G14104);
  nand GNAME14202(G14202,G14200,G14201);
  or GNAME14203(G14203,G7136,G14066);
  or GNAME14204(G14204,G7688,G14064);
  nand GNAME14205(G14205,G14065,G14077);
  or GNAME14206(G14206,G14065,G14077);
  or GNAME14207(G14207,G7137,G14062);
  or GNAME14208(G14208,G7687,G14063);
  nand GNAME14209(G14209,G14078,G14106);
  or GNAME14210(G14210,G14106,G14078);
  or GNAME14211(G14211,G7138,G14060);
  or GNAME14212(G14212,G7686,G14061);
  nand GNAME14213(G14213,G14079,G14108);
  or GNAME14214(G14214,G14108,G14079);
  or GNAME14215(G14215,G7139,G14058);
  or GNAME14216(G14216,G7685,G14059);
  nand GNAME14217(G14217,G14080,G14110);
  or GNAME14218(G14218,G14110,G14080);
  or GNAME14219(G14219,G7140,G14056);
  or GNAME14220(G14220,G7684,G14057);
  nand GNAME14221(G14221,G14081,G14112);
  or GNAME14222(G14222,G14112,G14081);
  or GNAME14223(G14223,G7141,G14054);
  or GNAME14224(G14224,G7683,G14055);
  nand GNAME14225(G14225,G14082,G14114);
  or GNAME14226(G14226,G14114,G14082);
  or GNAME14227(G14227,G7142,G14052);
  or GNAME14228(G14228,G7682,G14053);
  nand GNAME14229(G14229,G14083,G14116);
  or GNAME14230(G14230,G14116,G14083);
  or GNAME14231(G14231,G7143,G14050);
  or GNAME14232(G14232,G7681,G14051);
  nand GNAME14233(G14233,G14084,G14118);
  or GNAME14234(G14234,G14118,G14084);
  or GNAME14235(G14235,G7144,G14048);
  or GNAME14236(G14236,G7680,G14049);
  nand GNAME14237(G14237,G14085,G14120);
  or GNAME14238(G14238,G14120,G14085);
  nand GNAME14239(G14239,G14362,G14365,G14366);
  not GNAME14240(G14240,G7250);
  not GNAME14241(G14241,G7214);
  not GNAME14242(G14242,G7248);
  not GNAME14243(G14243,G7210);
  not GNAME14244(G14244,G7246);
  not GNAME14245(G14245,G7206);
  not GNAME14246(G14246,G7244);
  not GNAME14247(G14247,G7202);
  not GNAME14248(G14248,G7242);
  not GNAME14249(G14249,G7198);
  not GNAME14250(G14250,G7240);
  not GNAME14251(G14251,G7194);
  not GNAME14252(G14252,G7238);
  not GNAME14253(G14253,G7190);
  not GNAME14254(G14254,G7236);
  not GNAME14255(G14255,G7186);
  not GNAME14256(G14256,G7234);
  not GNAME14257(G14257,G7182);
  not GNAME14258(G14258,G7232);
  not GNAME14259(G14259,G7178);
  not GNAME14260(G14260,G7230);
  not GNAME14261(G14261,G7174);
  not GNAME14262(G14262,G7228);
  not GNAME14263(G14263,G7170);
  not GNAME14264(G14264,G7226);
  not GNAME14265(G14265,G7166);
  not GNAME14266(G14266,G7224);
  not GNAME14267(G14267,G7162);
  not GNAME14268(G14268,G7222);
  not GNAME14269(G14269,G7158);
  not GNAME14270(G14270,G7220);
  not GNAME14271(G14271,G7218);
  nand GNAME14272(G14272,G14240,G7216);
  nand GNAME14273(G14273,G7251,G14271,G14272);
  or GNAME14274(G14274,G7216,G14240);
  nand GNAME14275(G14275,G14241,G7249);
  nand GNAME14276(G14276,G14275,G14273,G14274);
  or GNAME14277(G14277,G7249,G14241);
  nand GNAME14278(G14278,G14242,G7212);
  nand GNAME14279(G14279,G14278,G14276,G14277);
  or GNAME14280(G14280,G7212,G14242);
  nand GNAME14281(G14281,G14243,G7247);
  nand GNAME14282(G14282,G14281,G14279,G14280);
  or GNAME14283(G14283,G7247,G14243);
  nand GNAME14284(G14284,G14244,G7208);
  nand GNAME14285(G14285,G14284,G14282,G14283);
  or GNAME14286(G14286,G7208,G14244);
  nand GNAME14287(G14287,G14245,G7245);
  nand GNAME14288(G14288,G14287,G14285,G14286);
  or GNAME14289(G14289,G7245,G14245);
  nand GNAME14290(G14290,G14246,G7204);
  nand GNAME14291(G14291,G14290,G14288,G14289);
  or GNAME14292(G14292,G7204,G14246);
  nand GNAME14293(G14293,G14247,G7243);
  nand GNAME14294(G14294,G14293,G14291,G14292);
  or GNAME14295(G14295,G7243,G14247);
  nand GNAME14296(G14296,G14248,G7200);
  nand GNAME14297(G14297,G14296,G14294,G14295);
  or GNAME14298(G14298,G7200,G14248);
  nand GNAME14299(G14299,G14249,G7241);
  nand GNAME14300(G14300,G14299,G14297,G14298);
  or GNAME14301(G14301,G7241,G14249);
  nand GNAME14302(G14302,G14250,G7196);
  nand GNAME14303(G14303,G14302,G14300,G14301);
  or GNAME14304(G14304,G7196,G14250);
  nand GNAME14305(G14305,G14251,G7239);
  nand GNAME14306(G14306,G14305,G14303,G14304);
  or GNAME14307(G14307,G7239,G14251);
  nand GNAME14308(G14308,G14252,G7192);
  nand GNAME14309(G14309,G14308,G14306,G14307);
  or GNAME14310(G14310,G7192,G14252);
  nand GNAME14311(G14311,G14253,G7237);
  nand GNAME14312(G14312,G14311,G14309,G14310);
  or GNAME14313(G14313,G7237,G14253);
  nand GNAME14314(G14314,G14254,G7188);
  nand GNAME14315(G14315,G14314,G14312,G14313);
  or GNAME14316(G14316,G7188,G14254);
  nand GNAME14317(G14317,G14255,G7235);
  nand GNAME14318(G14318,G14317,G14315,G14316);
  or GNAME14319(G14319,G7235,G14255);
  nand GNAME14320(G14320,G14256,G7184);
  nand GNAME14321(G14321,G14320,G14318,G14319);
  or GNAME14322(G14322,G7184,G14256);
  nand GNAME14323(G14323,G14257,G7233);
  nand GNAME14324(G14324,G14323,G14321,G14322);
  or GNAME14325(G14325,G7233,G14257);
  nand GNAME14326(G14326,G14258,G7180);
  nand GNAME14327(G14327,G14326,G14324,G14325);
  or GNAME14328(G14328,G7180,G14258);
  nand GNAME14329(G14329,G14259,G7231);
  nand GNAME14330(G14330,G14329,G14327,G14328);
  or GNAME14331(G14331,G7231,G14259);
  nand GNAME14332(G14332,G14260,G7176);
  nand GNAME14333(G14333,G14332,G14330,G14331);
  or GNAME14334(G14334,G7176,G14260);
  nand GNAME14335(G14335,G14261,G7229);
  nand GNAME14336(G14336,G14335,G14333,G14334);
  or GNAME14337(G14337,G7229,G14261);
  nand GNAME14338(G14338,G14262,G7172);
  nand GNAME14339(G14339,G14338,G14336,G14337);
  or GNAME14340(G14340,G7172,G14262);
  nand GNAME14341(G14341,G14263,G7227);
  nand GNAME14342(G14342,G14341,G14339,G14340);
  or GNAME14343(G14343,G7227,G14263);
  nand GNAME14344(G14344,G14264,G7168);
  nand GNAME14345(G14345,G14344,G14342,G14343);
  or GNAME14346(G14346,G7168,G14264);
  nand GNAME14347(G14347,G14265,G7225);
  nand GNAME14348(G14348,G14347,G14345,G14346);
  or GNAME14349(G14349,G7225,G14265);
  nand GNAME14350(G14350,G14266,G7164);
  nand GNAME14351(G14351,G14350,G14348,G14349);
  or GNAME14352(G14352,G7164,G14266);
  nand GNAME14353(G14353,G14267,G7223);
  nand GNAME14354(G14354,G14353,G14351,G14352);
  or GNAME14355(G14355,G7223,G14267);
  nand GNAME14356(G14356,G14268,G7160);
  nand GNAME14357(G14357,G14356,G14354,G14355);
  or GNAME14358(G14358,G7160,G14268);
  nand GNAME14359(G14359,G14269,G7221);
  nand GNAME14360(G14360,G14359,G14357,G14358);
  or GNAME14361(G14361,G7221,G14269);
  nand GNAME14362(G14362,G14363,G14364,G14360,G14361);
  nand GNAME14363(G14363,G14270,G7156);
  or GNAME14364(G14364,G7156,G14270);
  nand GNAME14365(G14365,G14270,G7156,G7155);
  or GNAME14366(G14366,G14270,G7156,G7155);
  and GNAME14367(G14367,G14386,G14431);
  and GNAME14368(G14368,G14387,G14429);
  and GNAME14369(G14369,G14388,G14428);
  and GNAME14370(G14370,G14389,G14427);
  and GNAME14371(G14371,G14390,G14426);
  and GNAME14372(G14372,G14391,G14425);
  and GNAME14373(G14373,G14392,G14424);
  and GNAME14374(G14374,G14393,G14423);
  and GNAME14375(G14375,G14394,G14422);
  and GNAME14376(G14376,G14395,G14421);
  and GNAME14377(G14377,G14396,G14420);
  and GNAME14378(G14378,G14382,G14419);
  and GNAME14379(G14379,G14383,G14417);
  and GNAME14380(G14380,G14384,G14416);
  and GNAME14381(G14381,G14385,G14415);
  or GNAME14382(G14382,G36464,G36465,G36463);
  or GNAME14383(G14383,G36466,G14382);
  or GNAME14384(G14384,G14438,G36468,G36469);
  or GNAME14385(G14385,G36470,G14384);
  or GNAME14386(G14386,G14434,G36473,G36472);
  or GNAME14387(G14387,G36474,G14386);
  or GNAME14388(G14388,G14462,G36476,G36477);
  or GNAME14389(G14389,G36478,G14388);
  or GNAME14390(G14390,G14458,G36480,G36481);
  or GNAME14391(G14391,G36482,G14390);
  or GNAME14392(G14392,G14452,G36484,G36485);
  or GNAME14393(G14393,G36486,G14392);
  or GNAME14394(G14394,G14448,G36488,G36489);
  or GNAME14395(G14395,G36490,G14394);
  or GNAME14396(G14396,G14395,G36491,G36492);
  nand GNAME14397(G14397,G14453,G14454);
  nand GNAME14398(G14398,G14439,G14440);
  and GNAME14399(G14399,G14430,G14432);
  and GNAME14400(G14400,G14433,G14434);
  and GNAME14401(G14401,G14435,G14436);
  and GNAME14402(G14402,G14437,G14438);
  not GNAME14403(G14403,G36494);
  and GNAME14404(G14404,G14441,G14442);
  and GNAME14405(G14405,G14443,G14444);
  and GNAME14406(G14406,G14445,G14446);
  and GNAME14407(G14407,G14447,G14448);
  and GNAME14408(G14408,G14449,G14450);
  and GNAME14409(G14409,G14451,G14452);
  not GNAME14410(G14410,G36463);
  and GNAME14411(G14411,G14455,G14456);
  and GNAME14412(G14412,G14457,G14458);
  and GNAME14413(G14413,G14459,G14460);
  and GNAME14414(G14414,G14461,G14462);
  nand GNAME14415(G14415,G14384,G36470);
  nand GNAME14416(G14416,G14436,G36469);
  nand GNAME14417(G14417,G14382,G36466);
  or GNAME14418(G14418,G36464,G36463);
  nand GNAME14419(G14419,G14418,G36465);
  nand GNAME14420(G14420,G14444,G36492);
  nand GNAME14421(G14421,G14394,G36490);
  nand GNAME14422(G14422,G14446,G36489);
  nand GNAME14423(G14423,G14392,G36486);
  nand GNAME14424(G14424,G14450,G36485);
  nand GNAME14425(G14425,G14390,G36482);
  nand GNAME14426(G14426,G14456,G36481);
  nand GNAME14427(G14427,G14388,G36478);
  nand GNAME14428(G14428,G14460,G36477);
  nand GNAME14429(G14429,G14386,G36474);
  or GNAME14430(G14430,G36472,G14434);
  nand GNAME14431(G14431,G14430,G36473);
  nand GNAME14432(G14432,G14434,G36472);
  nand GNAME14433(G14433,G14385,G36471);
  or GNAME14434(G14434,G36471,G14385);
  nand GNAME14435(G14435,G14438,G36468);
  or GNAME14436(G14436,G36468,G14438);
  nand GNAME14437(G14437,G14383,G36467);
  or GNAME14438(G14438,G36467,G14383);
  nand GNAME14439(G14439,G14403,G14442);
  or GNAME14440(G14440,G14403,G36493,G14396);
  nand GNAME14441(G14441,G14396,G36493);
  or GNAME14442(G14442,G36493,G14396);
  nand GNAME14443(G14443,G14395,G36491);
  or GNAME14444(G14444,G36491,G14395);
  nand GNAME14445(G14445,G14448,G36488);
  or GNAME14446(G14446,G36488,G14448);
  nand GNAME14447(G14447,G14393,G36487);
  or GNAME14448(G14448,G36487,G14393);
  nand GNAME14449(G14449,G14452,G36484);
  or GNAME14450(G14450,G36484,G14452);
  nand GNAME14451(G14451,G14391,G36483);
  or GNAME14452(G14452,G36483,G14391);
  or GNAME14453(G14453,G36464,G14410);
  nand GNAME14454(G14454,G14410,G36464);
  nand GNAME14455(G14455,G14458,G36480);
  or GNAME14456(G14456,G36480,G14458);
  nand GNAME14457(G14457,G14389,G36479);
  or GNAME14458(G14458,G36479,G14389);
  nand GNAME14459(G14459,G14462,G36476);
  or GNAME14460(G14460,G36476,G14462);
  nand GNAME14461(G14461,G14387,G36475);
  or GNAME14462(G14462,G36475,G14387);
  and GNAME14463(G14463,G14741,G14742);
  and GNAME14464(G14464,G14737,G14739);
  and GNAME14465(G14465,G14733,G14734);
  and GNAME14466(G14466,G14730,G14731);
  and GNAME14467(G14467,G14726,G14728);
  and GNAME14468(G14468,G14723,G14725);
  and GNAME14469(G14469,G14635,G14637);
  and GNAME14470(G14470,G14629,G14630);
  and GNAME14471(G14471,G14625,G14627);
  not GNAME14472(G14472,G7252);
  not GNAME14473(G14473,G7315);
  not GNAME14474(G14474,G7314);
  not GNAME14475(G14475,G7313);
  not GNAME14476(G14476,G7312);
  not GNAME14477(G14477,G7311);
  not GNAME14478(G14478,G7310);
  not GNAME14479(G14479,G7309);
  not GNAME14480(G14480,G7308);
  not GNAME14481(G14481,G7307);
  not GNAME14482(G14482,G7306);
  and GNAME14483(G14483,G14623,G14598);
  or GNAME14484(G14484,G14595,G14483);
  not GNAME14485(G14485,G7285);
  not GNAME14486(G14486,G7305);
  not GNAME14487(G14487,G7304);
  not GNAME14488(G14488,G7303);
  not GNAME14489(G14489,G7302);
  not GNAME14490(G14490,G7301);
  not GNAME14491(G14491,G7300);
  not GNAME14492(G14492,G7299);
  not GNAME14493(G14493,G7298);
  not GNAME14494(G14494,G7297);
  not GNAME14495(G14495,G7296);
  not GNAME14496(G14496,G7295);
  not GNAME14497(G14497,G7294);
  not GNAME14498(G14498,G7293);
  not GNAME14499(G14499,G7292);
  not GNAME14500(G14500,G7291);
  not GNAME14501(G14501,G7290);
  not GNAME14502(G14502,G7289);
  not GNAME14503(G14503,G7288);
  not GNAME14504(G14504,G7287);
  not GNAME14505(G14505,G7286);
  nor GNAME14506(G14506,G14719,G14507);
  and GNAME14507(G14507,G14718,G14717);
  and GNAME14508(G14508,G14633,G14604);
  or GNAME14509(G14509,G14601,G14508);
  and GNAME14510(G14510,G14659,G14658);
  nor GNAME14511(G14511,G14660,G14510);
  and GNAME14512(G14512,G14735,G14620);
  or GNAME14513(G14513,G14644,G14512);
  and GNAME14514(G14514,G14781,G14782);
  and GNAME14515(G14515,G14786,G14787);
  and GNAME14516(G14516,G14791,G14792);
  nand GNAME14517(G14517,G14903,G14904);
  nand GNAME14518(G14518,G14793,G14794);
  nand GNAME14519(G14519,G14795,G14796);
  nand GNAME14520(G14520,G14797,G14798);
  nand GNAME14521(G14521,G14799,G14800);
  nand GNAME14522(G14522,G14867,G14868);
  nand GNAME14523(G14523,G14869,G14870);
  nand GNAME14524(G14524,G14871,G14872);
  nand GNAME14525(G14525,G14873,G14874);
  nand GNAME14526(G14526,G14875,G14876);
  nand GNAME14527(G14527,G14877,G14878);
  nand GNAME14528(G14528,G14879,G14880);
  nand GNAME14529(G14529,G14881,G14882);
  nand GNAME14530(G14530,G14883,G14884);
  nand GNAME14531(G14531,G14885,G14886);
  nand GNAME14532(G14532,G14887,G14888);
  nand GNAME14533(G14533,G14889,G14890);
  nand GNAME14534(G14534,G14891,G14892);
  nand GNAME14535(G14535,G14893,G14894);
  nand GNAME14536(G14536,G14895,G14896);
  nand GNAME14537(G14537,G14897,G14898);
  nand GNAME14538(G14538,G14899,G14900);
  nand GNAME14539(G14539,G14901,G14902);
  not GNAME14540(G14540,G7274);
  not GNAME14541(G14541,G7276);
  not GNAME14542(G14542,G7277);
  not GNAME14543(G14543,G7278);
  not GNAME14544(G14544,G7280);
  not GNAME14545(G14545,G7281);
  not GNAME14546(G14546,G7282);
  nand GNAME14547(G14547,G14615,G14594);
  nand GNAME14548(G14548,G14621,G14592);
  nand GNAME14549(G14549,G14609,G14600);
  not GNAME14550(G14550,G7254);
  not GNAME14551(G14551,G7253);
  not GNAME14552(G14552,G7268);
  not GNAME14553(G14553,G7269);
  not GNAME14554(G14554,G7272);
  not GNAME14555(G14555,G7273);
  not GNAME14556(G14556,G7271);
  not GNAME14557(G14557,G7270);
  not GNAME14558(G14558,G7267);
  not GNAME14559(G14559,G7266);
  not GNAME14560(G14560,G7265);
  not GNAME14561(G14561,G7264);
  not GNAME14562(G14562,G7263);
  not GNAME14563(G14563,G7262);
  not GNAME14564(G14564,G7261);
  not GNAME14565(G14565,G7260);
  not GNAME14566(G14566,G7259);
  not GNAME14567(G14567,G7258);
  not GNAME14568(G14568,G7257);
  not GNAME14569(G14569,G7256);
  not GNAME14570(G14570,G7255);
  nand GNAME14571(G14571,G14714,G14713);
  nand GNAME14572(G14572,G14710,G14709);
  nand GNAME14573(G14573,G14706,G14705);
  nand GNAME14574(G14574,G14702,G14701);
  nand GNAME14575(G14575,G14698,G14697);
  nand GNAME14576(G14576,G14694,G14693);
  nand GNAME14577(G14577,G14690,G14689);
  nand GNAME14578(G14578,G14686,G14685);
  nand GNAME14579(G14579,G14682,G14681);
  nand GNAME14580(G14580,G14678,G14677);
  nand GNAME14581(G14581,G14631,G14591);
  nand GNAME14582(G14582,G14674,G14673);
  nand GNAME14583(G14583,G14670,G14669);
  nand GNAME14584(G14584,G14666,G14665);
  nand GNAME14585(G14585,G14662,G14640);
  or GNAME14586(G14586,G14511,G14641);
  nand GNAME14587(G14587,G14655,G14654);
  nand GNAME14588(G14588,G14651,G14643);
  nand GNAME14589(G14589,G14605,G14591);
  or GNAME14590(G14590,G14516,G14481);
  or GNAME14591(G14591,G14514,G14473);
  or GNAME14592(G14592,G14515,G14477);
  nand GNAME14593(G14593,G14480,G14769,G14770);
  nand GNAME14594(G14594,G14790,G7308);
  and GNAME14595(G14595,G14479,G14771,G14772);
  nand GNAME14596(G14596,G14789,G7309);
  nand GNAME14597(G14597,G14478,G14773,G14774);
  nand GNAME14598(G14598,G14788,G7310);
  nand GNAME14599(G14599,G14476,G14775,G14776);
  nand GNAME14600(G14600,G14785,G7312);
  and GNAME14601(G14601,G14475,G14777,G14778);
  nand GNAME14602(G14602,G14784,G7313);
  nand GNAME14603(G14603,G14474,G14779,G14780);
  nand GNAME14604(G14604,G14783,G7314);
  nand GNAME14605(G14605,G14473,G14514);
  nand GNAME14606(G14606,G14633,G14604);
  nand GNAME14607(G14607,G14906,G14606);
  nand GNAME14608(G14608,G14607,G14602);
  nand GNAME14609(G14609,G14599,G14608);
  not GNAME14610(G14610,G14549);
  nand GNAME14611(G14611,G14477,G14515);
  nand GNAME14612(G14612,G14623,G14598);
  nand GNAME14613(G14613,G14905,G14612);
  nand GNAME14614(G14614,G14613,G14596);
  nand GNAME14615(G14615,G14593,G14614);
  not GNAME14616(G14616,G14547);
  nand GNAME14617(G14617,G14481,G14516);
  not GNAME14618(G14618,G14647);
  nand GNAME14619(G14619,G14482,G14766,G14767);
  nand GNAME14620(G14620,G14768,G7306);
  nand GNAME14621(G14621,G14549,G14611);
  not GNAME14622(G14622,G14548);
  nand GNAME14623(G14623,G14597,G14548);
  nand GNAME14624(G14624,G14596,G14484);
  nand GNAME14625(G14625,G14624,G14593,G14594);
  nand GNAME14626(G14626,G14593,G14594);
  nand GNAME14627(G14627,G14626,G14596,G14484);
  or GNAME14628(G14628,G14595,G14908);
  nand GNAME14629(G14629,G14628,G14483);
  or GNAME14630(G14630,G14908,G14484);
  nand GNAME14631(G14631,G14605,G7252);
  not GNAME14632(G14632,G14581);
  nand GNAME14633(G14633,G14603,G14581);
  nand GNAME14634(G14634,G14602,G14509);
  nand GNAME14635(G14635,G14634,G14599,G14600);
  nand GNAME14636(G14636,G14599,G14600);
  nand GNAME14637(G14637,G14636,G14602,G14509);
  and GNAME14638(G14638,G14804,G7285);
  nand GNAME14639(G14639,G14491,G14807,G14808);
  nand GNAME14640(G14640,G14824,G7300);
  and GNAME14641(G14641,G14823,G7301);
  nand GNAME14642(G14642,G14487,G14811,G14812);
  nand GNAME14643(G14643,G14816,G7304);
  and GNAME14644(G14644,G14486,G14813,G14814);
  nand GNAME14645(G14645,G14815,G7305);
  nand GNAME14646(G14646,G14547,G14617);
  nand GNAME14647(G14647,G14646,G14590);
  nand GNAME14648(G14648,G14735,G14620);
  nand GNAME14649(G14649,G14907,G14648);
  nand GNAME14650(G14650,G14649,G14645);
  nand GNAME14651(G14651,G14642,G14650);
  not GNAME14652(G14652,G14588);
  nand GNAME14653(G14653,G14488,G14817,G14818);
  nand GNAME14654(G14654,G14819,G7303);
  nand GNAME14655(G14655,G14588,G14653);
  not GNAME14656(G14656,G14587);
  nand GNAME14657(G14657,G14489,G14820,G14821);
  nand GNAME14658(G14658,G14822,G7302);
  nand GNAME14659(G14659,G14587,G14657);
  and GNAME14660(G14660,G14490,G14809,G14810);
  not GNAME14661(G14661,G14586);
  nand GNAME14662(G14662,G14639,G14586);
  not GNAME14663(G14663,G14585);
  nand GNAME14664(G14664,G14492,G14825,G14826);
  nand GNAME14665(G14665,G14827,G7299);
  nand GNAME14666(G14666,G14585,G14664);
  not GNAME14667(G14667,G14584);
  nand GNAME14668(G14668,G14493,G14828,G14829);
  nand GNAME14669(G14669,G14830,G7298);
  nand GNAME14670(G14670,G14584,G14668);
  not GNAME14671(G14671,G14583);
  nand GNAME14672(G14672,G14494,G14831,G14832);
  nand GNAME14673(G14673,G14833,G7297);
  nand GNAME14674(G14674,G14583,G14672);
  not GNAME14675(G14675,G14582);
  nand GNAME14676(G14676,G14495,G14834,G14835);
  nand GNAME14677(G14677,G14836,G7296);
  nand GNAME14678(G14678,G14582,G14676);
  not GNAME14679(G14679,G14580);
  nand GNAME14680(G14680,G14496,G14837,G14838);
  nand GNAME14681(G14681,G14839,G7295);
  nand GNAME14682(G14682,G14580,G14680);
  not GNAME14683(G14683,G14579);
  nand GNAME14684(G14684,G14497,G14840,G14841);
  nand GNAME14685(G14685,G14842,G7294);
  nand GNAME14686(G14686,G14579,G14684);
  not GNAME14687(G14687,G14578);
  nand GNAME14688(G14688,G14498,G14843,G14844);
  nand GNAME14689(G14689,G14845,G7293);
  nand GNAME14690(G14690,G14578,G14688);
  not GNAME14691(G14691,G14577);
  nand GNAME14692(G14692,G14499,G14846,G14847);
  nand GNAME14693(G14693,G14848,G7292);
  nand GNAME14694(G14694,G14577,G14692);
  not GNAME14695(G14695,G14576);
  nand GNAME14696(G14696,G14500,G14849,G14850);
  nand GNAME14697(G14697,G14851,G7291);
  nand GNAME14698(G14698,G14576,G14696);
  not GNAME14699(G14699,G14575);
  nand GNAME14700(G14700,G14501,G14852,G14853);
  nand GNAME14701(G14701,G14854,G7290);
  nand GNAME14702(G14702,G14575,G14700);
  not GNAME14703(G14703,G14574);
  nand GNAME14704(G14704,G14502,G14855,G14856);
  nand GNAME14705(G14705,G14857,G7289);
  nand GNAME14706(G14706,G14574,G14704);
  not GNAME14707(G14707,G14573);
  nand GNAME14708(G14708,G14503,G14858,G14859);
  nand GNAME14709(G14709,G14860,G7288);
  nand GNAME14710(G14710,G14573,G14708);
  not GNAME14711(G14711,G14572);
  nand GNAME14712(G14712,G14504,G14861,G14862);
  nand GNAME14713(G14713,G14863,G7287);
  nand GNAME14714(G14714,G14572,G14712);
  not GNAME14715(G14715,G14571);
  nand GNAME14716(G14716,G14505,G14864,G14865);
  nand GNAME14717(G14717,G14866,G7286);
  nand GNAME14718(G14718,G14571,G14716);
  and GNAME14719(G14719,G14485,G14805,G14806);
  or GNAME14720(G14720,G14638,G14506);
  nand GNAME14721(G14721,G14720,G7284);
  or GNAME14722(G14722,G14506,G7284,G14638);
  nand GNAME14723(G14723,G14803,G14721,G14722);
  nand GNAME14724(G14724,G14721,G14722);
  nand GNAME14725(G14725,G14724,G14801,G14802);
  or GNAME14726(G14726,G14638,G14909);
  or GNAME14727(G14727,G14638,G14719);
  nand GNAME14728(G14728,G14727,G14507);
  or GNAME14729(G14729,G14601,G14910);
  nand GNAME14730(G14730,G14729,G14508);
  or GNAME14731(G14731,G14910,G14509);
  or GNAME14732(G14732,G14641,G14660);
  nand GNAME14733(G14733,G14732,G14510);
  or GNAME14734(G14734,G14641,G14911);
  nand GNAME14735(G14735,G14647,G14619);
  nand GNAME14736(G14736,G14645,G14513);
  nand GNAME14737(G14737,G14736,G14642,G14643);
  nand GNAME14738(G14738,G14642,G14643);
  nand GNAME14739(G14739,G14738,G14645,G14513);
  or GNAME14740(G14740,G14644,G14912);
  nand GNAME14741(G14741,G14740,G14512);
  or GNAME14742(G14742,G14912,G14513);
  not GNAME14743(G14743,G14589);
  nand GNAME14744(G14744,G14619,G14620);
  nand GNAME14745(G14745,G14590,G14617);
  nand GNAME14746(G14746,G14597,G14598);
  nand GNAME14747(G14747,G14592,G14611);
  nand GNAME14748(G14748,G14716,G14717);
  nand GNAME14749(G14749,G14712,G14713);
  nand GNAME14750(G14750,G14708,G14709);
  nand GNAME14751(G14751,G14704,G14705);
  nand GNAME14752(G14752,G14700,G14701);
  nand GNAME14753(G14753,G14696,G14697);
  nand GNAME14754(G14754,G14692,G14693);
  nand GNAME14755(G14755,G14688,G14689);
  nand GNAME14756(G14756,G14684,G14685);
  nand GNAME14757(G14757,G14680,G14681);
  nand GNAME14758(G14758,G14603,G14604);
  nand GNAME14759(G14759,G14676,G14677);
  nand GNAME14760(G14760,G14672,G14673);
  nand GNAME14761(G14761,G14668,G14669);
  nand GNAME14762(G14762,G14664,G14665);
  nand GNAME14763(G14763,G14639,G14640);
  nand GNAME14764(G14764,G14657,G14658);
  nand GNAME14765(G14765,G14653,G14654);
  nand GNAME14766(G14766,G14540,G7252);
  nand GNAME14767(G14767,G14472,G7274);
  nand GNAME14768(G14768,G14766,G14767);
  nand GNAME14769(G14769,G14541,G7252);
  nand GNAME14770(G14770,G14472,G7276);
  nand GNAME14771(G14771,G14542,G7252);
  nand GNAME14772(G14772,G14472,G7277);
  nand GNAME14773(G14773,G14543,G7252);
  nand GNAME14774(G14774,G14472,G7278);
  nand GNAME14775(G14775,G14544,G7252);
  nand GNAME14776(G14776,G14472,G7280);
  nand GNAME14777(G14777,G14545,G7252);
  nand GNAME14778(G14778,G14472,G7281);
  nand GNAME14779(G14779,G14546,G7252);
  nand GNAME14780(G14780,G14472,G7282);
  or GNAME14781(G14781,G7283,G14472);
  nand GNAME14782(G14782,G14472,G7283);
  nand GNAME14783(G14783,G14779,G14780);
  nand GNAME14784(G14784,G14777,G14778);
  nand GNAME14785(G14785,G14775,G14776);
  or GNAME14786(G14786,G7279,G14472);
  nand GNAME14787(G14787,G14472,G7279);
  nand GNAME14788(G14788,G14773,G14774);
  nand GNAME14789(G14789,G14771,G14772);
  nand GNAME14790(G14790,G14769,G14770);
  or GNAME14791(G14791,G7275,G14472);
  nand GNAME14792(G14792,G14472,G7275);
  nand GNAME14793(G14793,G14647,G14744);
  nand GNAME14794(G14794,G14618,G14619,G14620);
  nand GNAME14795(G14795,G14547,G14745);
  nand GNAME14796(G14796,G14616,G14590,G14617);
  nand GNAME14797(G14797,G14548,G14746);
  nand GNAME14798(G14798,G14622,G14597,G14598);
  nand GNAME14799(G14799,G14549,G14747);
  nand GNAME14800(G14800,G14610,G14592,G14611);
  nand GNAME14801(G14801,G14550,G7252);
  nand GNAME14802(G14802,G14472,G7254);
  nand GNAME14803(G14803,G14801,G14802);
  nand GNAME14804(G14804,G14805,G14806);
  nand GNAME14805(G14805,G14551,G7252);
  nand GNAME14806(G14806,G14472,G7253);
  nand GNAME14807(G14807,G14552,G7252);
  nand GNAME14808(G14808,G14472,G7268);
  nand GNAME14809(G14809,G14553,G7252);
  nand GNAME14810(G14810,G14472,G7269);
  nand GNAME14811(G14811,G14554,G7252);
  nand GNAME14812(G14812,G14472,G7272);
  nand GNAME14813(G14813,G14555,G7252);
  nand GNAME14814(G14814,G14472,G7273);
  nand GNAME14815(G14815,G14813,G14814);
  nand GNAME14816(G14816,G14811,G14812);
  nand GNAME14817(G14817,G14556,G7252);
  nand GNAME14818(G14818,G14472,G7271);
  nand GNAME14819(G14819,G14817,G14818);
  nand GNAME14820(G14820,G14557,G7252);
  nand GNAME14821(G14821,G14472,G7270);
  nand GNAME14822(G14822,G14820,G14821);
  nand GNAME14823(G14823,G14809,G14810);
  nand GNAME14824(G14824,G14807,G14808);
  nand GNAME14825(G14825,G14558,G7252);
  nand GNAME14826(G14826,G14472,G7267);
  nand GNAME14827(G14827,G14825,G14826);
  nand GNAME14828(G14828,G14559,G7252);
  nand GNAME14829(G14829,G14472,G7266);
  nand GNAME14830(G14830,G14828,G14829);
  nand GNAME14831(G14831,G14560,G7252);
  nand GNAME14832(G14832,G14472,G7265);
  nand GNAME14833(G14833,G14831,G14832);
  nand GNAME14834(G14834,G14561,G7252);
  nand GNAME14835(G14835,G14472,G7264);
  nand GNAME14836(G14836,G14834,G14835);
  nand GNAME14837(G14837,G14562,G7252);
  nand GNAME14838(G14838,G14472,G7263);
  nand GNAME14839(G14839,G14837,G14838);
  nand GNAME14840(G14840,G14563,G7252);
  nand GNAME14841(G14841,G14472,G7262);
  nand GNAME14842(G14842,G14840,G14841);
  nand GNAME14843(G14843,G14564,G7252);
  nand GNAME14844(G14844,G14472,G7261);
  nand GNAME14845(G14845,G14843,G14844);
  nand GNAME14846(G14846,G14565,G7252);
  nand GNAME14847(G14847,G14472,G7260);
  nand GNAME14848(G14848,G14846,G14847);
  nand GNAME14849(G14849,G14566,G7252);
  nand GNAME14850(G14850,G14472,G7259);
  nand GNAME14851(G14851,G14849,G14850);
  nand GNAME14852(G14852,G14567,G7252);
  nand GNAME14853(G14853,G14472,G7258);
  nand GNAME14854(G14854,G14852,G14853);
  nand GNAME14855(G14855,G14568,G7252);
  nand GNAME14856(G14856,G14472,G7257);
  nand GNAME14857(G14857,G14855,G14856);
  nand GNAME14858(G14858,G14569,G7252);
  nand GNAME14859(G14859,G14472,G7256);
  nand GNAME14860(G14860,G14858,G14859);
  nand GNAME14861(G14861,G14570,G7252);
  nand GNAME14862(G14862,G14472,G7255);
  nand GNAME14863(G14863,G14861,G14862);
  nand GNAME14864(G14864,G14550,G7252);
  nand GNAME14865(G14865,G14472,G7254);
  nand GNAME14866(G14866,G14864,G14865);
  nand GNAME14867(G14867,G14571,G14748);
  nand GNAME14868(G14868,G14715,G14716,G14717);
  nand GNAME14869(G14869,G14572,G14749);
  nand GNAME14870(G14870,G14711,G14712,G14713);
  nand GNAME14871(G14871,G14573,G14750);
  nand GNAME14872(G14872,G14707,G14708,G14709);
  nand GNAME14873(G14873,G14574,G14751);
  nand GNAME14874(G14874,G14703,G14704,G14705);
  nand GNAME14875(G14875,G14575,G14752);
  nand GNAME14876(G14876,G14699,G14700,G14701);
  nand GNAME14877(G14877,G14576,G14753);
  nand GNAME14878(G14878,G14695,G14696,G14697);
  nand GNAME14879(G14879,G14577,G14754);
  nand GNAME14880(G14880,G14691,G14692,G14693);
  nand GNAME14881(G14881,G14578,G14755);
  nand GNAME14882(G14882,G14687,G14688,G14689);
  nand GNAME14883(G14883,G14579,G14756);
  nand GNAME14884(G14884,G14683,G14684,G14685);
  nand GNAME14885(G14885,G14580,G14757);
  nand GNAME14886(G14886,G14679,G14680,G14681);
  nand GNAME14887(G14887,G14581,G14758);
  nand GNAME14888(G14888,G14632,G14603,G14604);
  nand GNAME14889(G14889,G14582,G14759);
  nand GNAME14890(G14890,G14675,G14676,G14677);
  nand GNAME14891(G14891,G14583,G14760);
  nand GNAME14892(G14892,G14671,G14672,G14673);
  nand GNAME14893(G14893,G14584,G14761);
  nand GNAME14894(G14894,G14667,G14668,G14669);
  nand GNAME14895(G14895,G14585,G14762);
  nand GNAME14896(G14896,G14663,G14664,G14665);
  nand GNAME14897(G14897,G14586,G14763);
  nand GNAME14898(G14898,G14661,G14639,G14640);
  nand GNAME14899(G14899,G14587,G14764);
  nand GNAME14900(G14900,G14656,G14657,G14658);
  nand GNAME14901(G14901,G14588,G14765);
  nand GNAME14902(G14902,G14652,G14653,G14654);
  nand GNAME14903(G14903,G14589,G7252);
  nand GNAME14904(G14904,G14472,G14743);
  not GNAME14905(G14905,G14595);
  not GNAME14906(G14906,G14601);
  not GNAME14907(G14907,G14644);
  not GNAME14908(G14908,G14596);
  not GNAME14909(G14909,G14506);
  not GNAME14910(G14910,G14602);
  not GNAME14911(G14911,G14511);
  not GNAME14912(G14912,G14645);
  not GNAME14913(G14913,G7159);
  and GNAME14914(G14914,G14915,G14916);
  nand GNAME14915(G14915,G14913,G7157);
  or GNAME14916(G14916,G7157,G14913);
  nand GNAME14917(G14917,G14979,G14962);
  nand GNAME14918(G14918,G14986,G14955);
  nand GNAME14919(G14919,G14971,G14945);
  nand GNAME14920(G14920,G14991,G14950);
  nand GNAME14921(G14921,G14978,G14963);
  nand GNAME14922(G14922,G14984,G14957);
  nand GNAME14923(G14923,G14969,G14947);
  nand GNAME14924(G14924,G14992,G14949);
  nand GNAME14925(G14925,G14968,G14948);
  nand GNAME14926(G14926,G14983,G14958);
  nand GNAME14927(G14927,G14977,G14964);
  nand GNAME14928(G14928,G14980,G14961);
  nand GNAME14929(G14929,G14970,G14946);
  nand GNAME14930(G14930,G14985,G14956);
  nand GNAME14931(G14931,G14982,G14959);
  nand GNAME14932(G14932,G14987,G14954);
  nand GNAME14933(G14933,G14972,G14944);
  nand GNAME14934(G14934,G14975,G14966);
  nand GNAME14935(G14935,G14990,G14951);
  nand GNAME14936(G14936,G14989,G14952);
  not GNAME14937(G14937,G36699);
  nand GNAME14938(G14938,G14976,G14965);
  nand GNAME14939(G14939,G14981,G14960);
  or GNAME14940(G14940,G14974,G14967);
  nand GNAME14941(G14941,G14973,G14943);
  nand GNAME14942(G14942,G14988,G14953);
  or GNAME14943(G14943,G36687,G36699);
  or GNAME14944(G14944,G36690,G14943);
  or GNAME14945(G14945,G36678,G14944);
  or GNAME14946(G14946,G36704,G14945);
  or GNAME14947(G14947,G36696,G14946);
  or GNAME14948(G14948,G36686,G14947);
  or GNAME14949(G14949,G36700,G14948);
  or GNAME14950(G14950,G36681,G14949);
  or GNAME14951(G14951,G36693,G14950);
  or GNAME14952(G14952,G36683,G14951);
  or GNAME14953(G14953,G36702,G14952);
  or GNAME14954(G14954,G36676,G14953);
  or GNAME14955(G14955,G36691,G14954);
  or GNAME14956(G14956,G36689,G14955);
  or GNAME14957(G14957,G36679,G14956);
  or GNAME14958(G14958,G36698,G14957);
  or GNAME14959(G14959,G36684,G14958);
  or GNAME14960(G14960,G36694,G14959);
  or GNAME14961(G14961,G36682,G14960);
  or GNAME14962(G14962,G36701,G14961);
  or GNAME14963(G14963,G36688,G14962);
  or GNAME14964(G14964,G36692,G14963);
  or GNAME14965(G14965,G36677,G14964);
  or GNAME14966(G14966,G36703,G14965);
  nor GNAME14967(G14967,G36697,G14966);
  nand GNAME14968(G14968,G14947,G36686);
  nand GNAME14969(G14969,G14946,G36696);
  nand GNAME14970(G14970,G14945,G36704);
  nand GNAME14971(G14971,G14944,G36678);
  nand GNAME14972(G14972,G14943,G36690);
  nand GNAME14973(G14973,G36699,G36687);
  and GNAME14974(G14974,G14966,G36697);
  nand GNAME14975(G14975,G14965,G36703);
  nand GNAME14976(G14976,G14964,G36677);
  nand GNAME14977(G14977,G14963,G36692);
  nand GNAME14978(G14978,G14962,G36688);
  nand GNAME14979(G14979,G14961,G36701);
  nand GNAME14980(G14980,G14960,G36682);
  nand GNAME14981(G14981,G14959,G36694);
  nand GNAME14982(G14982,G14958,G36684);
  nand GNAME14983(G14983,G14957,G36698);
  nand GNAME14984(G14984,G14956,G36679);
  nand GNAME14985(G14985,G14955,G36689);
  nand GNAME14986(G14986,G14954,G36691);
  nand GNAME14987(G14987,G14953,G36676);
  nand GNAME14988(G14988,G14952,G36702);
  nand GNAME14989(G14989,G14951,G36683);
  nand GNAME14990(G14990,G14950,G36693);
  nand GNAME14991(G14991,G14949,G36681);
  nand GNAME14992(G14992,G14948,G36700);
  nand GNAME14993(G14993,G1191,G1192);
  not GNAME14994(G14994,G7733);
  not GNAME14995(G14995,G7760);
  not GNAME14996(G14996,G7731);
  not GNAME14997(G14997,G7746);
  not GNAME14998(G14998,G7738);
  not GNAME14999(G14999,G7744);
  not GNAME15000(G15000,G7737);
  not GNAME15001(G15001,G7742);
  not GNAME15002(G15002,G7740);
  not GNAME15003(G15003,G7770);
  not GNAME15004(G15004,G7723);
  not GNAME15005(G15005,G7768);
  not GNAME15006(G15006,G7725);
  not GNAME15007(G15007,G7766);
  not GNAME15008(G15008,G7722);
  not GNAME15009(G15009,G7764);
  not GNAME15010(G15010,G7728);
  not GNAME15011(G15011,G7762);
  not GNAME15012(G15012,G7729);
  not GNAME15013(G15013,G7759);
  not GNAME15014(G15014,G7567);
  not GNAME15015(G15015,G7757);
  not GNAME15016(G15016,G7569);
  not GNAME15017(G15017,G7755);
  not GNAME15018(G15018,G7571);
  not GNAME15019(G15019,G7753);
  not GNAME15020(G15020,G7573);
  not GNAME15021(G15021,G7751);
  not GNAME15022(G15022,G7575);
  not GNAME15023(G15023,G7748);
  not GNAME15024(G15024,G7579);
  not GNAME15025(G15025,G7772);
  nand GNAME15026(G15026,G14994,G7771);
  nand GNAME15027(G15027,G7721,G15025,G15026);
  or GNAME15028(G15028,G7771,G14994);
  nand GNAME15029(G15029,G14995,G7735);
  nand GNAME15030(G15030,G15029,G15027,G15028);
  or GNAME15031(G15031,G7735,G14995);
  nand GNAME15032(G15032,G14996,G7749);
  nand GNAME15033(G15033,G15032,G15030,G15031);
  or GNAME15034(G15034,G7749,G14996);
  nand GNAME15035(G15035,G14997,G7734);
  nand GNAME15036(G15036,G15035,G15033,G15034);
  or GNAME15037(G15037,G7734,G14997);
  nand GNAME15038(G15038,G14998,G7745);
  nand GNAME15039(G15039,G15038,G15036,G15037);
  or GNAME15040(G15040,G7745,G14998);
  nand GNAME15041(G15041,G14999,G7736);
  nand GNAME15042(G15042,G15041,G15039,G15040);
  or GNAME15043(G15043,G7736,G14999);
  nand GNAME15044(G15044,G15000,G7743);
  nand GNAME15045(G15045,G15044,G15042,G15043);
  or GNAME15046(G15046,G7743,G15000);
  nand GNAME15047(G15047,G15001,G7732);
  nand GNAME15048(G15048,G15047,G15045,G15046);
  or GNAME15049(G15049,G7732,G15001);
  nand GNAME15050(G15050,G15002,G7741);
  nand GNAME15051(G15051,G15050,G15048,G15049);
  or GNAME15052(G15052,G7741,G15002);
  nand GNAME15053(G15053,G15003,G7739);
  nand GNAME15054(G15054,G15053,G15051,G15052);
  or GNAME15055(G15055,G7739,G15003);
  nand GNAME15056(G15056,G15004,G7769);
  nand GNAME15057(G15057,G15056,G15054,G15055);
  or GNAME15058(G15058,G7769,G15004);
  nand GNAME15059(G15059,G15005,G7727);
  nand GNAME15060(G15060,G15059,G15057,G15058);
  or GNAME15061(G15061,G7727,G15005);
  nand GNAME15062(G15062,G15006,G7767);
  nand GNAME15063(G15063,G15062,G15060,G15061);
  or GNAME15064(G15064,G7767,G15006);
  nand GNAME15065(G15065,G15007,G7724);
  nand GNAME15066(G15066,G15065,G15063,G15064);
  or GNAME15067(G15067,G7724,G15007);
  nand GNAME15068(G15068,G15008,G7765);
  nand GNAME15069(G15069,G15068,G15066,G15067);
  or GNAME15070(G15070,G7765,G15008);
  nand GNAME15071(G15071,G15009,G7726);

endmodule