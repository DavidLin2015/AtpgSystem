module b17s(CK,G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33,G34,G35,G36,G37,G59244,G59243,G59242,G59241,G59240,G59239,G59238,G59237,G59236,G59235,G59234,G59233,G59232,G59231,G59230,G59229,G59228,G59227,G59226,G59225,G59224,G59223,G59222,G59221,G59220,G59219,G59218,G59217,G59216,G59215,G59214,G59213,G59809,G59810,G59811,G59812,G59813,G59814,G59815,G59816,G59817,G59818,G59819,G59820,G59821,G59822,G59823,G59824,G59825,G59826,G59827,G59828,G59829,G59830,G59831,G59832,G59833,G59834,G59835,G59836,G59837,G59838,G1700,G1701,G1702,G1703,G1704,G1705,G1706,G1707,G1708,G1709,G1711,G1712,G1713,G1714,G1715,G1716,G1717,G1718,G1719,G1720,G1692,G1693,G1694,G1695,G1696,G1697,G1698,G1699,G1710,G1721,G59345,G59350,G59351,G60251,G59353);
input CK,G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33,G34,G35,G36,G37;
output G59244,G59243,G59242,G59241,G59240,G59239,G59238,G59237,G59236,G59235,G59234,G59233,G59232,G59231,G59230,G59229,G59228,G59227,G59226,G59225,G59224,G59223,G59222,G59221,G59220,G59219,G59218,G59217,G59216,G59215,G59214,G59213,G59809,G59810,G59811,G59812,G59813,G59814,G59815,G59816,G59817,G59818,G59819,G59820,G59821,G59822,G59823,G59824,G59825,G59826,G59827,G59828,G59829,G59830,G59831,G59832,G59833,G59834,G59835,G59836,G59837,G59838,G1700,G1701,G1702,G1703,G1704,G1705,G1706,G1707,G1708,G1709,G1711,G1712,G1713,G1714,G1715,G1716,G1717,G1718,G1719,G1720,G1692,G1693,G1694,G1695,G1696,G1697,G1698,G1699,G1710,G1721,G59345,G59350,G59351,G60251,G59353;

  wire G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,
       G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,G40,
       G41,G42,G43,G44,G45,G46,G47,G48,G49,G50,G51,G52,G53,G54,G55,G56,G57,G58,G59,G60,
       G61,G62,G63,G64,G65,G66,G67,G68,G69,G70,G71,G72,G73,G74,G75,G76,G77,G78,G79,G80,
       G81,G82,G83,G84,G85,G86,G87,G88,G89,G90,G91,G92,G93,G94,G95,G96,G97,G98,G99,G100,
       G101,G102,G103,G104,G105,G106,G107,G108,G109,G110,G111,G112,G113,G114,G115,G116,G117,G118,G119,G120,
       G121,G122,G123,G124,G125,G126,G127,G128,G129,G130,G131,G132,G133,G134,G135,G136,G137,G138,G139,G140,
       G141,G142,G143,G144,G145,G146,G147,G148,G149,G150,G151,G152,G153,G154,G155,G156,G157,G158,G159,G160,
       G161,G162,G163,G164,G165,G166,G167,G168,G169,G170,G171,G172,G173,G174,G175,G176,G177,G178,G179,G180,
       G181,G182,G183,G184,G185,G186,G187,G188,G189,G190,G191,G192,G193,G194,G195,G196,G197,G198,G199,G200,
       G201,G202,G203,G204,G205,G206,G207,G208,G209,G210,G211,G212,G213,G214,G215,G216,G217,G218,G219,G220,
       G221,G222,G223,G224,G225,G226,G227,G228,G229,G230,G231,G232,G233,G234,G235,G236,G237,G238,G239,G240,
       G241,G242,G243,G244,G245,G246,G247,G248,G249,G250,G251,G252,G253,G254,G255,G256,G257,G258,G259,G260,
       G261,G262,G263,G264,G265,G266,G267,G268,G269,G270,G271,G272,G273,G274,G275,G276,G277,G278,G279,G280,
       G281,G282,G283,G284,G285,G286,G287,G288,G289,G290,G291,G292,G293,G294,G295,G296,G297,G298,G299,G300,
       G301,G302,G303,G304,G305,G306,G307,G308,G309,G310,G311,G312,G313,G314,G315,G316,G317,G318,G319,G320,
       G321,G322,G323,G324,G325,G326,G327,G328,G329,G330,G331,G332,G333,G334,G335,G336,G337,G338,G339,G340,
       G341,G342,G343,G344,G345,G346,G347,G348,G349,G350,G351,G352,G353,G354,G355,G356,G357,G358,G359,G360,
       G361,G362,G363,G364,G365,G366,G367,G368,G369,G370,G371,G372,G373,G374,G375,G376,G377,G378,G379,G380,
       G381,G382,G383,G384,G385,G386,G387,G388,G389,G390,G391,G392,G393,G394,G395,G396,G397,G398,G399,G400,
       G401,G402,G403,G404,G405,G406,G407,G408,G409,G410,G411,G412,G413,G414,G415,G416,G417,G418,G419,G420,
       G421,G422,G423,G424,G425,G426,G427,G428,G429,G430,G431,G432,G433,G434,G435,G436,G437,G438,G439,G440,
       G441,G442,G443,G444,G445,G446,G447,G448,G449,G450,G451,G452,G453,G454,G455,G456,G457,G458,G459,G460,
       G461,G462,G463,G464,G465,G466,G467,G468,G469,G470,G471,G472,G473,G474,G475,G476,G477,G478,G479,G480,
       G481,G482,G483,G484,G485,G486,G487,G488,G489,G490,G491,G492,G493,G494,G495,G496,G497,G498,G499,G500,
       G501,G502,G503,G504,G505,G506,G507,G508,G509,G510,G511,G512,G513,G514,G515,G516,G517,G518,G519,G520,
       G521,G522,G523,G524,G525,G526,G527,G528,G529,G530,G531,G532,G533,G534,G535,G536,G537,G538,G539,G540,
       G541,G542,G543,G544,G545,G546,G547,G548,G549,G550,G551,G552,G553,G554,G555,G556,G557,G558,G559,G560,
       G561,G562,G563,G564,G565,G566,G567,G568,G569,G570,G571,G572,G573,G574,G575,G576,G577,G578,G579,G580,
       G581,G582,G583,G584,G585,G586,G587,G588,G589,G590,G591,G592,G593,G594,G595,G596,G597,G598,G599,G600,
       G601,G602,G603,G604,G605,G606,G607,G608,G609,G610,G611,G612,G613,G614,G615,G616,G617,G618,G619,G620,
       G621,G622,G623,G624,G625,G626,G627,G628,G629,G630,G631,G632,G633,G634,G635,G636,G637,G638,G639,G640,
       G641,G642,G643,G644,G645,G646,G647,G648,G649,G650,G651,G652,G653,G654,G655,G656,G657,G658,G659,G660,
       G661,G662,G663,G664,G665,G666,G667,G668,G669,G670,G671,G672,G673,G674,G675,G676,G677,G678,G679,G680,
       G681,G682,G683,G684,G685,G686,G687,G688,G689,G690,G691,G692,G693,G694,G695,G696,G697,G698,G699,G700,
       G701,G702,G703,G704,G705,G706,G707,G708,G709,G710,G711,G712,G713,G714,G715,G716,G717,G718,G719,G720,
       G721,G722,G723,G724,G725,G726,G727,G728,G729,G730,G731,G732,G733,G734,G735,G736,G737,G738,G739,G740,
       G741,G742,G743,G744,G745,G746,G747,G748,G749,G750,G751,G752,G753,G754,G755,G756,G757,G758,G759,G760,
       G761,G762,G763,G764,G765,G766,G767,G768,G769,G770,G771,G772,G773,G774,G775,G776,G777,G778,G779,G780,
       G781,G782,G783,G784,G785,G786,G787,G788,G789,G790,G791,G792,G793,G794,G795,G796,G797,G798,G799,G800,
       G801,G802,G803,G804,G805,G806,G807,G808,G809,G810,G811,G812,G813,G814,G815,G816,G817,G818,G819,G820,
       G821,G822,G823,G824,G825,G826,G827,G828,G829,G830,G831,G832,G833,G834,G835,G836,G837,G838,G839,G840,
       G841,G842,G843,G844,G845,G846,G847,G848,G849,G850,G851,G852,G853,G854,G855,G856,G857,G858,G859,G860,
       G861,G862,G863,G864,G865,G866,G867,G868,G869,G870,G871,G872,G873,G874,G875,G876,G877,G878,G879,G880,
       G881,G882,G883,G884,G885,G886,G887,G888,G889,G890,G891,G892,G893,G894,G895,G896,G897,G898,G899,G900,
       G901,G902,G903,G904,G905,G906,G907,G908,G909,G910,G911,G912,G913,G914,G915,G916,G917,G918,G919,G920,
       G921,G922,G923,G924,G925,G926,G927,G928,G929,G930,G931,G932,G933,G934,G935,G936,G937,G938,G939,G940,
       G941,G942,G943,G944,G945,G946,G947,G948,G949,G950,G951,G952,G953,G954,G955,G956,G957,G958,G959,G960,
       G961,G962,G963,G964,G965,G966,G967,G968,G969,G970,G971,G972,G973,G974,G975,G976,G977,G978,G979,G980,
       G981,G982,G983,G984,G985,G986,G987,G988,G989,G990,G991,G992,G993,G994,G995,G996,G997,G998,G999,G1000,
       G1001,G1002,G1003,G1004,G1005,G1006,G1007,G1008,G1009,G1010,G1011,G1012,G1013,G1014,G1015,G1016,G1017,G1018,G1019,G1020,
       G1021,G1022,G1023,G1024,G1025,G1026,G1027,G1028,G1029,G1030,G1031,G1032,G1033,G1034,G1035,G1036,G1037,G1038,G1039,G1040,
       G1041,G1042,G1043,G1044,G1045,G1046,G1047,G1048,G1049,G1050,G1051,G1052,G1053,G1054,G1055,G1056,G1057,G1058,G1059,G1060,
       G1061,G1062,G1063,G1064,G1065,G1066,G1067,G1068,G1069,G1070,G1071,G1072,G1073,G1074,G1075,G1076,G1077,G1078,G1079,G1080,
       G1081,G1082,G1083,G1084,G1085,G1086,G1087,G1088,G1089,G1090,G1091,G1092,G1093,G1094,G1095,G1096,G1097,G1098,G1099,G1100,
       G1101,G1102,G1103,G1104,G1105,G1106,G1107,G1108,G1109,G1110,G1111,G1112,G1113,G1114,G1115,G1116,G1117,G1118,G1119,G1120,
       G1121,G1122,G1123,G1124,G1125,G1126,G1127,G1128,G1129,G1130,G1131,G1132,G1133,G1134,G1135,G1136,G1137,G1138,G1139,G1140,
       G1141,G1142,G1143,G1144,G1145,G1146,G1147,G1148,G1149,G1150,G1151,G1152,G1153,G1154,G1155,G1156,G1157,G1158,G1159,G1160,
       G1161,G1162,G1163,G1164,G1165,G1166,G1167,G1168,G1169,G1170,G1171,G1172,G1173,G1174,G1175,G1176,G1177,G1178,G1179,G1180,
       G1181,G1182,G1183,G1184,G1185,G1186,G1187,G1188,G1189,G1190,G1191,G1192,G1193,G1194,G1195,G1196,G1197,G1198,G1199,G1200,
       G1201,G1202,G1203,G1204,G1205,G1206,G1207,G1208,G1209,G1210,G1211,G1212,G1213,G1214,G1215,G1216,G1217,G1218,G1219,G1220,
       G1221,G1222,G1223,G1224,G1225,G1226,G1227,G1228,G1229,G1230,G1231,G1232,G1233,G1234,G1235,G1236,G1237,G1238,G1239,G1240,
       G1241,G1242,G1243,G1244,G1245,G1246,G1247,G1248,G1249,G1250,G1251,G1252,G1253,G1254,G1255,G1256,G1257,G1258,G1259,G1260,
       G1261,G1262,G1263,G1264,G1265,G1266,G1267,G1268,G1269,G1270,G1271,G1272,G1273,G1274,G1275,G1276,G1277,G1278,G1279,G1280,
       G1281,G1282,G1283,G1284,G1285,G1286,G1287,G1288,G1289,G1290,G1291,G1292,G1293,G1294,G1295,G1296,G1297,G1298,G1299,G1300,
       G1301,G1302,G1303,G1304,G1305,G1306,G1307,G1308,G1309,G1310,G1311,G1312,G1313,G1314,G1315,G1316,G1317,G1318,G1319,G1320,
       G1321,G1322,G1323,G1324,G1325,G1326,G1327,G1328,G1329,G1330,G1331,G1332,G1333,G1334,G1335,G1336,G1337,G1338,G1339,G1340,
       G1341,G1342,G1343,G1344,G1345,G1346,G1347,G1348,G1349,G1350,G1351,G1352,G1353,G1354,G1355,G1356,G1357,G1358,G1359,G1360,
       G1361,G1362,G1363,G1364,G1365,G1366,G1367,G1368,G1369,G1370,G1371,G1372,G1373,G1374,G1375,G1376,G1377,G1378,G1379,G1380,
       G1381,G1382,G1383,G1384,G1385,G1386,G1387,G1388,G1389,G1390,G1391,G1392,G1393,G1394,G1395,G1396,G1397,G1398,G1399,G1400,
       G1401,G1402,G1403,G1404,G1405,G1406,G1407,G1408,G1409,G1410,G1411,G1412,G1413,G1414,G1415,G1416,G1417,G1418,G1419,G1420,
       G1421,G1422,G1423,G1424,G1425,G1426,G1427,G1428,G1429,G1430,G1431,G1432,G1433,G1434,G1435,G1436,G1437,G1438,G1439,G1440,
       G1441,G1442,G1443,G1444,G1445,G1446,G1447,G1448,G1449,G1450,G1451,G1452,G1453,G1454,G1455,G1456,G1457,G1458,G1459,G1460,
       G1461,G1462,G1463,G1464,G1465,G1466,G1467,G1468,G1469,G1470,G1471,G1472,G1473,G1474,G1475,G1476,G1477,G1478,G1479,G1480,
       G1481,G1482,G1483,G1484,G1485,G1486,G1487,G1488,G1489,G1490,G1491,G1492,G1493,G1494,G1495,G1496,G1497,G1498,G1499,G1500,
       G1501,G1502,G1503,G1504,G1505,G1506,G1507,G1508,G1509,G1510,G1511,G1512,G1513,G1514,G1515,G1516,G1517,G1518,G1519,G1520,
       G1521,G1522,G1523,G1524,G1525,G1526,G1527,G1528,G1529,G1530,G1531,G1532,G1533,G1534,G1535,G1536,G1537,G1538,G1539,G1540,
       G1541,G1542,G1543,G1544,G1545,G1546,G1547,G1548,G1549,G1550,G1551,G1552,G1553,G1554,G1555,G1556,G1557,G1558,G1559,G1560,
       G1561,G1562,G1563,G1564,G1565,G1566,G1567,G1568,G1569,G1570,G1571,G1572,G1573,G1574,G1575,G1576,G1577,G1578,G1579,G1580,
       G1581,G1582,G1583,G1584,G1585,G1586,G1587,G1588,G1589,G1590,G1591,G1592,G1593,G1594,G1595,G1596,G1597,G1598,G1599,G1600,
       G1601,G1602,G1603,G1604,G1605,G1606,G1607,G1608,G1609,G1610,G1611,G1612,G1613,G1614,G1615,G1616,G1617,G1618,G1619,G1620,
       G1621,G1622,G1623,G1624,G1625,G1626,G1627,G1628,G1629,G1630,G1631,G1632,G1633,G1634,G1635,G1636,G1637,G1638,G1639,G1640,
       G1641,G1642,G1643,G1644,G1645,G1646,G1647,G1648,G1649,G1650,G1651,G1652,G1653,G1654,G1655,G1656,G1657,G1658,G1659,G1660,
       G1661,G1662,G1663,G1664,G1665,G1666,G1667,G1668,G1669,G1670,G1671,G1672,G1673,G1674,G1675,G1676,G1677,G1678,G1679,G1680,
       G1681,G1682,G1683,G1684,G1685,G1686,G1687,G1688,G1689,G1690,G1691,G1692,G1693,G1694,G1695,G1696,G1697,G1698,G1699,G1700,
       G1701,G1702,G1703,G1704,G1705,G1706,G1707,G1708,G1709,G1710,G1711,G1712,G1713,G1714,G1715,G1716,G1717,G1718,G1719,G1720,
       G1721,G1722,G1723,G1724,G1725,G1726,G1727,G1728,G1729,G1730,G1731,G1732,G1733,G1734,G1735,G1736,G1737,G1738,G1739,G1740,
       G1741,G1742,G1743,G1744,G1745,G1746,G1747,G1748,G1749,G1750,G1751,G1752,G1753,G1754,G1755,G1756,G1757,G1758,G1759,G1760,
       G1761,G1762,G1763,G1764,G1765,G1766,G1767,G1768,G1769,G1770,G1771,G1772,G1773,G1774,G1775,G1776,G1777,G1778,G1779,G1780,
       G1781,G1782,G1783,G1784,G1785,G1786,G1787,G1788,G1789,G1790,G1791,G1792,G1793,G1794,G1795,G1796,G1797,G1798,G1799,G1800,
       G1801,G1802,G1803,G1804,G1805,G1806,G1807,G1808,G1809,G1810,G1811,G1812,G1813,G1814,G1815,G1816,G1817,G1818,G1819,G1820,
       G1821,G1822,G1823,G1824,G1825,G1826,G1827,G1828,G1829,G1830,G1831,G1832,G1833,G1834,G1835,G1836,G1837,G1838,G1839,G1840,
       G1841,G1842,G1843,G1844,G1845,G1846,G1847,G1848,G1849,G1850,G1851,G1852,G1853,G1854,G1855,G1856,G1857,G1858,G1859,G1860,
       G1861,G1862,G1863,G1864,G1865,G1866,G1867,G1868,G1869,G1870,G1871,G1872,G1873,G1874,G1875,G1876,G1877,G1878,G1879,G1880,
       G1881,G1882,G1883,G1884,G1885,G1886,G1887,G1888,G1889,G1890,G1891,G1892,G1893,G1894,G1895,G1896,G1897,G1898,G1899,G1900,
       G1901,G1902,G1903,G1904,G1905,G1906,G1907,G1908,G1909,G1910,G1911,G1912,G1913,G1914,G1915,G1916,G1917,G1918,G1919,G1920,
       G1921,G1922,G1923,G1924,G1925,G1926,G1927,G1928,G1929,G1930,G1931,G1932,G1933,G1934,G1935,G1936,G1937,G1938,G1939,G1940,
       G1941,G1942,G1943,G1944,G1945,G1946,G1947,G1948,G1949,G1950,G1951,G1952,G1953,G1954,G1955,G1956,G1957,G1958,G1959,G1960,
       G1961,G1962,G1963,G1964,G1965,G1966,G1967,G1968,G1969,G1970,G1971,G1972,G1973,G1974,G1975,G1976,G1977,G1978,G1979,G1980,
       G1981,G1982,G1983,G1984,G1985,G1986,G1987,G1988,G1989,G1990,G1991,G1992,G1993,G1994,G1995,G1996,G1997,G1998,G1999,G2000,
       G2001,G2002,G2003,G2004,G2005,G2006,G2007,G2008,G2009,G2010,G2011,G2012,G2013,G2014,G2015,G2016,G2017,G2018,G2019,G2020,
       G2021,G2022,G2023,G2024,G2025,G2026,G2027,G2028,G2029,G2030,G2031,G2032,G2033,G2034,G2035,G2036,G2037,G2038,G2039,G2040,
       G2041,G2042,G2043,G2044,G2045,G2046,G2047,G2048,G2049,G2050,G2051,G2052,G2053,G2054,G2055,G2056,G2057,G2058,G2059,G2060,
       G2061,G2062,G2063,G2064,G2065,G2066,G2067,G2068,G2069,G2070,G2071,G2072,G2073,G2074,G2075,G2076,G2077,G2078,G2079,G2080,
       G2081,G2082,G2083,G2084,G2085,G2086,G2087,G2088,G2089,G2090,G2091,G2092,G2093,G2094,G2095,G2096,G2097,G2098,G2099,G2100,
       G2101,G2102,G2103,G2104,G2105,G2106,G2107,G2108,G2109,G2110,G2111,G2112,G2113,G2114,G2115,G2116,G2117,G2118,G2119,G2120,
       G2121,G2122,G2123,G2124,G2125,G2126,G2127,G2128,G2129,G2130,G2131,G2132,G2133,G2134,G2135,G2136,G2137,G2138,G2139,G2140,
       G2141,G2142,G2143,G2144,G2145,G2146,G2147,G2148,G2149,G2150,G2151,G2152,G2153,G2154,G2155,G2156,G2157,G2158,G2159,G2160,
       G2161,G2162,G2163,G2164,G2165,G2166,G2167,G2168,G2169,G2170,G2171,G2172,G2173,G2174,G2175,G2176,G2177,G2178,G2179,G2180,
       G2181,G2182,G2183,G2184,G2185,G2186,G2187,G2188,G2189,G2190,G2191,G2192,G2193,G2194,G2195,G2196,G2197,G2198,G2199,G2200,
       G2201,G2202,G2203,G2204,G2205,G2206,G2207,G2208,G2209,G2210,G2211,G2212,G2213,G2214,G2215,G2216,G2217,G2218,G2219,G2220,
       G2221,G2222,G2223,G2224,G2225,G2226,G2227,G2228,G2229,G2230,G2231,G2232,G2233,G2234,G2235,G2236,G2237,G2238,G2239,G2240,
       G2241,G2242,G2243,G2244,G2245,G2246,G2247,G2248,G2249,G2250,G2251,G2252,G2253,G2254,G2255,G2256,G2257,G2258,G2259,G2260,
       G2261,G2262,G2263,G2264,G2265,G2266,G2267,G2268,G2269,G2270,G2271,G2272,G2273,G2274,G2275,G2276,G2277,G2278,G2279,G2280,
       G2281,G2282,G2283,G2284,G2285,G2286,G2287,G2288,G2289,G2290,G2291,G2292,G2293,G2294,G2295,G2296,G2297,G2298,G2299,G2300,
       G2301,G2302,G2303,G2304,G2305,G2306,G2307,G2308,G2309,G2310,G2311,G2312,G2313,G2314,G2315,G2316,G2317,G2318,G2319,G2320,
       G2321,G2322,G2323,G2324,G2325,G2326,G2327,G2328,G2329,G2330,G2331,G2332,G2333,G2334,G2335,G2336,G2337,G2338,G2339,G2340,
       G2341,G2342,G2343,G2344,G2345,G2346,G2347,G2348,G2349,G2350,G2351,G2352,G2353,G2354,G2355,G2356,G2357,G2358,G2359,G2360,
       G2361,G2362,G2363,G2364,G2365,G2366,G2367,G2368,G2369,G2370,G2371,G2372,G2373,G2374,G2375,G2376,G2377,G2378,G2379,G2380,
       G2381,G2382,G2383,G2384,G2385,G2386,G2387,G2388,G2389,G2390,G2391,G2392,G2393,G2394,G2395,G2396,G2397,G2398,G2399,G2400,
       G2401,G2402,G2403,G2404,G2405,G2406,G2407,G2408,G2409,G2410,G2411,G2412,G2413,G2414,G2415,G2416,G2417,G2418,G2419,G2420,
       G2421,G2422,G2423,G2424,G2425,G2426,G2427,G2428,G2429,G2430,G2431,G2432,G2433,G2434,G2435,G2436,G2437,G2438,G2439,G2440,
       G2441,G2442,G2443,G2444,G2445,G2446,G2447,G2448,G2449,G2450,G2451,G2452,G2453,G2454,G2455,G2456,G2457,G2458,G2459,G2460,
       G2461,G2462,G2463,G2464,G2465,G2466,G2467,G2468,G2469,G2470,G2471,G2472,G2473,G2474,G2475,G2476,G2477,G2478,G2479,G2480,
       G2481,G2482,G2483,G2484,G2485,G2486,G2487,G2488,G2489,G2490,G2491,G2492,G2493,G2494,G2495,G2496,G2497,G2498,G2499,G2500,
       G2501,G2502,G2503,G2504,G2505,G2506,G2507,G2508,G2509,G2510,G2511,G2512,G2513,G2514,G2515,G2516,G2517,G2518,G2519,G2520,
       G2521,G2522,G2523,G2524,G2525,G2526,G2527,G2528,G2529,G2530,G2531,G2532,G2533,G2534,G2535,G2536,G2537,G2538,G2539,G2540,
       G2541,G2542,G2543,G2544,G2545,G2546,G2547,G2548,G2549,G2550,G2551,G2552,G2553,G2554,G2555,G2556,G2557,G2558,G2559,G2560,
       G2561,G2562,G2563,G2564,G2565,G2566,G2567,G2568,G2569,G2570,G2571,G2572,G2573,G2574,G2575,G2576,G2577,G2578,G2579,G2580,
       G2581,G2582,G2583,G2584,G2585,G2586,G2587,G2588,G2589,G2590,G2591,G2592,G2593,G2594,G2595,G2596,G2597,G2598,G2599,G2600,
       G2601,G2602,G2603,G2604,G2605,G2606,G2607,G2608,G2609,G2610,G2611,G2612,G2613,G2614,G2615,G2616,G2617,G2618,G2619,G2620,
       G2621,G2622,G2623,G2624,G2625,G2626,G2627,G2628,G2629,G2630,G2631,G2632,G2633,G2634,G2635,G2636,G2637,G2638,G2639,G2640,
       G2641,G2642,G2643,G2644,G2645,G2646,G2647,G2648,G2649,G2650,G2651,G2652,G2653,G2654,G2655,G2656,G2657,G2658,G2659,G2660,
       G2661,G2662,G2663,G2664,G2665,G2666,G2667,G2668,G2669,G2670,G2671,G2672,G2673,G2674,G2675,G2676,G2677,G2678,G2679,G2680,
       G2681,G2682,G2683,G2684,G2685,G2686,G2687,G2688,G2689,G2690,G2691,G2692,G2693,G2694,G2695,G2696,G2697,G2698,G2699,G2700,
       G2701,G2702,G2703,G2704,G2705,G2706,G2707,G2708,G2709,G2710,G2711,G2712,G2713,G2714,G2715,G2716,G2717,G2718,G2719,G2720,
       G2721,G2722,G2723,G2724,G2725,G2726,G2727,G2728,G2729,G2730,G2731,G2732,G2733,G2734,G2735,G2736,G2737,G2738,G2739,G2740,
       G2741,G2742,G2743,G2744,G2745,G2746,G2747,G2748,G2749,G2750,G2751,G2752,G2753,G2754,G2755,G2756,G2757,G2758,G2759,G2760,
       G2761,G2762,G2763,G2764,G2765,G2766,G2767,G2768,G2769,G2770,G2771,G2772,G2773,G2774,G2775,G2776,G2777,G2778,G2779,G2780,
       G2781,G2782,G2783,G2784,G2785,G2786,G2787,G2788,G2789,G2790,G2791,G2792,G2793,G2794,G2795,G2796,G2797,G2798,G2799,G2800,
       G2801,G2802,G2803,G2804,G2805,G2806,G2807,G2808,G2809,G2810,G2811,G2812,G2813,G2814,G2815,G2816,G2817,G2818,G2819,G2820,
       G2821,G2822,G2823,G2824,G2825,G2826,G2827,G2828,G2829,G2830,G2831,G2832,G2833,G2834,G2835,G2836,G2837,G2838,G2839,G2840,
       G2841,G2842,G2843,G2844,G2845,G2846,G2847,G2848,G2849,G2850,G2851,G2852,G2853,G2854,G2855,G2856,G2857,G2858,G2859,G2860,
       G2861,G2862,G2863,G2864,G2865,G2866,G2867,G2868,G2869,G2870,G2871,G2872,G2873,G2874,G2875,G2876,G2877,G2878,G2879,G2880,
       G2881,G2882,G2883,G2884,G2885,G2886,G2887,G2888,G2889,G2890,G2891,G2892,G2893,G2894,G2895,G2896,G2897,G2898,G2899,G2900,
       G2901,G2902,G2903,G2904,G2905,G2906,G2907,G2908,G2909,G2910,G2911,G2912,G2913,G2914,G2915,G2916,G2917,G2918,G2919,G2920,
       G2921,G2922,G2923,G2924,G2925,G2926,G2927,G2928,G2929,G2930,G2931,G2932,G2933,G2934,G2935,G2936,G2937,G2938,G2939,G2940,
       G2941,G2942,G2943,G2944,G2945,G2946,G2947,G2948,G2949,G2950,G2951,G2952,G2953,G2954,G2955,G2956,G2957,G2958,G2959,G2960,
       G2961,G2962,G2963,G2964,G2965,G2966,G2967,G2968,G2969,G2970,G2971,G2972,G2973,G2974,G2975,G2976,G2977,G2978,G2979,G2980,
       G2981,G2982,G2983,G2984,G2985,G2986,G2987,G2988,G2989,G2990,G2991,G2992,G2993,G2994,G2995,G2996,G2997,G2998,G2999,G3000,
       G3001,G3002,G3003,G3004,G3005,G3006,G3007,G3008,G3009,G3010,G3011,G3012,G3013,G3014,G3015,G3016,G3017,G3018,G3019,G3020,
       G3021,G3022,G3023,G3024,G3025,G3026,G3027,G3028,G3029,G3030,G3031,G3032,G3033,G3034,G3035,G3036,G3037,G3038,G3039,G3040,
       G3041,G3042,G3043,G3044,G3045,G3046,G3047,G3048,G3049,G3050,G3051,G3052,G3053,G3054,G3055,G3056,G3057,G3058,G3059,G3060,
       G3061,G3062,G3063,G3064,G3065,G3066,G3067,G3068,G3069,G3070,G3071,G3072,G3073,G3074,G3075,G3076,G3077,G3078,G3079,G3080,
       G3081,G3082,G3083,G3084,G3085,G3086,G3087,G3088,G3089,G3090,G3091,G3092,G3093,G3094,G3095,G3096,G3097,G3098,G3099,G3100,
       G3101,G3102,G3103,G3104,G3105,G3106,G3107,G3108,G3109,G3110,G3111,G3112,G3113,G3114,G3115,G3116,G3117,G3118,G3119,G3120,
       G3121,G3122,G3123,G3124,G3125,G3126,G3127,G3128,G3129,G3130,G3131,G3132,G3133,G3134,G3135,G3136,G3137,G3138,G3139,G3140,
       G3141,G3142,G3143,G3144,G3145,G3146,G3147,G3148,G3149,G3150,G3151,G3152,G3153,G3154,G3155,G3156,G3157,G3158,G3159,G3160,
       G3161,G3162,G3163,G3164,G3165,G3166,G3167,G3168,G3169,G3170,G3171,G3172,G3173,G3174,G3175,G3176,G3177,G3178,G3179,G3180,
       G3181,G3182,G3183,G3184,G3185,G3186,G3187,G3188,G3189,G3190,G3191,G3192,G3193,G3194,G3195,G3196,G3197,G3198,G3199,G3200,
       G3201,G3202,G3203,G3204,G3205,G3206,G3207,G3208,G3209,G3210,G3211,G3212,G3213,G3214,G3215,G3216,G3217,G3218,G3219,G3220,
       G3221,G3222,G3223,G3224,G3225,G3226,G3227,G3228,G3229,G3230,G3231,G3232,G3233,G3234,G3235,G3236,G3237,G3238,G3239,G3240,
       G3241,G3242,G3243,G3244,G3245,G3246,G3247,G3248,G3249,G3250,G3251,G3252,G3253,G3254,G3255,G3256,G3257,G3258,G3259,G3260,
       G3261,G3262,G3263,G3264,G3265,G3266,G3267,G3268,G3269,G3270,G3271,G3272,G3273,G3274,G3275,G3276,G3277,G3278,G3279,G3280,
       G3281,G3282,G3283,G3284,G3285,G3286,G3287,G3288,G3289,G3290,G3291,G3292,G3293,G3294,G3295,G3296,G3297,G3298,G3299,G3300,
       G3301,G3302,G3303,G3304,G3305,G3306,G3307,G3308,G3309,G3310,G3311,G3312,G3313,G3314,G3315,G3316,G3317,G3318,G3319,G3320,
       G3321,G3322,G3323,G3324,G3325,G3326,G3327,G3328,G3329,G3330,G3331,G3332,G3333,G3334,G3335,G3336,G3337,G3338,G3339,G3340,
       G3341,G3342,G3343,G3344,G3345,G3346,G3347,G3348,G3349,G3350,G3351,G3352,G3353,G3354,G3355,G3356,G3357,G3358,G3359,G3360,
       G3361,G3362,G3363,G3364,G3365,G3366,G3367,G3368,G3369,G3370,G3371,G3372,G3373,G3374,G3375,G3376,G3377,G3378,G3379,G3380,
       G3381,G3382,G3383,G3384,G3385,G3386,G3387,G3388,G3389,G3390,G3391,G3392,G3393,G3394,G3395,G3396,G3397,G3398,G3399,G3400,
       G3401,G3402,G3403,G3404,G3405,G3406,G3407,G3408,G3409,G3410,G3411,G3412,G3413,G3414,G3415,G3416,G3417,G3418,G3419,G3420,
       G3421,G3422,G3423,G3424,G3425,G3426,G3427,G3428,G3429,G3430,G3431,G3432,G3433,G3434,G3435,G3436,G3437,G3438,G3439,G3440,
       G3441,G3442,G3443,G3444,G3445,G3446,G3447,G3448,G3449,G3450,G3451,G3452,G3453,G3454,G3455,G3456,G3457,G3458,G3459,G3460,
       G3461,G3462,G3463,G3464,G3465,G3466,G3467,G3468,G3469,G3470,G3471,G3472,G3473,G3474,G3475,G3476,G3477,G3478,G3479,G3480,
       G3481,G3482,G3483,G3484,G3485,G3486,G3487,G3488,G3489,G3490,G3491,G3492,G3493,G3494,G3495,G3496,G3497,G3498,G3499,G3500,
       G3501,G3502,G3503,G3504,G3505,G3506,G3507,G3508,G3509,G3510,G3511,G3512,G3513,G3514,G3515,G3516,G3517,G3518,G3519,G3520,
       G3521,G3522,G3523,G3524,G3525,G3526,G3527,G3528,G3529,G3530,G3531,G3532,G3533,G3534,G3535,G3536,G3537,G3538,G3539,G3540,
       G3541,G3542,G3543,G3544,G3545,G3546,G3547,G3548,G3549,G3550,G3551,G3552,G3553,G3554,G3555,G3556,G3557,G3558,G3559,G3560,
       G3561,G3562,G3563,G3564,G3565,G3566,G3567,G3568,G3569,G3570,G3571,G3572,G3573,G3574,G3575,G3576,G3577,G3578,G3579,G3580,
       G3581,G3582,G3583,G3584,G3585,G3586,G3587,G3588,G3589,G3590,G3591,G3592,G3593,G3594,G3595,G3596,G3597,G3598,G3599,G3600,
       G3601,G3602,G3603,G3604,G3605,G3606,G3607,G3608,G3609,G3610,G3611,G3612,G3613,G3614,G3615,G3616,G3617,G3618,G3619,G3620,
       G3621,G3622,G3623,G3624,G3625,G3626,G3627,G3628,G3629,G3630,G3631,G3632,G3633,G3634,G3635,G3636,G3637,G3638,G3639,G3640,
       G3641,G3642,G3643,G3644,G3645,G3646,G3647,G3648,G3649,G3650,G3651,G3652,G3653,G3654,G3655,G3656,G3657,G3658,G3659,G3660,
       G3661,G3662,G3663,G3664,G3665,G3666,G3667,G3668,G3669,G3670,G3671,G3672,G3673,G3674,G3675,G3676,G3677,G3678,G3679,G3680,
       G3681,G3682,G3683,G3684,G3685,G3686,G3687,G3688,G3689,G3690,G3691,G3692,G3693,G3694,G3695,G3696,G3697,G3698,G3699,G3700,
       G3701,G3702,G3703,G3704,G3705,G3706,G3707,G3708,G3709,G3710,G3711,G3712,G3713,G3714,G3715,G3716,G3717,G3718,G3719,G3720,
       G3721,G3722,G3723,G3724,G3725,G3726,G3727,G3728,G3729,G3730,G3731,G3732,G3733,G3734,G3735,G3736,G3737,G3738,G3739,G3740,
       G3741,G3742,G3743,G3744,G3745,G3746,G3747,G3748,G3749,G3750,G3751,G3752,G3753,G3754,G3755,G3756,G3757,G3758,G3759,G3760,
       G3761,G3762,G3763,G3764,G3765,G3766,G3767,G3768,G3769,G3770,G3771,G3772,G3773,G3774,G3775,G3776,G3777,G3778,G3779,G3780,
       G3781,G3782,G3783,G3784,G3785,G3786,G3787,G3788,G3789,G3790,G3791,G3792,G3793,G3794,G3795,G3796,G3797,G3798,G3799,G3800,
       G3801,G3802,G3803,G3804,G3805,G3806,G3807,G3808,G3809,G3810,G3811,G3812,G3813,G3814,G3815,G3816,G3817,G3818,G3819,G3820,
       G3821,G3822,G3823,G3824,G3825,G3826,G3827,G3828,G3829,G3830,G3831,G3832,G3833,G3834,G3835,G3836,G3837,G3838,G3839,G3840,
       G3841,G3842,G3843,G3844,G3845,G3846,G3847,G3848,G3849,G3850,G3851,G3852,G3853,G3854,G3855,G3856,G3857,G3858,G3859,G3860,
       G3861,G3862,G3863,G3864,G3865,G3866,G3867,G3868,G3869,G3870,G3871,G3872,G3873,G3874,G3875,G3876,G3877,G3878,G3879,G3880,
       G3881,G3882,G3883,G3884,G3885,G3886,G3887,G3888,G3889,G3890,G3891,G3892,G3893,G3894,G3895,G3896,G3897,G3898,G3899,G3900,
       G3901,G3902,G3903,G3904,G3905,G3906,G3907,G3908,G3909,G3910,G3911,G3912,G3913,G3914,G3915,G3916,G3917,G3918,G3919,G3920,
       G3921,G3922,G3923,G3924,G3925,G3926,G3927,G3928,G3929,G3930,G3931,G3932,G3933,G3934,G3935,G3936,G3937,G3938,G3939,G3940,
       G3941,G3942,G3943,G3944,G3945,G3946,G3947,G3948,G3949,G3950,G3951,G3952,G3953,G3954,G3955,G3956,G3957,G3958,G3959,G3960,
       G3961,G3962,G3963,G3964,G3965,G3966,G3967,G3968,G3969,G3970,G3971,G3972,G3973,G3974,G3975,G3976,G3977,G3978,G3979,G3980,
       G3981,G3982,G3983,G3984,G3985,G3986,G3987,G3988,G3989,G3990,G3991,G3992,G3993,G3994,G3995,G3996,G3997,G3998,G3999,G4000,
       G4001,G4002,G4003,G4004,G4005,G4006,G4007,G4008,G4009,G4010,G4011,G4012,G4013,G4014,G4015,G4016,G4017,G4018,G4019,G4020,
       G4021,G4022,G4023,G4024,G4025,G4026,G4027,G4028,G4029,G4030,G4031,G4032,G4033,G4034,G4035,G4036,G4037,G4038,G4039,G4040,
       G4041,G4042,G4043,G4044,G4045,G4046,G4047,G4048,G4049,G4050,G4051,G4052,G4053,G4054,G4055,G4056,G4057,G4058,G4059,G4060,
       G4061,G4062,G4063,G4064,G4065,G4066,G4067,G4068,G4069,G4070,G4071,G4072,G4073,G4074,G4075,G4076,G4077,G4078,G4079,G4080,
       G4081,G4082,G4083,G4084,G4085,G4086,G4087,G4088,G4089,G4090,G4091,G4092,G4093,G4094,G4095,G4096,G4097,G4098,G4099,G4100,
       G4101,G4102,G4103,G4104,G4105,G4106,G4107,G4108,G4109,G4110,G4111,G4112,G4113,G4114,G4115,G4116,G4117,G4118,G4119,G4120,
       G4121,G4122,G4123,G4124,G4125,G4126,G4127,G4128,G4129,G4130,G4131,G4132,G4133,G4134,G4135,G4136,G4137,G4138,G4139,G4140,
       G4141,G4142,G4143,G4144,G4145,G4146,G4147,G4148,G4149,G4150,G4151,G4152,G4153,G4154,G4155,G4156,G4157,G4158,G4159,G4160,
       G4161,G4162,G4163,G4164,G4165,G4166,G4167,G4168,G4169,G4170,G4171,G4172,G4173,G4174,G4175,G4176,G4177,G4178,G4179,G4180,
       G4181,G4182,G4183,G4184,G4185,G4186,G4187,G4188,G4189,G4190,G4191,G4192,G4193,G4194,G4195,G4196,G4197,G4198,G4199,G4200,
       G4201,G4202,G4203,G4204,G4205,G4206,G4207,G4208,G4209,G4210,G4211,G4212,G4213,G4214,G4215,G4216,G4217,G4218,G4219,G4220,
       G4221,G4222,G4223,G4224,G4225,G4226,G4227,G4228,G4229,G4230,G4231,G4232,G4233,G4234,G4235,G4236,G4237,G4238,G4239,G4240,
       G4241,G4242,G4243,G4244,G4245,G4246,G4247,G4248,G4249,G4250,G4251,G4252,G4253,G4254,G4255,G4256,G4257,G4258,G4259,G4260,
       G4261,G4262,G4263,G4264,G4265,G4266,G4267,G4268,G4269,G4270,G4271,G4272,G4273,G4274,G4275,G4276,G4277,G4278,G4279,G4280,
       G4281,G4282,G4283,G4284,G4285,G4286,G4287,G4288,G4289,G4290,G4291,G4292,G4293,G4294,G4295,G4296,G4297,G4298,G4299,G4300,
       G4301,G4302,G4303,G4304,G4305,G4306,G4307,G4308,G4309,G4310,G4311,G4312,G4313,G4314,G4315,G4316,G4317,G4318,G4319,G4320,
       G4321,G4322,G4323,G4324,G4325,G4326,G4327,G4328,G4329,G4330,G4331,G4332,G4333,G4334,G4335,G4336,G4337,G4338,G4339,G4340,
       G4341,G4342,G4343,G4344,G4345,G4346,G4347,G4348,G4349,G4350,G4351,G4352,G4353,G4354,G4355,G4356,G4357,G4358,G4359,G4360,
       G4361,G4362,G4363,G4364,G4365,G4366,G4367,G4368,G4369,G4370,G4371,G4372,G4373,G4374,G4375,G4376,G4377,G4378,G4379,G4380,
       G4381,G4382,G4383,G4384,G4385,G4386,G4387,G4388,G4389,G4390,G4391,G4392,G4393,G4394,G4395,G4396,G4397,G4398,G4399,G4400,
       G4401,G4402,G4403,G4404,G4405,G4406,G4407,G4408,G4409,G4410,G4411,G4412,G4413,G4414,G4415,G4416,G4417,G4418,G4419,G4420,
       G4421,G4422,G4423,G4424,G4425,G4426,G4427,G4428,G4429,G4430,G4431,G4432,G4433,G4434,G4435,G4436,G4437,G4438,G4439,G4440,
       G4441,G4442,G4443,G4444,G4445,G4446,G4447,G4448,G4449,G4450,G4451,G4452,G4453,G4454,G4455,G4456,G4457,G4458,G4459,G4460,
       G4461,G4462,G4463,G4464,G4465,G4466,G4467,G4468,G4469,G4470,G4471,G4472,G4473,G4474,G4475,G4476,G4477,G4478,G4479,G4480,
       G4481,G4482,G4483,G4484,G4485,G4486,G4487,G4488,G4489,G4490,G4491,G4492,G4493,G4494,G4495,G4496,G4497,G4498,G4499,G4500,
       G4501,G4502,G4503,G4504,G4505,G4506,G4507,G4508,G4509,G4510,G4511,G4512,G4513,G4514,G4515,G4516,G4517,G4518,G4519,G4520,
       G4521,G4522,G4523,G4524,G4525,G4526,G4527,G4528,G4529,G4530,G4531,G4532,G4533,G4534,G4535,G4536,G4537,G4538,G4539,G4540,
       G4541,G4542,G4543,G4544,G4545,G4546,G4547,G4548,G4549,G4550,G4551,G4552,G4553,G4554,G4555,G4556,G4557,G4558,G4559,G4560,
       G4561,G4562,G4563,G4564,G4565,G4566,G4567,G4568,G4569,G4570,G4571,G4572,G4573,G4574,G4575,G4576,G4577,G4578,G4579,G4580,
       G4581,G4582,G4583,G4584,G4585,G4586,G4587,G4588,G4589,G4590,G4591,G4592,G4593,G4594,G4595,G4596,G4597,G4598,G4599,G4600,
       G4601,G4602,G4603,G4604,G4605,G4606,G4607,G4608,G4609,G4610,G4611,G4612,G4613,G4614,G4615,G4616,G4617,G4618,G4619,G4620,
       G4621,G4622,G4623,G4624,G4625,G4626,G4627,G4628,G4629,G4630,G4631,G4632,G4633,G4634,G4635,G4636,G4637,G4638,G4639,G4640,
       G4641,G4642,G4643,G4644,G4645,G4646,G4647,G4648,G4649,G4650,G4651,G4652,G4653,G4654,G4655,G4656,G4657,G4658,G4659,G4660,
       G4661,G4662,G4663,G4664,G4665,G4666,G4667,G4668,G4669,G4670,G4671,G4672,G4673,G4674,G4675,G4676,G4677,G4678,G4679,G4680,
       G4681,G4682,G4683,G4684,G4685,G4686,G4687,G4688,G4689,G4690,G4691,G4692,G4693,G4694,G4695,G4696,G4697,G4698,G4699,G4700,
       G4701,G4702,G4703,G4704,G4705,G4706,G4707,G4708,G4709,G4710,G4711,G4712,G4713,G4714,G4715,G4716,G4717,G4718,G4719,G4720,
       G4721,G4722,G4723,G4724,G4725,G4726,G4727,G4728,G4729,G4730,G4731,G4732,G4733,G4734,G4735,G4736,G4737,G4738,G4739,G4740,
       G4741,G4742,G4743,G4744,G4745,G4746,G4747,G4748,G4749,G4750,G4751,G4752,G4753,G4754,G4755,G4756,G4757,G4758,G4759,G4760,
       G4761,G4762,G4763,G4764,G4765,G4766,G4767,G4768,G4769,G4770,G4771,G4772,G4773,G4774,G4775,G4776,G4777,G4778,G4779,G4780,
       G4781,G4782,G4783,G4784,G4785,G4786,G4787,G4788,G4789,G4790,G4791,G4792,G4793,G4794,G4795,G4796,G4797,G4798,G4799,G4800,
       G4801,G4802,G4803,G4804,G4805,G4806,G4807,G4808,G4809,G4810,G4811,G4812,G4813,G4814,G4815,G4816,G4817,G4818,G4819,G4820,
       G4821,G4822,G4823,G4824,G4825,G4826,G4827,G4828,G4829,G4830,G4831,G4832,G4833,G4834,G4835,G4836,G4837,G4838,G4839,G4840,
       G4841,G4842,G4843,G4844,G4845,G4846,G4847,G4848,G4849,G4850,G4851,G4852,G4853,G4854,G4855,G4856,G4857,G4858,G4859,G4860,
       G4861,G4862,G4863,G4864,G4865,G4866,G4867,G4868,G4869,G4870,G4871,G4872,G4873,G4874,G4875,G4876,G4877,G4878,G4879,G4880,
       G4881,G4882,G4883,G4884,G4885,G4886,G4887,G4888,G4889,G4890,G4891,G4892,G4893,G4894,G4895,G4896,G4897,G4898,G4899,G4900,
       G4901,G4902,G4903,G4904,G4905,G4906,G4907,G4908,G4909,G4910,G4911,G4912,G4913,G4914,G4915,G4916,G4917,G4918,G4919,G4920,
       G4921,G4922,G4923,G4924,G4925,G4926,G4927,G4928,G4929,G4930,G4931,G4932,G4933,G4934,G4935,G4936,G4937,G4938,G4939,G4940,
       G4941,G4942,G4943,G4944,G4945,G4946,G4947,G4948,G4949,G4950,G4951,G4952,G4953,G4954,G4955,G4956,G4957,G4958,G4959,G4960,
       G4961,G4962,G4963,G4964,G4965,G4966,G4967,G4968,G4969,G4970,G4971,G4972,G4973,G4974,G4975,G4976,G4977,G4978,G4979,G4980,
       G4981,G4982,G4983,G4984,G4985,G4986,G4987,G4988,G4989,G4990,G4991,G4992,G4993,G4994,G4995,G4996,G4997,G4998,G4999,G5000,
       G5001,G5002,G5003,G5004,G5005,G5006,G5007,G5008,G5009,G5010,G5011,G5012,G5013,G5014,G5015,G5016,G5017,G5018,G5019,G5020,
       G5021,G5022,G5023,G5024,G5025,G5026,G5027,G5028,G5029,G5030,G5031,G5032,G5033,G5034,G5035,G5036,G5037,G5038,G5039,G5040,
       G5041,G5042,G5043,G5044,G5045,G5046,G5047,G5048,G5049,G5050,G5051,G5052,G5053,G5054,G5055,G5056,G5057,G5058,G5059,G5060,
       G5061,G5062,G5063,G5064,G5065,G5066,G5067,G5068,G5069,G5070,G5071,G5072,G5073,G5074,G5075,G5076,G5077,G5078,G5079,G5080,
       G5081,G5082,G5083,G5084,G5085,G5086,G5087,G5088,G5089,G5090,G5091,G5092,G5093,G5094,G5095,G5096,G5097,G5098,G5099,G5100,
       G5101,G5102,G5103,G5104,G5105,G5106,G5107,G5108,G5109,G5110,G5111,G5112,G5113,G5114,G5115,G5116,G5117,G5118,G5119,G5120,
       G5121,G5122,G5123,G5124,G5125,G5126,G5127,G5128,G5129,G5130,G5131,G5132,G5133,G5134,G5135,G5136,G5137,G5138,G5139,G5140,
       G5141,G5142,G5143,G5144,G5145,G5146,G5147,G5148,G5149,G5150,G5151,G5152,G5153,G5154,G5155,G5156,G5157,G5158,G5159,G5160,
       G5161,G5162,G5163,G5164,G5165,G5166,G5167,G5168,G5169,G5170,G5171,G5172,G5173,G5174,G5175,G5176,G5177,G5178,G5179,G5180,
       G5181,G5182,G5183,G5184,G5185,G5186,G5187,G5188,G5189,G5190,G5191,G5192,G5193,G5194,G5195,G5196,G5197,G5198,G5199,G5200,
       G5201,G5202,G5203,G5204,G5205,G5206,G5207,G5208,G5209,G5210,G5211,G5212,G5213,G5214,G5215,G5216,G5217,G5218,G5219,G5220,
       G5221,G5222,G5223,G5224,G5225,G5226,G5227,G5228,G5229,G5230,G5231,G5232,G5233,G5234,G5235,G5236,G5237,G5238,G5239,G5240,
       G5241,G5242,G5243,G5244,G5245,G5246,G5247,G5248,G5249,G5250,G5251,G5252,G5253,G5254,G5255,G5256,G5257,G5258,G5259,G5260,
       G5261,G5262,G5263,G5264,G5265,G5266,G5267,G5268,G5269,G5270,G5271,G5272,G5273,G5274,G5275,G5276,G5277,G5278,G5279,G5280,
       G5281,G5282,G5283,G5284,G5285,G5286,G5287,G5288,G5289,G5290,G5291,G5292,G5293,G5294,G5295,G5296,G5297,G5298,G5299,G5300,
       G5301,G5302,G5303,G5304,G5305,G5306,G5307,G5308,G5309,G5310,G5311,G5312,G5313,G5314,G5315,G5316,G5317,G5318,G5319,G5320,
       G5321,G5322,G5323,G5324,G5325,G5326,G5327,G5328,G5329,G5330,G5331,G5332,G5333,G5334,G5335,G5336,G5337,G5338,G5339,G5340,
       G5341,G5342,G5343,G5344,G5345,G5346,G5347,G5348,G5349,G5350,G5351,G5352,G5353,G5354,G5355,G5356,G5357,G5358,G5359,G5360,
       G5361,G5362,G5363,G5364,G5365,G5366,G5367,G5368,G5369,G5370,G5371,G5372,G5373,G5374,G5375,G5376,G5377,G5378,G5379,G5380,
       G5381,G5382,G5383,G5384,G5385,G5386,G5387,G5388,G5389,G5390,G5391,G5392,G5393,G5394,G5395,G5396,G5397,G5398,G5399,G5400,
       G5401,G5402,G5403,G5404,G5405,G5406,G5407,G5408,G5409,G5410,G5411,G5412,G5413,G5414,G5415,G5416,G5417,G5418,G5419,G5420,
       G5421,G5422,G5423,G5424,G5425,G5426,G5427,G5428,G5429,G5430,G5431,G5432,G5433,G5434,G5435,G5436,G5437,G5438,G5439,G5440,
       G5441,G5442,G5443,G5444,G5445,G5446,G5447,G5448,G5449,G5450,G5451,G5452,G5453,G5454,G5455,G5456,G5457,G5458,G5459,G5460,
       G5461,G5462,G5463,G5464,G5465,G5466,G5467,G5468,G5469,G5470,G5471,G5472,G5473,G5474,G5475,G5476,G5477,G5478,G5479,G5480,
       G5481,G5482,G5483,G5484,G5485,G5486,G5487,G5488,G5489,G5490,G5491,G5492,G5493,G5494,G5495,G5496,G5497,G5498,G5499,G5500,
       G5501,G5502,G5503,G5504,G5505,G5506,G5507,G5508,G5509,G5510,G5511,G5512,G5513,G5514,G5515,G5516,G5517,G5518,G5519,G5520,
       G5521,G5522,G5523,G5524,G5525,G5526,G5527,G5528,G5529,G5530,G5531,G5532,G5533,G5534,G5535,G5536,G5537,G5538,G5539,G5540,
       G5541,G5542,G5543,G5544,G5545,G5546,G5547,G5548,G5549,G5550,G5551,G5552,G5553,G5554,G5555,G5556,G5557,G5558,G5559,G5560,
       G5561,G5562,G5563,G5564,G5565,G5566,G5567,G5568,G5569,G5570,G5571,G5572,G5573,G5574,G5575,G5576,G5577,G5578,G5579,G5580,
       G5581,G5582,G5583,G5584,G5585,G5586,G5587,G5588,G5589,G5590,G5591,G5592,G5593,G5594,G5595,G5596,G5597,G5598,G5599,G5600,
       G5601,G5602,G5603,G5604,G5605,G5606,G5607,G5608,G5609,G5610,G5611,G5612,G5613,G5614,G5615,G5616,G5617,G5618,G5619,G5620,
       G5621,G5622,G5623,G5624,G5625,G5626,G5627,G5628,G5629,G5630,G5631,G5632,G5633,G5634,G5635,G5636,G5637,G5638,G5639,G5640,
       G5641,G5642,G5643,G5644,G5645,G5646,G5647,G5648,G5649,G5650,G5651,G5652,G5653,G5654,G5655,G5656,G5657,G5658,G5659,G5660,
       G5661,G5662,G5663,G5664,G5665,G5666,G5667,G5668,G5669,G5670,G5671,G5672,G5673,G5674,G5675,G5676,G5677,G5678,G5679,G5680,
       G5681,G5682,G5683,G5684,G5685,G5686,G5687,G5688,G5689,G5690,G5691,G5692,G5693,G5694,G5695,G5696,G5697,G5698,G5699,G5700,
       G5701,G5702,G5703,G5704,G5705,G5706,G5707,G5708,G5709,G5710,G5711,G5712,G5713,G5714,G5715,G5716,G5717,G5718,G5719,G5720,
       G5721,G5722,G5723,G5724,G5725,G5726,G5727,G5728,G5729,G5730,G5731,G5732,G5733,G5734,G5735,G5736,G5737,G5738,G5739,G5740,
       G5741,G5742,G5743,G5744,G5745,G5746,G5747,G5748,G5749,G5750,G5751,G5752,G5753,G5754,G5755,G5756,G5757,G5758,G5759,G5760,
       G5761,G5762,G5763,G5764,G5765,G5766,G5767,G5768,G5769,G5770,G5771,G5772,G5773,G5774,G5775,G5776,G5777,G5778,G5779,G5780,
       G5781,G5782,G5783,G5784,G5785,G5786,G5787,G5788,G5789,G5790,G5791,G5792,G5793,G5794,G5795,G5796,G5797,G5798,G5799,G5800,
       G5801,G5802,G5803,G5804,G5805,G5806,G5807,G5808,G5809,G5810,G5811,G5812,G5813,G5814,G5815,G5816,G5817,G5818,G5819,G5820,
       G5821,G5822,G5823,G5824,G5825,G5826,G5827,G5828,G5829,G5830,G5831,G5832,G5833,G5834,G5835,G5836,G5837,G5838,G5839,G5840,
       G5841,G5842,G5843,G5844,G5845,G5846,G5847,G5848,G5849,G5850,G5851,G5852,G5853,G5854,G5855,G5856,G5857,G5858,G5859,G5860,
       G5861,G5862,G5863,G5864,G5865,G5866,G5867,G5868,G5869,G5870,G5871,G5872,G5873,G5874,G5875,G5876,G5877,G5878,G5879,G5880,
       G5881,G5882,G5883,G5884,G5885,G5886,G5887,G5888,G5889,G5890,G5891,G5892,G5893,G5894,G5895,G5896,G5897,G5898,G5899,G5900,
       G5901,G5902,G5903,G5904,G5905,G5906,G5907,G5908,G5909,G5910,G5911,G5912,G5913,G5914,G5915,G5916,G5917,G5918,G5919,G5920,
       G5921,G5922,G5923,G5924,G5925,G5926,G5927,G5928,G5929,G5930,G5931,G5932,G5933,G5934,G5935,G5936,G5937,G5938,G5939,G5940,
       G5941,G5942,G5943,G5944,G5945,G5946,G5947,G5948,G5949,G5950,G5951,G5952,G5953,G5954,G5955,G5956,G5957,G5958,G5959,G5960,
       G5961,G5962,G5963,G5964,G5965,G5966,G5967,G5968,G5969,G5970,G5971,G5972,G5973,G5974,G5975,G5976,G5977,G5978,G5979,G5980,
       G5981,G5982,G5983,G5984,G5985,G5986,G5987,G5988,G5989,G5990,G5991,G5992,G5993,G5994,G5995,G5996,G5997,G5998,G5999,G6000,
       G6001,G6002,G6003,G6004,G6005,G6006,G6007,G6008,G6009,G6010,G6011,G6012,G6013,G6014,G6015,G6016,G6017,G6018,G6019,G6020,
       G6021,G6022,G6023,G6024,G6025,G6026,G6027,G6028,G6029,G6030,G6031,G6032,G6033,G6034,G6035,G6036,G6037,G6038,G6039,G6040,
       G6041,G6042,G6043,G6044,G6045,G6046,G6047,G6048,G6049,G6050,G6051,G6052,G6053,G6054,G6055,G6056,G6057,G6058,G6059,G6060,
       G6061,G6062,G6063,G6064,G6065,G6066,G6067,G6068,G6069,G6070,G6071,G6072,G6073,G6074,G6075,G6076,G6077,G6078,G6079,G6080,
       G6081,G6082,G6083,G6084,G6085,G6086,G6087,G6088,G6089,G6090,G6091,G6092,G6093,G6094,G6095,G6096,G6097,G6098,G6099,G6100,
       G6101,G6102,G6103,G6104,G6105,G6106,G6107,G6108,G6109,G6110,G6111,G6112,G6113,G6114,G6115,G6116,G6117,G6118,G6119,G6120,
       G6121,G6122,G6123,G6124,G6125,G6126,G6127,G6128,G6129,G6130,G6131,G6132,G6133,G6134,G6135,G6136,G6137,G6138,G6139,G6140,
       G6141,G6142,G6143,G6144,G6145,G6146,G6147,G6148,G6149,G6150,G6151,G6152,G6153,G6154,G6155,G6156,G6157,G6158,G6159,G6160,
       G6161,G6162,G6163,G6164,G6165,G6166,G6167,G6168,G6169,G6170,G6171,G6172,G6173,G6174,G6175,G6176,G6177,G6178,G6179,G6180,
       G6181,G6182,G6183,G6184,G6185,G6186,G6187,G6188,G6189,G6190,G6191,G6192,G6193,G6194,G6195,G6196,G6197,G6198,G6199,G6200,
       G6201,G6202,G6203,G6204,G6205,G6206,G6207,G6208,G6209,G6210,G6211,G6212,G6213,G6214,G6215,G6216,G6217,G6218,G6219,G6220,
       G6221,G6222,G6223,G6224,G6225,G6226,G6227,G6228,G6229,G6230,G6231,G6232,G6233,G6234,G6235,G6236,G6237,G6238,G6239,G6240,
       G6241,G6242,G6243,G6244,G6245,G6246,G6247,G6248,G6249,G6250,G6251,G6252,G6253,G6254,G6255,G6256,G6257,G6258,G6259,G6260,
       G6261,G6262,G6263,G6264,G6265,G6266,G6267,G6268,G6269,G6270,G6271,G6272,G6273,G6274,G6275,G6276,G6277,G6278,G6279,G6280,
       G6281,G6282,G6283,G6284,G6285,G6286,G6287,G6288,G6289,G6290,G6291,G6292,G6293,G6294,G6295,G6296,G6297,G6298,G6299,G6300,
       G6301,G6302,G6303,G6304,G6305,G6306,G6307,G6308,G6309,G6310,G6311,G6312,G6313,G6314,G6315,G6316,G6317,G6318,G6319,G6320,
       G6321,G6322,G6323,G6324,G6325,G6326,G6327,G6328,G6329,G6330,G6331,G6332,G6333,G6334,G6335,G6336,G6337,G6338,G6339,G6340,
       G6341,G6342,G6343,G6344,G6345,G6346,G6347,G6348,G6349,G6350,G6351,G6352,G6353,G6354,G6355,G6356,G6357,G6358,G6359,G6360,
       G6361,G6362,G6363,G6364,G6365,G6366,G6367,G6368,G6369,G6370,G6371,G6372,G6373,G6374,G6375,G6376,G6377,G6378,G6379,G6380,
       G6381,G6382,G6383,G6384,G6385,G6386,G6387,G6388,G6389,G6390,G6391,G6392,G6393,G6394,G6395,G6396,G6397,G6398,G6399,G6400,
       G6401,G6402,G6403,G6404,G6405,G6406,G6407,G6408,G6409,G6410,G6411,G6412,G6413,G6414,G6415,G6416,G6417,G6418,G6419,G6420,
       G6421,G6422,G6423,G6424,G6425,G6426,G6427,G6428,G6429,G6430,G6431,G6432,G6433,G6434,G6435,G6436,G6437,G6438,G6439,G6440,
       G6441,G6442,G6443,G6444,G6445,G6446,G6447,G6448,G6449,G6450,G6451,G6452,G6453,G6454,G6455,G6456,G6457,G6458,G6459,G6460,
       G6461,G6462,G6463,G6464,G6465,G6466,G6467,G6468,G6469,G6470,G6471,G6472,G6473,G6474,G6475,G6476,G6477,G6478,G6479,G6480,
       G6481,G6482,G6483,G6484,G6485,G6486,G6487,G6488,G6489,G6490,G6491,G6492,G6493,G6494,G6495,G6496,G6497,G6498,G6499,G6500,
       G6501,G6502,G6503,G6504,G6505,G6506,G6507,G6508,G6509,G6510,G6511,G6512,G6513,G6514,G6515,G6516,G6517,G6518,G6519,G6520,
       G6521,G6522,G6523,G6524,G6525,G6526,G6527,G6528,G6529,G6530,G6531,G6532,G6533,G6534,G6535,G6536,G6537,G6538,G6539,G6540,
       G6541,G6542,G6543,G6544,G6545,G6546,G6547,G6548,G6549,G6550,G6551,G6552,G6553,G6554,G6555,G6556,G6557,G6558,G6559,G6560,
       G6561,G6562,G6563,G6564,G6565,G6566,G6567,G6568,G6569,G6570,G6571,G6572,G6573,G6574,G6575,G6576,G6577,G6578,G6579,G6580,
       G6581,G6582,G6583,G6584,G6585,G6586,G6587,G6588,G6589,G6590,G6591,G6592,G6593,G6594,G6595,G6596,G6597,G6598,G6599,G6600,
       G6601,G6602,G6603,G6604,G6605,G6606,G6607,G6608,G6609,G6610,G6611,G6612,G6613,G6614,G6615,G6616,G6617,G6618,G6619,G6620,
       G6621,G6622,G6623,G6624,G6625,G6626,G6627,G6628,G6629,G6630,G6631,G6632,G6633,G6634,G6635,G6636,G6637,G6638,G6639,G6640,
       G6641,G6642,G6643,G6644,G6645,G6646,G6647,G6648,G6649,G6650,G6651,G6652,G6653,G6654,G6655,G6656,G6657,G6658,G6659,G6660,
       G6661,G6662,G6663,G6664,G6665,G6666,G6667,G6668,G6669,G6670,G6671,G6672,G6673,G6674,G6675,G6676,G6677,G6678,G6679,G6680,
       G6681,G6682,G6683,G6684,G6685,G6686,G6687,G6688,G6689,G6690,G6691,G6692,G6693,G6694,G6695,G6696,G6697,G6698,G6699,G6700,
       G6701,G6702,G6703,G6704,G6705,G6706,G6707,G6708,G6709,G6710,G6711,G6712,G6713,G6714,G6715,G6716,G6717,G6718,G6719,G6720,
       G6721,G6722,G6723,G6724,G6725,G6726,G6727,G6728,G6729,G6730,G6731,G6732,G6733,G6734,G6735,G6736,G6737,G6738,G6739,G6740,
       G6741,G6742,G6743,G6744,G6745,G6746,G6747,G6748,G6749,G6750,G6751,G6752,G6753,G6754,G6755,G6756,G6757,G6758,G6759,G6760,
       G6761,G6762,G6763,G6764,G6765,G6766,G6767,G6768,G6769,G6770,G6771,G6772,G6773,G6774,G6775,G6776,G6777,G6778,G6779,G6780,
       G6781,G6782,G6783,G6784,G6785,G6786,G6787,G6788,G6789,G6790,G6791,G6792,G6793,G6794,G6795,G6796,G6797,G6798,G6799,G6800,
       G6801,G6802,G6803,G6804,G6805,G6806,G6807,G6808,G6809,G6810,G6811,G6812,G6813,G6814,G6815,G6816,G6817,G6818,G6819,G6820,
       G6821,G6822,G6823,G6824,G6825,G6826,G6827,G6828,G6829,G6830,G6831,G6832,G6833,G6834,G6835,G6836,G6837,G6838,G6839,G6840,
       G6841,G6842,G6843,G6844,G6845,G6846,G6847,G6848,G6849,G6850,G6851,G6852,G6853,G6854,G6855,G6856,G6857,G6858,G6859,G6860,
       G6861,G6862,G6863,G6864,G6865,G6866,G6867,G6868,G6869,G6870,G6871,G6872,G6873,G6874,G6875,G6876,G6877,G6878,G6879,G6880,
       G6881,G6882,G6883,G6884,G6885,G6886,G6887,G6888,G6889,G6890,G6891,G6892,G6893,G6894,G6895,G6896,G6897,G6898,G6899,G6900,
       G6901,G6902,G6903,G6904,G6905,G6906,G6907,G6908,G6909,G6910,G6911,G6912,G6913,G6914,G6915,G6916,G6917,G6918,G6919,G6920,
       G6921,G6922,G6923,G6924,G6925,G6926,G6927,G6928,G6929,G6930,G6931,G6932,G6933,G6934,G6935,G6936,G6937,G6938,G6939,G6940,
       G6941,G6942,G6943,G6944,G6945,G6946,G6947,G6948,G6949,G6950,G6951,G6952,G6953,G6954,G6955,G6956,G6957,G6958,G6959,G6960,
       G6961,G6962,G6963,G6964,G6965,G6966,G6967,G6968,G6969,G6970,G6971,G6972,G6973,G6974,G6975,G6976,G6977,G6978,G6979,G6980,
       G6981,G6982,G6983,G6984,G6985,G6986,G6987,G6988,G6989,G6990,G6991,G6992,G6993,G6994,G6995,G6996,G6997,G6998,G6999,G7000,
       G7001,G7002,G7003,G7004,G7005,G7006,G7007,G7008,G7009,G7010,G7011,G7012,G7013,G7014,G7015,G7016,G7017,G7018,G7019,G7020,
       G7021,G7022,G7023,G7024,G7025,G7026,G7027,G7028,G7029,G7030,G7031,G7032,G7033,G7034,G7035,G7036,G7037,G7038,G7039,G7040,
       G7041,G7042,G7043,G7044,G7045,G7046,G7047,G7048,G7049,G7050,G7051,G7052,G7053,G7054,G7055,G7056,G7057,G7058,G7059,G7060,
       G7061,G7062,G7063,G7064,G7065,G7066,G7067,G7068,G7069,G7070,G7071,G7072,G7073,G7074,G7075,G7076,G7077,G7078,G7079,G7080,
       G7081,G7082,G7083,G7084,G7085,G7086,G7087,G7088,G7089,G7090,G7091,G7092,G7093,G7094,G7095,G7096,G7097,G7098,G7099,G7100,
       G7101,G7102,G7103,G7104,G7105,G7106,G7107,G7108,G7109,G7110,G7111,G7112,G7113,G7114,G7115,G7116,G7117,G7118,G7119,G7120,
       G7121,G7122,G7123,G7124,G7125,G7126,G7127,G7128,G7129,G7130,G7131,G7132,G7133,G7134,G7135,G7136,G7137,G7138,G7139,G7140,
       G7141,G7142,G7143,G7144,G7145,G7146,G7147,G7148,G7149,G7150,G7151,G7152,G7153,G7154,G7155,G7156,G7157,G7158,G7159,G7160,
       G7161,G7162,G7163,G7164,G7165,G7166,G7167,G7168,G7169,G7170,G7171,G7172,G7173,G7174,G7175,G7176,G7177,G7178,G7179,G7180,
       G7181,G7182,G7183,G7184,G7185,G7186,G7187,G7188,G7189,G7190,G7191,G7192,G7193,G7194,G7195,G7196,G7197,G7198,G7199,G7200,
       G7201,G7202,G7203,G7204,G7205,G7206,G7207,G7208,G7209,G7210,G7211,G7212,G7213,G7214,G7215,G7216,G7217,G7218,G7219,G7220,
       G7221,G7222,G7223,G7224,G7225,G7226,G7227,G7228,G7229,G7230,G7231,G7232,G7233,G7234,G7235,G7236,G7237,G7238,G7239,G7240,
       G7241,G7242,G7243,G7244,G7245,G7246,G7247,G7248,G7249,G7250,G7251,G7252,G7253,G7254,G7255,G7256,G7257,G7258,G7259,G7260,
       G7261,G7262,G7263,G7264,G7265,G7266,G7267,G7268,G7269,G7270,G7271,G7272,G7273,G7274,G7275,G7276,G7277,G7278,G7279,G7280,
       G7281,G7282,G7283,G7284,G7285,G7286,G7287,G7288,G7289,G7290,G7291,G7292,G7293,G7294,G7295,G7296,G7297,G7298,G7299,G7300,
       G7301,G7302,G7303,G7304,G7305,G7306,G7307,G7308,G7309,G7310,G7311,G7312,G7313,G7314,G7315,G7316,G7317,G7318,G7319,G7320,
       G7321,G7322,G7323,G7324,G7325,G7326,G7327,G7328,G7329,G7330,G7331,G7332,G7333,G7334,G7335,G7336,G7337,G7338,G7339,G7340,
       G7341,G7342,G7343,G7344,G7345,G7346,G7347,G7348,G7349,G7350,G7351,G7352,G7353,G7354,G7355,G7356,G7357,G7358,G7359,G7360,
       G7361,G7362,G7363,G7364,G7365,G7366,G7367,G7368,G7369,G7370,G7371,G7372,G7373,G7374,G7375,G7376,G7377,G7378,G7379,G7380,
       G7381,G7382,G7383,G7384,G7385,G7386,G7387,G7388,G7389,G7390,G7391,G7392,G7393,G7394,G7395,G7396,G7397,G7398,G7399,G7400,
       G7401,G7402,G7403,G7404,G7405,G7406,G7407,G7408,G7409,G7410,G7411,G7412,G7413,G7414,G7415,G7416,G7417,G7418,G7419,G7420,
       G7421,G7422,G7423,G7424,G7425,G7426,G7427,G7428,G7429,G7430,G7431,G7432,G7433,G7434,G7435,G7436,G7437,G7438,G7439,G7440,
       G7441,G7442,G7443,G7444,G7445,G7446,G7447,G7448,G7449,G7450,G7451,G7452,G7453,G7454,G7455,G7456,G7457,G7458,G7459,G7460,
       G7461,G7462,G7463,G7464,G7465,G7466,G7467,G7468,G7469,G7470,G7471,G7472,G7473,G7474,G7475,G7476,G7477,G7478,G7479,G7480,
       G7481,G7482,G7483,G7484,G7485,G7486,G7487,G7488,G7489,G7490,G7491,G7492,G7493,G7494,G7495,G7496,G7497,G7498,G7499,G7500,
       G7501,G7502,G7503,G7504,G7505,G7506,G7507,G7508,G7509,G7510,G7511,G7512,G7513,G7514,G7515,G7516,G7517,G7518,G7519,G7520,
       G7521,G7522,G7523,G7524,G7525,G7526,G7527,G7528,G7529,G7530,G7531,G7532,G7533,G7534,G7535,G7536,G7537,G7538,G7539,G7540,
       G7541,G7542,G7543,G7544,G7545,G7546,G7547,G7548,G7549,G7550,G7551,G7552,G7553,G7554,G7555,G7556,G7557,G7558,G7559,G7560,
       G7561,G7562,G7563,G7564,G7565,G7566,G7567,G7568,G7569,G7570,G7571,G7572,G7573,G7574,G7575,G7576,G7577,G7578,G7579,G7580,
       G7581,G7582,G7583,G7584,G7585,G7586,G7587,G7588,G7589,G7590,G7591,G7592,G7593,G7594,G7595,G7596,G7597,G7598,G7599,G7600,
       G7601,G7602,G7603,G7604,G7605,G7606,G7607,G7608,G7609,G7610,G7611,G7612,G7613,G7614,G7615,G7616,G7617,G7618,G7619,G7620,
       G7621,G7622,G7623,G7624,G7625,G7626,G7627,G7628,G7629,G7630,G7631,G7632,G7633,G7634,G7635,G7636,G7637,G7638,G7639,G7640,
       G7641,G7642,G7643,G7644,G7645,G7646,G7647,G7648,G7649,G7650,G7651,G7652,G7653,G7654,G7655,G7656,G7657,G7658,G7659,G7660,
       G7661,G7662,G7663,G7664,G7665,G7666,G7667,G7668,G7669,G7670,G7671,G7672,G7673,G7674,G7675,G7676,G7677,G7678,G7679,G7680,
       G7681,G7682,G7683,G7684,G7685,G7686,G7687,G7688,G7689,G7690,G7691,G7692,G7693,G7694,G7695,G7696,G7697,G7698,G7699,G7700,
       G7701,G7702,G7703,G7704,G7705,G7706,G7707,G7708,G7709,G7710,G7711,G7712,G7713,G7714,G7715,G7716,G7717,G7718,G7719,G7720,
       G7721,G7722,G7723,G7724,G7725,G7726,G7727,G7728,G7729,G7730,G7731,G7732,G7733,G7734,G7735,G7736,G7737,G7738,G7739,G7740,
       G7741,G7742,G7743,G7744,G7745,G7746,G7747,G7748,G7749,G7750,G7751,G7752,G7753,G7754,G7755,G7756,G7757,G7758,G7759,G7760,
       G7761,G7762,G7763,G7764,G7765,G7766,G7767,G7768,G7769,G7770,G7771,G7772,G7773,G7774,G7775,G7776,G7777,G7778,G7779,G7780,
       G7781,G7782,G7783,G7784,G7785,G7786,G7787,G7788,G7789,G7790,G7791,G7792,G7793,G7794,G7795,G7796,G7797,G7798,G7799,G7800,
       G7801,G7802,G7803,G7804,G7805,G7806,G7807,G7808,G7809,G7810,G7811,G7812,G7813,G7814,G7815,G7816,G7817,G7818,G7819,G7820,
       G7821,G7822,G7823,G7824,G7825,G7826,G7827,G7828,G7829,G7830,G7831,G7832,G7833,G7834,G7835,G7836,G7837,G7838,G7839,G7840,
       G7841,G7842,G7843,G7844,G7845,G7846,G7847,G7848,G7849,G7850,G7851,G7852,G7853,G7854,G7855,G7856,G7857,G7858,G7859,G7860,
       G7861,G7862,G7863,G7864,G7865,G7866,G7867,G7868,G7869,G7870,G7871,G7872,G7873,G7874,G7875,G7876,G7877,G7878,G7879,G7880,
       G7881,G7882,G7883,G7884,G7885,G7886,G7887,G7888,G7889,G7890,G7891,G7892,G7893,G7894,G7895,G7896,G7897,G7898,G7899,G7900,
       G7901,G7902,G7903,G7904,G7905,G7906,G7907,G7908,G7909,G7910,G7911,G7912,G7913,G7914,G7915,G7916,G7917,G7918,G7919,G7920,
       G7921,G7922,G7923,G7924,G7925,G7926,G7927,G7928,G7929,G7930,G7931,G7932,G7933,G7934,G7935,G7936,G7937,G7938,G7939,G7940,
       G7941,G7942,G7943,G7944,G7945,G7946,G7947,G7948,G7949,G7950,G7951,G7952,G7953,G7954,G7955,G7956,G7957,G7958,G7959,G7960,
       G7961,G7962,G7963,G7964,G7965,G7966,G7967,G7968,G7969,G7970,G7971,G7972,G7973,G7974,G7975,G7976,G7977,G7978,G7979,G7980,
       G7981,G7982,G7983,G7984,G7985,G7986,G7987,G7988,G7989,G7990,G7991,G7992,G7993,G7994,G7995,G7996,G7997,G7998,G7999,G8000,
       G8001,G8002,G8003,G8004,G8005,G8006,G8007,G8008,G8009,G8010,G8011,G8012,G8013,G8014,G8015,G8016,G8017,G8018,G8019,G8020,
       G8021,G8022,G8023,G8024,G8025,G8026,G8027,G8028,G8029,G8030,G8031,G8032,G8033,G8034,G8035,G8036,G8037,G8038,G8039,G8040,
       G8041,G8042,G8043,G8044,G8045,G8046,G8047,G8048,G8049,G8050,G8051,G8052,G8053,G8054,G8055,G8056,G8057,G8058,G8059,G8060,
       G8061,G8062,G8063,G8064,G8065,G8066,G8067,G8068,G8069,G8070,G8071,G8072,G8073,G8074,G8075,G8076,G8077,G8078,G8079,G8080,
       G8081,G8082,G8083,G8084,G8085,G8086,G8087,G8088,G8089,G8090,G8091,G8092,G8093,G8094,G8095,G8096,G8097,G8098,G8099,G8100,
       G8101,G8102,G8103,G8104,G8105,G8106,G8107,G8108,G8109,G8110,G8111,G8112,G8113,G8114,G8115,G8116,G8117,G8118,G8119,G8120,
       G8121,G8122,G8123,G8124,G8125,G8126,G8127,G8128,G8129,G8130,G8131,G8132,G8133,G8134,G8135,G8136,G8137,G8138,G8139,G8140,
       G8141,G8142,G8143,G8144,G8145,G8146,G8147,G8148,G8149,G8150,G8151,G8152,G8153,G8154,G8155,G8156,G8157,G8158,G8159,G8160,
       G8161,G8162,G8163,G8164,G8165,G8166,G8167,G8168,G8169,G8170,G8171,G8172,G8173,G8174,G8175,G8176,G8177,G8178,G8179,G8180,
       G8181,G8182,G8183,G8184,G8185,G8186,G8187,G8188,G8189,G8190,G8191,G8192,G8193,G8194,G8195,G8196,G8197,G8198,G8199,G8200,
       G8201,G8202,G8203,G8204,G8205,G8206,G8207,G8208,G8209,G8210,G8211,G8212,G8213,G8214,G8215,G8216,G8217,G8218,G8219,G8220,
       G8221,G8222,G8223,G8224,G8225,G8226,G8227,G8228,G8229,G8230,G8231,G8232,G8233,G8234,G8235,G8236,G8237,G8238,G8239,G8240,
       G8241,G8242,G8243,G8244,G8245,G8246,G8247,G8248,G8249,G8250,G8251,G8252,G8253,G8254,G8255,G8256,G8257,G8258,G8259,G8260,
       G8261,G8262,G8263,G8264,G8265,G8266,G8267,G8268,G8269,G8270,G8271,G8272,G8273,G8274,G8275,G8276,G8277,G8278,G8279,G8280,
       G8281,G8282,G8283,G8284,G8285,G8286,G8287,G8288,G8289,G8290,G8291,G8292,G8293,G8294,G8295,G8296,G8297,G8298,G8299,G8300,
       G8301,G8302,G8303,G8304,G8305,G8306,G8307,G8308,G8309,G8310,G8311,G8312,G8313,G8314,G8315,G8316,G8317,G8318,G8319,G8320,
       G8321,G8322,G8323,G8324,G8325,G8326,G8327,G8328,G8329,G8330,G8331,G8332,G8333,G8334,G8335,G8336,G8337,G8338,G8339,G8340,
       G8341,G8342,G8343,G8344,G8345,G8346,G8347,G8348,G8349,G8350,G8351,G8352,G8353,G8354,G8355,G8356,G8357,G8358,G8359,G8360,
       G8361,G8362,G8363,G8364,G8365,G8366,G8367,G8368,G8369,G8370,G8371,G8372,G8373,G8374,G8375,G8376,G8377,G8378,G8379,G8380,
       G8381,G8382,G8383,G8384,G8385,G8386,G8387,G8388,G8389,G8390,G8391,G8392,G8393,G8394,G8395,G8396,G8397,G8398,G8399,G8400,
       G8401,G8402,G8403,G8404,G8405,G8406,G8407,G8408,G8409,G8410,G8411,G8412,G8413,G8414,G8415,G8416,G8417,G8418,G8419,G8420,
       G8421,G8422,G8423,G8424,G8425,G8426,G8427,G8428,G8429,G8430,G8431,G8432,G8433,G8434,G8435,G8436,G8437,G8438,G8439,G8440,
       G8441,G8442,G8443,G8444,G8445,G8446,G8447,G8448,G8449,G8450,G8451,G8452,G8453,G8454,G8455,G8456,G8457,G8458,G8459,G8460,
       G8461,G8462,G8463,G8464,G8465,G8466,G8467,G8468,G8469,G8470,G8471,G8472,G8473,G8474,G8475,G8476,G8477,G8478,G8479,G8480,
       G8481,G8482,G8483,G8484,G8485,G8486,G8487,G8488,G8489,G8490,G8491,G8492,G8493,G8494,G8495,G8496,G8497,G8498,G8499,G8500,
       G8501,G8502,G8503,G8504,G8505,G8506,G8507,G8508,G8509,G8510,G8511,G8512,G8513,G8514,G8515,G8516,G8517,G8518,G8519,G8520,
       G8521,G8522,G8523,G8524,G8525,G8526,G8527,G8528,G8529,G8530,G8531,G8532,G8533,G8534,G8535,G8536,G8537,G8538,G8539,G8540,
       G8541,G8542,G8543,G8544,G8545,G8546,G8547,G8548,G8549,G8550,G8551,G8552,G8553,G8554,G8555,G8556,G8557,G8558,G8559,G8560,
       G8561,G8562,G8563,G8564,G8565,G8566,G8567,G8568,G8569,G8570,G8571,G8572,G8573,G8574,G8575,G8576,G8577,G8578,G8579,G8580,
       G8581,G8582,G8583,G8584,G8585,G8586,G8587,G8588,G8589,G8590,G8591,G8592,G8593,G8594,G8595,G8596,G8597,G8598,G8599,G8600,
       G8601,G8602,G8603,G8604,G8605,G8606,G8607,G8608,G8609,G8610,G8611,G8612,G8613,G8614,G8615,G8616,G8617,G8618,G8619,G8620,
       G8621,G8622,G8623,G8624,G8625,G8626,G8627,G8628,G8629,G8630,G8631,G8632,G8633,G8634,G8635,G8636,G8637,G8638,G8639,G8640,
       G8641,G8642,G8643,G8644,G8645,G8646,G8647,G8648,G8649,G8650,G8651,G8652,G8653,G8654,G8655,G8656,G8657,G8658,G8659,G8660,
       G8661,G8662,G8663,G8664,G8665,G8666,G8667,G8668,G8669,G8670,G8671,G8672,G8673,G8674,G8675,G8676,G8677,G8678,G8679,G8680,
       G8681,G8682,G8683,G8684,G8685,G8686,G8687,G8688,G8689,G8690,G8691,G8692,G8693,G8694,G8695,G8696,G8697,G8698,G8699,G8700,
       G8701,G8702,G8703,G8704,G8705,G8706,G8707,G8708,G8709,G8710,G8711,G8712,G8713,G8714,G8715,G8716,G8717,G8718,G8719,G8720,
       G8721,G8722,G8723,G8724,G8725,G8726,G8727,G8728,G8729,G8730,G8731,G8732,G8733,G8734,G8735,G8736,G8737,G8738,G8739,G8740,
       G8741,G8742,G8743,G8744,G8745,G8746,G8747,G8748,G8749,G8750,G8751,G8752,G8753,G8754,G8755,G8756,G8757,G8758,G8759,G8760,
       G8761,G8762,G8763,G8764,G8765,G8766,G8767,G8768,G8769,G8770,G8771,G8772,G8773,G8774,G8775,G8776,G8777,G8778,G8779,G8780,
       G8781,G8782,G8783,G8784,G8785,G8786,G8787,G8788,G8789,G8790,G8791,G8792,G8793,G8794,G8795,G8796,G8797,G8798,G8799,G8800,
       G8801,G8802,G8803,G8804,G8805,G8806,G8807,G8808,G8809,G8810,G8811,G8812,G8813,G8814,G8815,G8816,G8817,G8818,G8819,G8820,
       G8821,G8822,G8823,G8824,G8825,G8826,G8827,G8828,G8829,G8830,G8831,G8832,G8833,G8834,G8835,G8836,G8837,G8838,G8839,G8840,
       G8841,G8842,G8843,G8844,G8845,G8846,G8847,G8848,G8849,G8850,G8851,G8852,G8853,G8854,G8855,G8856,G8857,G8858,G8859,G8860,
       G8861,G8862,G8863,G8864,G8865,G8866,G8867,G8868,G8869,G8870,G8871,G8872,G8873,G8874,G8875,G8876,G8877,G8878,G8879,G8880,
       G8881,G8882,G8883,G8884,G8885,G8886,G8887,G8888,G8889,G8890,G8891,G8892,G8893,G8894,G8895,G8896,G8897,G8898,G8899,G8900,
       G8901,G8902,G8903,G8904,G8905,G8906,G8907,G8908,G8909,G8910,G8911,G8912,G8913,G8914,G8915,G8916,G8917,G8918,G8919,G8920,
       G8921,G8922,G8923,G8924,G8925,G8926,G8927,G8928,G8929,G8930,G8931,G8932,G8933,G8934,G8935,G8936,G8937,G8938,G8939,G8940,
       G8941,G8942,G8943,G8944,G8945,G8946,G8947,G8948,G8949,G8950,G8951,G8952,G8953,G8954,G8955,G8956,G8957,G8958,G8959,G8960,
       G8961,G8962,G8963,G8964,G8965,G8966,G8967,G8968,G8969,G8970,G8971,G8972,G8973,G8974,G8975,G8976,G8977,G8978,G8979,G8980,
       G8981,G8982,G8983,G8984,G8985,G8986,G8987,G8988,G8989,G8990,G8991,G8992,G8993,G8994,G8995,G8996,G8997,G8998,G8999,G9000,
       G9001,G9002,G9003,G9004,G9005,G9006,G9007,G9008,G9009,G9010,G9011,G9012,G9013,G9014,G9015,G9016,G9017,G9018,G9019,G9020,
       G9021,G9022,G9023,G9024,G9025,G9026,G9027,G9028,G9029,G9030,G9031,G9032,G9033,G9034,G9035,G9036,G9037,G9038,G9039,G9040,
       G9041,G9042,G9043,G9044,G9045,G9046,G9047,G9048,G9049,G9050,G9051,G9052,G9053,G9054,G9055,G9056,G9057,G9058,G9059,G9060,
       G9061,G9062,G9063,G9064,G9065,G9066,G9067,G9068,G9069,G9070,G9071,G9072,G9073,G9074,G9075,G9076,G9077,G9078,G9079,G9080,
       G9081,G9082,G9083,G9084,G9085,G9086,G9087,G9088,G9089,G9090,G9091,G9092,G9093,G9094,G9095,G9096,G9097,G9098,G9099,G9100,
       G9101,G9102,G9103,G9104,G9105,G9106,G9107,G9108,G9109,G9110,G9111,G9112,G9113,G9114,G9115,G9116,G9117,G9118,G9119,G9120,
       G9121,G9122,G9123,G9124,G9125,G9126,G9127,G9128,G9129,G9130,G9131,G9132,G9133,G9134,G9135,G9136,G9137,G9138,G9139,G9140,
       G9141,G9142,G9143,G9144,G9145,G9146,G9147,G9148,G9149,G9150,G9151,G9152,G9153,G9154,G9155,G9156,G9157,G9158,G9159,G9160,
       G9161,G9162,G9163,G9164,G9165,G9166,G9167,G9168,G9169,G9170,G9171,G9172,G9173,G9174,G9175,G9176,G9177,G9178,G9179,G9180,
       G9181,G9182,G9183,G9184,G9185,G9186,G9187,G9188,G9189,G9190,G9191,G9192,G9193,G9194,G9195,G9196,G9197,G9198,G9199,G9200,
       G9201,G9202,G9203,G9204,G9205,G9206,G9207,G9208,G9209,G9210,G9211,G9212,G9213,G9214,G9215,G9216,G9217,G9218,G9219,G9220,
       G9221,G9222,G9223,G9224,G9225,G9226,G9227,G9228,G9229,G9230,G9231,G9232,G9233,G9234,G9235,G9236,G9237,G9238,G9239,G9240,
       G9241,G9242,G9243,G9244,G9245,G9246,G9247,G9248,G9249,G9250,G9251,G9252,G9253,G9254,G9255,G9256,G9257,G9258,G9259,G9260,
       G9261,G9262,G9263,G9264,G9265,G9266,G9267,G9268,G9269,G9270,G9271,G9272,G9273,G9274,G9275,G9276,G9277,G9278,G9279,G9280,
       G9281,G9282,G9283,G9284,G9285,G9286,G9287,G9288,G9289,G9290,G9291,G9292,G9293,G9294,G9295,G9296,G9297,G9298,G9299,G9300,
       G9301,G9302,G9303,G9304,G9305,G9306,G9307,G9308,G9309,G9310,G9311,G9312,G9313,G9314,G9315,G9316,G9317,G9318,G9319,G9320,
       G9321,G9322,G9323,G9324,G9325,G9326,G9327,G9328,G9329,G9330,G9331,G9332,G9333,G9334,G9335,G9336,G9337,G9338,G9339,G9340,
       G9341,G9342,G9343,G9344,G9345,G9346,G9347,G9348,G9349,G9350,G9351,G9352,G9353,G9354,G9355,G9356,G9357,G9358,G9359,G9360,
       G9361,G9362,G9363,G9364,G9365,G9366,G9367,G9368,G9369,G9370,G9371,G9372,G9373,G9374,G9375,G9376,G9377,G9378,G9379,G9380,
       G9381,G9382,G9383,G9384,G9385,G9386,G9387,G9388,G9389,G9390,G9391,G9392,G9393,G9394,G9395,G9396,G9397,G9398,G9399,G9400,
       G9401,G9402,G9403,G9404,G9405,G9406,G9407,G9408,G9409,G9410,G9411,G9412,G9413,G9414,G9415,G9416,G9417,G9418,G9419,G9420,
       G9421,G9422,G9423,G9424,G9425,G9426,G9427,G9428,G9429,G9430,G9431,G9432,G9433,G9434,G9435,G9436,G9437,G9438,G9439,G9440,
       G9441,G9442,G9443,G9444,G9445,G9446,G9447,G9448,G9449,G9450,G9451,G9452,G9453,G9454,G9455,G9456,G9457,G9458,G9459,G9460,
       G9461,G9462,G9463,G9464,G9465,G9466,G9467,G9468,G9469,G9470,G9471,G9472,G9473,G9474,G9475,G9476,G9477,G9478,G9479,G9480,
       G9481,G9482,G9483,G9484,G9485,G9486,G9487,G9488,G9489,G9490,G9491,G9492,G9493,G9494,G9495,G9496,G9497,G9498,G9499,G9500,
       G9501,G9502,G9503,G9504,G9505,G9506,G9507,G9508,G9509,G9510,G9511,G9512,G9513,G9514,G9515,G9516,G9517,G9518,G9519,G9520,
       G9521,G9522,G9523,G9524,G9525,G9526,G9527,G9528,G9529,G9530,G9531,G9532,G9533,G9534,G9535,G9536,G9537,G9538,G9539,G9540,
       G9541,G9542,G9543,G9544,G9545,G9546,G9547,G9548,G9549,G9550,G9551,G9552,G9553,G9554,G9555,G9556,G9557,G9558,G9559,G9560,
       G9561,G9562,G9563,G9564,G9565,G9566,G9567,G9568,G9569,G9570,G9571,G9572,G9573,G9574,G9575,G9576,G9577,G9578,G9579,G9580,
       G9581,G9582,G9583,G9584,G9585,G9586,G9587,G9588,G9589,G9590,G9591,G9592,G9593,G9594,G9595,G9596,G9597,G9598,G9599,G9600,
       G9601,G9602,G9603,G9604,G9605,G9606,G9607,G9608,G9609,G9610,G9611,G9612,G9613,G9614,G9615,G9616,G9617,G9618,G9619,G9620,
       G9621,G9622,G9623,G9624,G9625,G9626,G9627,G9628,G9629,G9630,G9631,G9632,G9633,G9634,G9635,G9636,G9637,G9638,G9639,G9640,
       G9641,G9642,G9643,G9644,G9645,G9646,G9647,G9648,G9649,G9650,G9651,G9652,G9653,G9654,G9655,G9656,G9657,G9658,G9659,G9660,
       G9661,G9662,G9663,G9664,G9665,G9666,G9667,G9668,G9669,G9670,G9671,G9672,G9673,G9674,G9675,G9676,G9677,G9678,G9679,G9680,
       G9681,G9682,G9683,G9684,G9685,G9686,G9687,G9688,G9689,G9690,G9691,G9692,G9693,G9694,G9695,G9696,G9697,G9698,G9699,G9700,
       G9701,G9702,G9703,G9704,G9705,G9706,G9707,G9708,G9709,G9710,G9711,G9712,G9713,G9714,G9715,G9716,G9717,G9718,G9719,G9720,
       G9721,G9722,G9723,G9724,G9725,G9726,G9727,G9728,G9729,G9730,G9731,G9732,G9733,G9734,G9735,G9736,G9737,G9738,G9739,G9740,
       G9741,G9742,G9743,G9744,G9745,G9746,G9747,G9748,G9749,G9750,G9751,G9752,G9753,G9754,G9755,G9756,G9757,G9758,G9759,G9760,
       G9761,G9762,G9763,G9764,G9765,G9766,G9767,G9768,G9769,G9770,G9771,G9772,G9773,G9774,G9775,G9776,G9777,G9778,G9779,G9780,
       G9781,G9782,G9783,G9784,G9785,G9786,G9787,G9788,G9789,G9790,G9791,G9792,G9793,G9794,G9795,G9796,G9797,G9798,G9799,G9800,
       G9801,G9802,G9803,G9804,G9805,G9806,G9807,G9808,G9809,G9810,G9811,G9812,G9813,G9814,G9815,G9816,G9817,G9818,G9819,G9820,
       G9821,G9822,G9823,G9824,G9825,G9826,G9827,G9828,G9829,G9830,G9831,G9832,G9833,G9834,G9835,G9836,G9837,G9838,G9839,G9840,
       G9841,G9842,G9843,G9844,G9845,G9846,G9847,G9848,G9849,G9850,G9851,G9852,G9853,G9854,G9855,G9856,G9857,G9858,G9859,G9860,
       G9861,G9862,G9863,G9864,G9865,G9866,G9867,G9868,G9869,G9870,G9871,G9872,G9873,G9874,G9875,G9876,G9877,G9878,G9879,G9880,
       G9881,G9882,G9883,G9884,G9885,G9886,G9887,G9888,G9889,G9890,G9891,G9892,G9893,G9894,G9895,G9896,G9897,G9898,G9899,G9900,
       G9901,G9902,G9903,G9904,G9905,G9906,G9907,G9908,G9909,G9910,G9911,G9912,G9913,G9914,G9915,G9916,G9917,G9918,G9919,G9920,
       G9921,G9922,G9923,G9924,G9925,G9926,G9927,G9928,G9929,G9930,G9931,G9932,G9933,G9934,G9935,G9936,G9937,G9938,G9939,G9940,
       G9941,G9942,G9943,G9944,G9945,G9946,G9947,G9948,G9949,G9950,G9951,G9952,G9953,G9954,G9955,G9956,G9957,G9958,G9959,G9960,
       G9961,G9962,G9963,G9964,G9965,G9966,G9967,G9968,G9969,G9970,G9971,G9972,G9973,G9974,G9975,G9976,G9977,G9978,G9979,G9980,
       G9981,G9982,G9983,G9984,G9985,G9986,G9987,G9988,G9989,G9990,G9991,G9992,G9993,G9994,G9995,G9996,G9997,G9998,G9999,G10000,
       G10001,G10002,G10003,G10004,G10005,G10006,G10007,G10008,G10009,G10010,G10011,G10012,G10013,G10014,G10015,G10016,G10017,G10018,G10019,G10020,
       G10021,G10022,G10023,G10024,G10025,G10026,G10027,G10028,G10029,G10030,G10031,G10032,G10033,G10034,G10035,G10036,G10037,G10038,G10039,G10040,
       G10041,G10042,G10043,G10044,G10045,G10046,G10047,G10048,G10049,G10050,G10051,G10052,G10053,G10054,G10055,G10056,G10057,G10058,G10059,G10060,
       G10061,G10062,G10063,G10064,G10065,G10066,G10067,G10068,G10069,G10070,G10071,G10072,G10073,G10074,G10075,G10076,G10077,G10078,G10079,G10080,
       G10081,G10082,G10083,G10084,G10085,G10086,G10087,G10088,G10089,G10090,G10091,G10092,G10093,G10094,G10095,G10096,G10097,G10098,G10099,G10100,
       G10101,G10102,G10103,G10104,G10105,G10106,G10107,G10108,G10109,G10110,G10111,G10112,G10113,G10114,G10115,G10116,G10117,G10118,G10119,G10120,
       G10121,G10122,G10123,G10124,G10125,G10126,G10127,G10128,G10129,G10130,G10131,G10132,G10133,G10134,G10135,G10136,G10137,G10138,G10139,G10140,
       G10141,G10142,G10143,G10144,G10145,G10146,G10147,G10148,G10149,G10150,G10151,G10152,G10153,G10154,G10155,G10156,G10157,G10158,G10159,G10160,
       G10161,G10162,G10163,G10164,G10165,G10166,G10167,G10168,G10169,G10170,G10171,G10172,G10173,G10174,G10175,G10176,G10177,G10178,G10179,G10180,
       G10181,G10182,G10183,G10184,G10185,G10186,G10187,G10188,G10189,G10190,G10191,G10192,G10193,G10194,G10195,G10196,G10197,G10198,G10199,G10200,
       G10201,G10202,G10203,G10204,G10205,G10206,G10207,G10208,G10209,G10210,G10211,G10212,G10213,G10214,G10215,G10216,G10217,G10218,G10219,G10220,
       G10221,G10222,G10223,G10224,G10225,G10226,G10227,G10228,G10229,G10230,G10231,G10232,G10233,G10234,G10235,G10236,G10237,G10238,G10239,G10240,
       G10241,G10242,G10243,G10244,G10245,G10246,G10247,G10248,G10249,G10250,G10251,G10252,G10253,G10254,G10255,G10256,G10257,G10258,G10259,G10260,
       G10261,G10262,G10263,G10264,G10265,G10266,G10267,G10268,G10269,G10270,G10271,G10272,G10273,G10274,G10275,G10276,G10277,G10278,G10279,G10280,
       G10281,G10282,G10283,G10284,G10285,G10286,G10287,G10288,G10289,G10290,G10291,G10292,G10293,G10294,G10295,G10296,G10297,G10298,G10299,G10300,
       G10301,G10302,G10303,G10304,G10305,G10306,G10307,G10308,G10309,G10310,G10311,G10312,G10313,G10314,G10315,G10316,G10317,G10318,G10319,G10320,
       G10321,G10322,G10323,G10324,G10325,G10326,G10327,G10328,G10329,G10330,G10331,G10332,G10333,G10334,G10335,G10336,G10337,G10338,G10339,G10340,
       G10341,G10342,G10343,G10344,G10345,G10346,G10347,G10348,G10349,G10350,G10351,G10352,G10353,G10354,G10355,G10356,G10357,G10358,G10359,G10360,
       G10361,G10362,G10363,G10364,G10365,G10366,G10367,G10368,G10369,G10370,G10371,G10372,G10373,G10374,G10375,G10376,G10377,G10378,G10379,G10380,
       G10381,G10382,G10383,G10384,G10385,G10386,G10387,G10388,G10389,G10390,G10391,G10392,G10393,G10394,G10395,G10396,G10397,G10398,G10399,G10400,
       G10401,G10402,G10403,G10404,G10405,G10406,G10407,G10408,G10409,G10410,G10411,G10412,G10413,G10414,G10415,G10416,G10417,G10418,G10419,G10420,
       G10421,G10422,G10423,G10424,G10425,G10426,G10427,G10428,G10429,G10430,G10431,G10432,G10433,G10434,G10435,G10436,G10437,G10438,G10439,G10440,
       G10441,G10442,G10443,G10444,G10445,G10446,G10447,G10448,G10449,G10450,G10451,G10452,G10453,G10454,G10455,G10456,G10457,G10458,G10459,G10460,
       G10461,G10462,G10463,G10464,G10465,G10466,G10467,G10468,G10469,G10470,G10471,G10472,G10473,G10474,G10475,G10476,G10477,G10478,G10479,G10480,
       G10481,G10482,G10483,G10484,G10485,G10486,G10487,G10488,G10489,G10490,G10491,G10492,G10493,G10494,G10495,G10496,G10497,G10498,G10499,G10500,
       G10501,G10502,G10503,G10504,G10505,G10506,G10507,G10508,G10509,G10510,G10511,G10512,G10513,G10514,G10515,G10516,G10517,G10518,G10519,G10520,
       G10521,G10522,G10523,G10524,G10525,G10526,G10527,G10528,G10529,G10530,G10531,G10532,G10533,G10534,G10535,G10536,G10537,G10538,G10539,G10540,
       G10541,G10542,G10543,G10544,G10545,G10546,G10547,G10548,G10549,G10550,G10551,G10552,G10553,G10554,G10555,G10556,G10557,G10558,G10559,G10560,
       G10561,G10562,G10563,G10564,G10565,G10566,G10567,G10568,G10569,G10570,G10571,G10572,G10573,G10574,G10575,G10576,G10577,G10578,G10579,G10580,
       G10581,G10582,G10583,G10584,G10585,G10586,G10587,G10588,G10589,G10590,G10591,G10592,G10593,G10594,G10595,G10596,G10597,G10598,G10599,G10600,
       G10601,G10602,G10603,G10604,G10605,G10606,G10607,G10608,G10609,G10610,G10611,G10612,G10613,G10614,G10615,G10616,G10617,G10618,G10619,G10620,
       G10621,G10622,G10623,G10624,G10625,G10626,G10627,G10628,G10629,G10630,G10631,G10632,G10633,G10634,G10635,G10636,G10637,G10638,G10639,G10640,
       G10641,G10642,G10643,G10644,G10645,G10646,G10647,G10648,G10649,G10650,G10651,G10652,G10653,G10654,G10655,G10656,G10657,G10658,G10659,G10660,
       G10661,G10662,G10663,G10664,G10665,G10666,G10667,G10668,G10669,G10670,G10671,G10672,G10673,G10674,G10675,G10676,G10677,G10678,G10679,G10680,
       G10681,G10682,G10683,G10684,G10685,G10686,G10687,G10688,G10689,G10690,G10691,G10692,G10693,G10694,G10695,G10696,G10697,G10698,G10699,G10700,
       G10701,G10702,G10703,G10704,G10705,G10706,G10707,G10708,G10709,G10710,G10711,G10712,G10713,G10714,G10715,G10716,G10717,G10718,G10719,G10720,
       G10721,G10722,G10723,G10724,G10725,G10726,G10727,G10728,G10729,G10730,G10731,G10732,G10733,G10734,G10735,G10736,G10737,G10738,G10739,G10740,
       G10741,G10742,G10743,G10744,G10745,G10746,G10747,G10748,G10749,G10750,G10751,G10752,G10753,G10754,G10755,G10756,G10757,G10758,G10759,G10760,
       G10761,G10762,G10763,G10764,G10765,G10766,G10767,G10768,G10769,G10770,G10771,G10772,G10773,G10774,G10775,G10776,G10777,G10778,G10779,G10780,
       G10781,G10782,G10783,G10784,G10785,G10786,G10787,G10788,G10789,G10790,G10791,G10792,G10793,G10794,G10795,G10796,G10797,G10798,G10799,G10800,
       G10801,G10802,G10803,G10804,G10805,G10806,G10807,G10808,G10809,G10810,G10811,G10812,G10813,G10814,G10815,G10816,G10817,G10818,G10819,G10820,
       G10821,G10822,G10823,G10824,G10825,G10826,G10827,G10828,G10829,G10830,G10831,G10832,G10833,G10834,G10835,G10836,G10837,G10838,G10839,G10840,
       G10841,G10842,G10843,G10844,G10845,G10846,G10847,G10848,G10849,G10850,G10851,G10852,G10853,G10854,G10855,G10856,G10857,G10858,G10859,G10860,
       G10861,G10862,G10863,G10864,G10865,G10866,G10867,G10868,G10869,G10870,G10871,G10872,G10873,G10874,G10875,G10876,G10877,G10878,G10879,G10880,
       G10881,G10882,G10883,G10884,G10885,G10886,G10887,G10888,G10889,G10890,G10891,G10892,G10893,G10894,G10895,G10896,G10897,G10898,G10899,G10900,
       G10901,G10902,G10903,G10904,G10905,G10906,G10907,G10908,G10909,G10910,G10911,G10912,G10913,G10914,G10915,G10916,G10917,G10918,G10919,G10920,
       G10921,G10922,G10923,G10924,G10925,G10926,G10927,G10928,G10929,G10930,G10931,G10932,G10933,G10934,G10935,G10936,G10937,G10938,G10939,G10940,
       G10941,G10942,G10943,G10944,G10945,G10946,G10947,G10948,G10949,G10950,G10951,G10952,G10953,G10954,G10955,G10956,G10957,G10958,G10959,G10960,
       G10961,G10962,G10963,G10964,G10965,G10966,G10967,G10968,G10969,G10970,G10971,G10972,G10973,G10974,G10975,G10976,G10977,G10978,G10979,G10980,
       G10981,G10982,G10983,G10984,G10985,G10986,G10987,G10988,G10989,G10990,G10991,G10992,G10993,G10994,G10995,G10996,G10997,G10998,G10999,G11000,
       G11001,G11002,G11003,G11004,G11005,G11006,G11007,G11008,G11009,G11010,G11011,G11012,G11013,G11014,G11015,G11016,G11017,G11018,G11019,G11020,
       G11021,G11022,G11023,G11024,G11025,G11026,G11027,G11028,G11029,G11030,G11031,G11032,G11033,G11034,G11035,G11036,G11037,G11038,G11039,G11040,
       G11041,G11042,G11043,G11044,G11045,G11046,G11047,G11048,G11049,G11050,G11051,G11052,G11053,G11054,G11055,G11056,G11057,G11058,G11059,G11060,
       G11061,G11062,G11063,G11064,G11065,G11066,G11067,G11068,G11069,G11070,G11071,G11072,G11073,G11074,G11075,G11076,G11077,G11078,G11079,G11080,
       G11081,G11082,G11083,G11084,G11085,G11086,G11087,G11088,G11089,G11090,G11091,G11092,G11093,G11094,G11095,G11096,G11097,G11098,G11099,G11100,
       G11101,G11102,G11103,G11104,G11105,G11106,G11107,G11108,G11109,G11110,G11111,G11112,G11113,G11114,G11115,G11116,G11117,G11118,G11119,G11120,
       G11121,G11122,G11123,G11124,G11125,G11126,G11127,G11128,G11129,G11130,G11131,G11132,G11133,G11134,G11135,G11136,G11137,G11138,G11139,G11140,
       G11141,G11142,G11143,G11144,G11145,G11146,G11147,G11148,G11149,G11150,G11151,G11152,G11153,G11154,G11155,G11156,G11157,G11158,G11159,G11160,
       G11161,G11162,G11163,G11164,G11165,G11166,G11167,G11168,G11169,G11170,G11171,G11172,G11173,G11174,G11175,G11176,G11177,G11178,G11179,G11180,
       G11181,G11182,G11183,G11184,G11185,G11186,G11187,G11188,G11189,G11190,G11191,G11192,G11193,G11194,G11195,G11196,G11197,G11198,G11199,G11200,
       G11201,G11202,G11203,G11204,G11205,G11206,G11207,G11208,G11209,G11210,G11211,G11212,G11213,G11214,G11215,G11216,G11217,G11218,G11219,G11220,
       G11221,G11222,G11223,G11224,G11225,G11226,G11227,G11228,G11229,G11230,G11231,G11232,G11233,G11234,G11235,G11236,G11237,G11238,G11239,G11240,
       G11241,G11242,G11243,G11244,G11245,G11246,G11247,G11248,G11249,G11250,G11251,G11252,G11253,G11254,G11255,G11256,G11257,G11258,G11259,G11260,
       G11261,G11262,G11263,G11264,G11265,G11266,G11267,G11268,G11269,G11270,G11271,G11272,G11273,G11274,G11275,G11276,G11277,G11278,G11279,G11280,
       G11281,G11282,G11283,G11284,G11285,G11286,G11287,G11288,G11289,G11290,G11291,G11292,G11293,G11294,G11295,G11296,G11297,G11298,G11299,G11300,
       G11301,G11302,G11303,G11304,G11305,G11306,G11307,G11308,G11309,G11310,G11311,G11312,G11313,G11314,G11315,G11316,G11317,G11318,G11319,G11320,
       G11321,G11322,G11323,G11324,G11325,G11326,G11327,G11328,G11329,G11330,G11331,G11332,G11333,G11334,G11335,G11336,G11337,G11338,G11339,G11340,
       G11341,G11342,G11343,G11344,G11345,G11346,G11347,G11348,G11349,G11350,G11351,G11352,G11353,G11354,G11355,G11356,G11357,G11358,G11359,G11360,
       G11361,G11362,G11363,G11364,G11365,G11366,G11367,G11368,G11369,G11370,G11371,G11372,G11373,G11374,G11375,G11376,G11377,G11378,G11379,G11380,
       G11381,G11382,G11383,G11384,G11385,G11386,G11387,G11388,G11389,G11390,G11391,G11392,G11393,G11394,G11395,G11396,G11397,G11398,G11399,G11400,
       G11401,G11402,G11403,G11404,G11405,G11406,G11407,G11408,G11409,G11410,G11411,G11412,G11413,G11414,G11415,G11416,G11417,G11418,G11419,G11420,
       G11421,G11422,G11423,G11424,G11425,G11426,G11427,G11428,G11429,G11430,G11431,G11432,G11433,G11434,G11435,G11436,G11437,G11438,G11439,G11440,
       G11441,G11442,G11443,G11444,G11445,G11446,G11447,G11448,G11449,G11450,G11451,G11452,G11453,G11454,G11455,G11456,G11457,G11458,G11459,G11460,
       G11461,G11462,G11463,G11464,G11465,G11466,G11467,G11468,G11469,G11470,G11471,G11472,G11473,G11474,G11475,G11476,G11477,G11478,G11479,G11480,
       G11481,G11482,G11483,G11484,G11485,G11486,G11487,G11488,G11489,G11490,G11491,G11492,G11493,G11494,G11495,G11496,G11497,G11498,G11499,G11500,
       G11501,G11502,G11503,G11504,G11505,G11506,G11507,G11508,G11509,G11510,G11511,G11512,G11513,G11514,G11515,G11516,G11517,G11518,G11519,G11520,
       G11521,G11522,G11523,G11524,G11525,G11526,G11527,G11528,G11529,G11530,G11531,G11532,G11533,G11534,G11535,G11536,G11537,G11538,G11539,G11540,
       G11541,G11542,G11543,G11544,G11545,G11546,G11547,G11548,G11549,G11550,G11551,G11552,G11553,G11554,G11555,G11556,G11557,G11558,G11559,G11560,
       G11561,G11562,G11563,G11564,G11565,G11566,G11567,G11568,G11569,G11570,G11571,G11572,G11573,G11574,G11575,G11576,G11577,G11578,G11579,G11580,
       G11581,G11582,G11583,G11584,G11585,G11586,G11587,G11588,G11589,G11590,G11591,G11592,G11593,G11594,G11595,G11596,G11597,G11598,G11599,G11600,
       G11601,G11602,G11603,G11604,G11605,G11606,G11607,G11608,G11609,G11610,G11611,G11612,G11613,G11614,G11615,G11616,G11617,G11618,G11619,G11620,
       G11621,G11622,G11623,G11624,G11625,G11626,G11627,G11628,G11629,G11630,G11631,G11632,G11633,G11634,G11635,G11636,G11637,G11638,G11639,G11640,
       G11641,G11642,G11643,G11644,G11645,G11646,G11647,G11648,G11649,G11650,G11651,G11652,G11653,G11654,G11655,G11656,G11657,G11658,G11659,G11660,
       G11661,G11662,G11663,G11664,G11665,G11666,G11667,G11668,G11669,G11670,G11671,G11672,G11673,G11674,G11675,G11676,G11677,G11678,G11679,G11680,
       G11681,G11682,G11683,G11684,G11685,G11686,G11687,G11688,G11689,G11690,G11691,G11692,G11693,G11694,G11695,G11696,G11697,G11698,G11699,G11700,
       G11701,G11702,G11703,G11704,G11705,G11706,G11707,G11708,G11709,G11710,G11711,G11712,G11713,G11714,G11715,G11716,G11717,G11718,G11719,G11720,
       G11721,G11722,G11723,G11724,G11725,G11726,G11727,G11728,G11729,G11730,G11731,G11732,G11733,G11734,G11735,G11736,G11737,G11738,G11739,G11740,
       G11741,G11742,G11743,G11744,G11745,G11746,G11747,G11748,G11749,G11750,G11751,G11752,G11753,G11754,G11755,G11756,G11757,G11758,G11759,G11760,
       G11761,G11762,G11763,G11764,G11765,G11766,G11767,G11768,G11769,G11770,G11771,G11772,G11773,G11774,G11775,G11776,G11777,G11778,G11779,G11780,
       G11781,G11782,G11783,G11784,G11785,G11786,G11787,G11788,G11789,G11790,G11791,G11792,G11793,G11794,G11795,G11796,G11797,G11798,G11799,G11800,
       G11801,G11802,G11803,G11804,G11805,G11806,G11807,G11808,G11809,G11810,G11811,G11812,G11813,G11814,G11815,G11816,G11817,G11818,G11819,G11820,
       G11821,G11822,G11823,G11824,G11825,G11826,G11827,G11828,G11829,G11830,G11831,G11832,G11833,G11834,G11835,G11836,G11837,G11838,G11839,G11840,
       G11841,G11842,G11843,G11844,G11845,G11846,G11847,G11848,G11849,G11850,G11851,G11852,G11853,G11854,G11855,G11856,G11857,G11858,G11859,G11860,
       G11861,G11862,G11863,G11864,G11865,G11866,G11867,G11868,G11869,G11870,G11871,G11872,G11873,G11874,G11875,G11876,G11877,G11878,G11879,G11880,
       G11881,G11882,G11883,G11884,G11885,G11886,G11887,G11888,G11889,G11890,G11891,G11892,G11893,G11894,G11895,G11896,G11897,G11898,G11899,G11900,
       G11901,G11902,G11903,G11904,G11905,G11906,G11907,G11908,G11909,G11910,G11911,G11912,G11913,G11914,G11915,G11916,G11917,G11918,G11919,G11920,
       G11921,G11922,G11923,G11924,G11925,G11926,G11927,G11928,G11929,G11930,G11931,G11932,G11933,G11934,G11935,G11936,G11937,G11938,G11939,G11940,
       G11941,G11942,G11943,G11944,G11945,G11946,G11947,G11948,G11949,G11950,G11951,G11952,G11953,G11954,G11955,G11956,G11957,G11958,G11959,G11960,
       G11961,G11962,G11963,G11964,G11965,G11966,G11967,G11968,G11969,G11970,G11971,G11972,G11973,G11974,G11975,G11976,G11977,G11978,G11979,G11980,
       G11981,G11982,G11983,G11984,G11985,G11986,G11987,G11988,G11989,G11990,G11991,G11992,G11993,G11994,G11995,G11996,G11997,G11998,G11999,G12000,
       G12001,G12002,G12003,G12004,G12005,G12006,G12007,G12008,G12009,G12010,G12011,G12012,G12013,G12014,G12015,G12016,G12017,G12018,G12019,G12020,
       G12021,G12022,G12023,G12024,G12025,G12026,G12027,G12028,G12029,G12030,G12031,G12032,G12033,G12034,G12035,G12036,G12037,G12038,G12039,G12040,
       G12041,G12042,G12043,G12044,G12045,G12046,G12047,G12048,G12049,G12050,G12051,G12052,G12053,G12054,G12055,G12056,G12057,G12058,G12059,G12060,
       G12061,G12062,G12063,G12064,G12065,G12066,G12067,G12068,G12069,G12070,G12071,G12072,G12073,G12074,G12075,G12076,G12077,G12078,G12079,G12080,
       G12081,G12082,G12083,G12084,G12085,G12086,G12087,G12088,G12089,G12090,G12091,G12092,G12093,G12094,G12095,G12096,G12097,G12098,G12099,G12100,
       G12101,G12102,G12103,G12104,G12105,G12106,G12107,G12108,G12109,G12110,G12111,G12112,G12113,G12114,G12115,G12116,G12117,G12118,G12119,G12120,
       G12121,G12122,G12123,G12124,G12125,G12126,G12127,G12128,G12129,G12130,G12131,G12132,G12133,G12134,G12135,G12136,G12137,G12138,G12139,G12140,
       G12141,G12142,G12143,G12144,G12145,G12146,G12147,G12148,G12149,G12150,G12151,G12152,G12153,G12154,G12155,G12156,G12157,G12158,G12159,G12160,
       G12161,G12162,G12163,G12164,G12165,G12166,G12167,G12168,G12169,G12170,G12171,G12172,G12173,G12174,G12175,G12176,G12177,G12178,G12179,G12180,
       G12181,G12182,G12183,G12184,G12185,G12186,G12187,G12188,G12189,G12190,G12191,G12192,G12193,G12194,G12195,G12196,G12197,G12198,G12199,G12200,
       G12201,G12202,G12203,G12204,G12205,G12206,G12207,G12208,G12209,G12210,G12211,G12212,G12213,G12214,G12215,G12216,G12217,G12218,G12219,G12220,
       G12221,G12222,G12223,G12224,G12225,G12226,G12227,G12228,G12229,G12230,G12231,G12232,G12233,G12234,G12235,G12236,G12237,G12238,G12239,G12240,
       G12241,G12242,G12243,G12244,G12245,G12246,G12247,G12248,G12249,G12250,G12251,G12252,G12253,G12254,G12255,G12256,G12257,G12258,G12259,G12260,
       G12261,G12262,G12263,G12264,G12265,G12266,G12267,G12268,G12269,G12270,G12271,G12272,G12273,G12274,G12275,G12276,G12277,G12278,G12279,G12280,
       G12281,G12282,G12283,G12284,G12285,G12286,G12287,G12288,G12289,G12290,G12291,G12292,G12293,G12294,G12295,G12296,G12297,G12298,G12299,G12300,
       G12301,G12302,G12303,G12304,G12305,G12306,G12307,G12308,G12309,G12310,G12311,G12312,G12313,G12314,G12315,G12316,G12317,G12318,G12319,G12320,
       G12321,G12322,G12323,G12324,G12325,G12326,G12327,G12328,G12329,G12330,G12331,G12332,G12333,G12334,G12335,G12336,G12337,G12338,G12339,G12340,
       G12341,G12342,G12343,G12344,G12345,G12346,G12347,G12348,G12349,G12350,G12351,G12352,G12353,G12354,G12355,G12356,G12357,G12358,G12359,G12360,
       G12361,G12362,G12363,G12364,G12365,G12366,G12367,G12368,G12369,G12370,G12371,G12372,G12373,G12374,G12375,G12376,G12377,G12378,G12379,G12380,
       G12381,G12382,G12383,G12384,G12385,G12386,G12387,G12388,G12389,G12390,G12391,G12392,G12393,G12394,G12395,G12396,G12397,G12398,G12399,G12400,
       G12401,G12402,G12403,G12404,G12405,G12406,G12407,G12408,G12409,G12410,G12411,G12412,G12413,G12414,G12415,G12416,G12417,G12418,G12419,G12420,
       G12421,G12422,G12423,G12424,G12425,G12426,G12427,G12428,G12429,G12430,G12431,G12432,G12433,G12434,G12435,G12436,G12437,G12438,G12439,G12440,
       G12441,G12442,G12443,G12444,G12445,G12446,G12447,G12448,G12449,G12450,G12451,G12452,G12453,G12454,G12455,G12456,G12457,G12458,G12459,G12460,
       G12461,G12462,G12463,G12464,G12465,G12466,G12467,G12468,G12469,G12470,G12471,G12472,G12473,G12474,G12475,G12476,G12477,G12478,G12479,G12480,
       G12481,G12482,G12483,G12484,G12485,G12486,G12487,G12488,G12489,G12490,G12491,G12492,G12493,G12494,G12495,G12496,G12497,G12498,G12499,G12500,
       G12501,G12502,G12503,G12504,G12505,G12506,G12507,G12508,G12509,G12510,G12511,G12512,G12513,G12514,G12515,G12516,G12517,G12518,G12519,G12520,
       G12521,G12522,G12523,G12524,G12525,G12526,G12527,G12528,G12529,G12530,G12531,G12532,G12533,G12534,G12535,G12536,G12537,G12538,G12539,G12540,
       G12541,G12542,G12543,G12544,G12545,G12546,G12547,G12548,G12549,G12550,G12551,G12552,G12553,G12554,G12555,G12556,G12557,G12558,G12559,G12560,
       G12561,G12562,G12563,G12564,G12565,G12566,G12567,G12568,G12569,G12570,G12571,G12572,G12573,G12574,G12575,G12576,G12577,G12578,G12579,G12580,
       G12581,G12582,G12583,G12584,G12585,G12586,G12587,G12588,G12589,G12590,G12591,G12592,G12593,G12594,G12595,G12596,G12597,G12598,G12599,G12600,
       G12601,G12602,G12603,G12604,G12605,G12606,G12607,G12608,G12609,G12610,G12611,G12612,G12613,G12614,G12615,G12616,G12617,G12618,G12619,G12620,
       G12621,G12622,G12623,G12624,G12625,G12626,G12627,G12628,G12629,G12630,G12631,G12632,G12633,G12634,G12635,G12636,G12637,G12638,G12639,G12640,
       G12641,G12642,G12643,G12644,G12645,G12646,G12647,G12648,G12649,G12650,G12651,G12652,G12653,G12654,G12655,G12656,G12657,G12658,G12659,G12660,
       G12661,G12662,G12663,G12664,G12665,G12666,G12667,G12668,G12669,G12670,G12671,G12672,G12673,G12674,G12675,G12676,G12677,G12678,G12679,G12680,
       G12681,G12682,G12683,G12684,G12685,G12686,G12687,G12688,G12689,G12690,G12691,G12692,G12693,G12694,G12695,G12696,G12697,G12698,G12699,G12700,
       G12701,G12702,G12703,G12704,G12705,G12706,G12707,G12708,G12709,G12710,G12711,G12712,G12713,G12714,G12715,G12716,G12717,G12718,G12719,G12720,
       G12721,G12722,G12723,G12724,G12725,G12726,G12727,G12728,G12729,G12730,G12731,G12732,G12733,G12734,G12735,G12736,G12737,G12738,G12739,G12740,
       G12741,G12742,G12743,G12744,G12745,G12746,G12747,G12748,G12749,G12750,G12751,G12752,G12753,G12754,G12755,G12756,G12757,G12758,G12759,G12760,
       G12761,G12762,G12763,G12764,G12765,G12766,G12767,G12768,G12769,G12770,G12771,G12772,G12773,G12774,G12775,G12776,G12777,G12778,G12779,G12780,
       G12781,G12782,G12783,G12784,G12785,G12786,G12787,G12788,G12789,G12790,G12791,G12792,G12793,G12794,G12795,G12796,G12797,G12798,G12799,G12800,
       G12801,G12802,G12803,G12804,G12805,G12806,G12807,G12808,G12809,G12810,G12811,G12812,G12813,G12814,G12815,G12816,G12817,G12818,G12819,G12820,
       G12821,G12822,G12823,G12824,G12825,G12826,G12827,G12828,G12829,G12830,G12831,G12832,G12833,G12834,G12835,G12836,G12837,G12838,G12839,G12840,
       G12841,G12842,G12843,G12844,G12845,G12846,G12847,G12848,G12849,G12850,G12851,G12852,G12853,G12854,G12855,G12856,G12857,G12858,G12859,G12860,
       G12861,G12862,G12863,G12864,G12865,G12866,G12867,G12868,G12869,G12870,G12871,G12872,G12873,G12874,G12875,G12876,G12877,G12878,G12879,G12880,
       G12881,G12882,G12883,G12884,G12885,G12886,G12887,G12888,G12889,G12890,G12891,G12892,G12893,G12894,G12895,G12896,G12897,G12898,G12899,G12900,
       G12901,G12902,G12903,G12904,G12905,G12906,G12907,G12908,G12909,G12910,G12911,G12912,G12913,G12914,G12915,G12916,G12917,G12918,G12919,G12920,
       G12921,G12922,G12923,G12924,G12925,G12926,G12927,G12928,G12929,G12930,G12931,G12932,G12933,G12934,G12935,G12936,G12937,G12938,G12939,G12940,
       G12941,G12942,G12943,G12944,G12945,G12946,G12947,G12948,G12949,G12950,G12951,G12952,G12953,G12954,G12955,G12956,G12957,G12958,G12959,G12960,
       G12961,G12962,G12963,G12964,G12965,G12966,G12967,G12968,G12969,G12970,G12971,G12972,G12973,G12974,G12975,G12976,G12977,G12978,G12979,G12980,
       G12981,G12982,G12983,G12984,G12985,G12986,G12987,G12988,G12989,G12990,G12991,G12992,G12993,G12994,G12995,G12996,G12997,G12998,G12999,G13000,
       G13001,G13002,G13003,G13004,G13005,G13006,G13007,G13008,G13009,G13010,G13011,G13012,G13013,G13014,G13015,G13016,G13017,G13018,G13019,G13020,
       G13021,G13022,G13023,G13024,G13025,G13026,G13027,G13028,G13029,G13030,G13031,G13032,G13033,G13034,G13035,G13036,G13037,G13038,G13039,G13040,
       G13041,G13042,G13043,G13044,G13045,G13046,G13047,G13048,G13049,G13050,G13051,G13052,G13053,G13054,G13055,G13056,G13057,G13058,G13059,G13060,
       G13061,G13062,G13063,G13064,G13065,G13066,G13067,G13068,G13069,G13070,G13071,G13072,G13073,G13074,G13075,G13076,G13077,G13078,G13079,G13080,
       G13081,G13082,G13083,G13084,G13085,G13086,G13087,G13088,G13089,G13090,G13091,G13092,G13093,G13094,G13095,G13096,G13097,G13098,G13099,G13100,
       G13101,G13102,G13103,G13104,G13105,G13106,G13107,G13108,G13109,G13110,G13111,G13112,G13113,G13114,G13115,G13116,G13117,G13118,G13119,G13120,
       G13121,G13122,G13123,G13124,G13125,G13126,G13127,G13128,G13129,G13130,G13131,G13132,G13133,G13134,G13135,G13136,G13137,G13138,G13139,G13140,
       G13141,G13142,G13143,G13144,G13145,G13146,G13147,G13148,G13149,G13150,G13151,G13152,G13153,G13154,G13155,G13156,G13157,G13158,G13159,G13160,
       G13161,G13162,G13163,G13164,G13165,G13166,G13167,G13168,G13169,G13170,G13171,G13172,G13173,G13174,G13175,G13176,G13177,G13178,G13179,G13180,
       G13181,G13182,G13183,G13184,G13185,G13186,G13187,G13188,G13189,G13190,G13191,G13192,G13193,G13194,G13195,G13196,G13197,G13198,G13199,G13200,
       G13201,G13202,G13203,G13204,G13205,G13206,G13207,G13208,G13209,G13210,G13211,G13212,G13213,G13214,G13215,G13216,G13217,G13218,G13219,G13220,
       G13221,G13222,G13223,G13224,G13225,G13226,G13227,G13228,G13229,G13230,G13231,G13232,G13233,G13234,G13235,G13236,G13237,G13238,G13239,G13240,
       G13241,G13242,G13243,G13244,G13245,G13246,G13247,G13248,G13249,G13250,G13251,G13252,G13253,G13254,G13255,G13256,G13257,G13258,G13259,G13260,
       G13261,G13262,G13263,G13264,G13265,G13266,G13267,G13268,G13269,G13270,G13271,G13272,G13273,G13274,G13275,G13276,G13277,G13278,G13279,G13280,
       G13281,G13282,G13283,G13284,G13285,G13286,G13287,G13288,G13289,G13290,G13291,G13292,G13293,G13294,G13295,G13296,G13297,G13298,G13299,G13300,
       G13301,G13302,G13303,G13304,G13305,G13306,G13307,G13308,G13309,G13310,G13311,G13312,G13313,G13314,G13315,G13316,G13317,G13318,G13319,G13320,
       G13321,G13322,G13323,G13324,G13325,G13326,G13327,G13328,G13329,G13330,G13331,G13332,G13333,G13334,G13335,G13336,G13337,G13338,G13339,G13340,
       G13341,G13342,G13343,G13344,G13345,G13346,G13347,G13348,G13349,G13350,G13351,G13352,G13353,G13354,G13355,G13356,G13357,G13358,G13359,G13360,
       G13361,G13362,G13363,G13364,G13365,G13366,G13367,G13368,G13369,G13370,G13371,G13372,G13373,G13374,G13375,G13376,G13377,G13378,G13379,G13380,
       G13381,G13382,G13383,G13384,G13385,G13386,G13387,G13388,G13389,G13390,G13391,G13392,G13393,G13394,G13395,G13396,G13397,G13398,G13399,G13400,
       G13401,G13402,G13403,G13404,G13405,G13406,G13407,G13408,G13409,G13410,G13411,G13412,G13413,G13414,G13415,G13416,G13417,G13418,G13419,G13420,
       G13421,G13422,G13423,G13424,G13425,G13426,G13427,G13428,G13429,G13430,G13431,G13432,G13433,G13434,G13435,G13436,G13437,G13438,G13439,G13440,
       G13441,G13442,G13443,G13444,G13445,G13446,G13447,G13448,G13449,G13450,G13451,G13452,G13453,G13454,G13455,G13456,G13457,G13458,G13459,G13460,
       G13461,G13462,G13463,G13464,G13465,G13466,G13467,G13468,G13469,G13470,G13471,G13472,G13473,G13474,G13475,G13476,G13477,G13478,G13479,G13480,
       G13481,G13482,G13483,G13484,G13485,G13486,G13487,G13488,G13489,G13490,G13491,G13492,G13493,G13494,G13495,G13496,G13497,G13498,G13499,G13500,
       G13501,G13502,G13503,G13504,G13505,G13506,G13507,G13508,G13509,G13510,G13511,G13512,G13513,G13514,G13515,G13516,G13517,G13518,G13519,G13520,
       G13521,G13522,G13523,G13524,G13525,G13526,G13527,G13528,G13529,G13530,G13531,G13532,G13533,G13534,G13535,G13536,G13537,G13538,G13539,G13540,
       G13541,G13542,G13543,G13544,G13545,G13546,G13547,G13548,G13549,G13550,G13551,G13552,G13553,G13554,G13555,G13556,G13557,G13558,G13559,G13560,
       G13561,G13562,G13563,G13564,G13565,G13566,G13567,G13568,G13569,G13570,G13571,G13572,G13573,G13574,G13575,G13576,G13577,G13578,G13579,G13580,
       G13581,G13582,G13583,G13584,G13585,G13586,G13587,G13588,G13589,G13590,G13591,G13592,G13593,G13594,G13595,G13596,G13597,G13598,G13599,G13600,
       G13601,G13602,G13603,G13604,G13605,G13606,G13607,G13608,G13609,G13610,G13611,G13612,G13613,G13614,G13615,G13616,G13617,G13618,G13619,G13620,
       G13621,G13622,G13623,G13624,G13625,G13626,G13627,G13628,G13629,G13630,G13631,G13632,G13633,G13634,G13635,G13636,G13637,G13638,G13639,G13640,
       G13641,G13642,G13643,G13644,G13645,G13646,G13647,G13648,G13649,G13650,G13651,G13652,G13653,G13654,G13655,G13656,G13657,G13658,G13659,G13660,
       G13661,G13662,G13663,G13664,G13665,G13666,G13667,G13668,G13669,G13670,G13671,G13672,G13673,G13674,G13675,G13676,G13677,G13678,G13679,G13680,
       G13681,G13682,G13683,G13684,G13685,G13686,G13687,G13688,G13689,G13690,G13691,G13692,G13693,G13694,G13695,G13696,G13697,G13698,G13699,G13700,
       G13701,G13702,G13703,G13704,G13705,G13706,G13707,G13708,G13709,G13710,G13711,G13712,G13713,G13714,G13715,G13716,G13717,G13718,G13719,G13720,
       G13721,G13722,G13723,G13724,G13725,G13726,G13727,G13728,G13729,G13730,G13731,G13732,G13733,G13734,G13735,G13736,G13737,G13738,G13739,G13740,
       G13741,G13742,G13743,G13744,G13745,G13746,G13747,G13748,G13749,G13750,G13751,G13752,G13753,G13754,G13755,G13756,G13757,G13758,G13759,G13760,
       G13761,G13762,G13763,G13764,G13765,G13766,G13767,G13768,G13769,G13770,G13771,G13772,G13773,G13774,G13775,G13776,G13777,G13778,G13779,G13780,
       G13781,G13782,G13783,G13784,G13785,G13786,G13787,G13788,G13789,G13790,G13791,G13792,G13793,G13794,G13795,G13796,G13797,G13798,G13799,G13800,
       G13801,G13802,G13803,G13804,G13805,G13806,G13807,G13808,G13809,G13810,G13811,G13812,G13813,G13814,G13815,G13816,G13817,G13818,G13819,G13820,
       G13821,G13822,G13823,G13824,G13825,G13826,G13827,G13828,G13829,G13830,G13831,G13832,G13833,G13834,G13835,G13836,G13837,G13838,G13839,G13840,
       G13841,G13842,G13843,G13844,G13845,G13846,G13847,G13848,G13849,G13850,G13851,G13852,G13853,G13854,G13855,G13856,G13857,G13858,G13859,G13860,
       G13861,G13862,G13863,G13864,G13865,G13866,G13867,G13868,G13869,G13870,G13871,G13872,G13873,G13874,G13875,G13876,G13877,G13878,G13879,G13880,
       G13881,G13882,G13883,G13884,G13885,G13886,G13887,G13888,G13889,G13890,G13891,G13892,G13893,G13894,G13895,G13896,G13897,G13898,G13899,G13900,
       G13901,G13902,G13903,G13904,G13905,G13906,G13907,G13908,G13909,G13910,G13911,G13912,G13913,G13914,G13915,G13916,G13917,G13918,G13919,G13920,
       G13921,G13922,G13923,G13924,G13925,G13926,G13927,G13928,G13929,G13930,G13931,G13932,G13933,G13934,G13935,G13936,G13937,G13938,G13939,G13940,
       G13941,G13942,G13943,G13944,G13945,G13946,G13947,G13948,G13949,G13950,G13951,G13952,G13953,G13954,G13955,G13956,G13957,G13958,G13959,G13960,
       G13961,G13962,G13963,G13964,G13965,G13966,G13967,G13968,G13969,G13970,G13971,G13972,G13973,G13974,G13975,G13976,G13977,G13978,G13979,G13980,
       G13981,G13982,G13983,G13984,G13985,G13986,G13987,G13988,G13989,G13990,G13991,G13992,G13993,G13994,G13995,G13996,G13997,G13998,G13999,G14000,
       G14001,G14002,G14003,G14004,G14005,G14006,G14007,G14008,G14009,G14010,G14011,G14012,G14013,G14014,G14015,G14016,G14017,G14018,G14019,G14020,
       G14021,G14022,G14023,G14024,G14025,G14026,G14027,G14028,G14029,G14030,G14031,G14032,G14033,G14034,G14035,G14036,G14037,G14038,G14039,G14040,
       G14041,G14042,G14043,G14044,G14045,G14046,G14047,G14048,G14049,G14050,G14051,G14052,G14053,G14054,G14055,G14056,G14057,G14058,G14059,G14060,
       G14061,G14062,G14063,G14064,G14065,G14066,G14067,G14068,G14069,G14070,G14071,G14072,G14073,G14074,G14075,G14076,G14077,G14078,G14079,G14080,
       G14081,G14082,G14083,G14084,G14085,G14086,G14087,G14088,G14089,G14090,G14091,G14092,G14093,G14094,G14095,G14096,G14097,G14098,G14099,G14100,
       G14101,G14102,G14103,G14104,G14105,G14106,G14107,G14108,G14109,G14110,G14111,G14112,G14113,G14114,G14115,G14116,G14117,G14118,G14119,G14120,
       G14121,G14122,G14123,G14124,G14125,G14126,G14127,G14128,G14129,G14130,G14131,G14132,G14133,G14134,G14135,G14136,G14137,G14138,G14139,G14140,
       G14141,G14142,G14143,G14144,G14145,G14146,G14147,G14148,G14149,G14150,G14151,G14152,G14153,G14154,G14155,G14156,G14157,G14158,G14159,G14160,
       G14161,G14162,G14163,G14164,G14165,G14166,G14167,G14168,G14169,G14170,G14171,G14172,G14173,G14174,G14175,G14176,G14177,G14178,G14179,G14180,
       G14181,G14182,G14183,G14184,G14185,G14186,G14187,G14188,G14189,G14190,G14191,G14192,G14193,G14194,G14195,G14196,G14197,G14198,G14199,G14200,
       G14201,G14202,G14203,G14204,G14205,G14206,G14207,G14208,G14209,G14210,G14211,G14212,G14213,G14214,G14215,G14216,G14217,G14218,G14219,G14220,
       G14221,G14222,G14223,G14224,G14225,G14226,G14227,G14228,G14229,G14230,G14231,G14232,G14233,G14234,G14235,G14236,G14237,G14238,G14239,G14240,
       G14241,G14242,G14243,G14244,G14245,G14246,G14247,G14248,G14249,G14250,G14251,G14252,G14253,G14254,G14255,G14256,G14257,G14258,G14259,G14260,
       G14261,G14262,G14263,G14264,G14265,G14266,G14267,G14268,G14269,G14270,G14271,G14272,G14273,G14274,G14275,G14276,G14277,G14278,G14279,G14280,
       G14281,G14282,G14283,G14284,G14285,G14286,G14287,G14288,G14289,G14290,G14291,G14292,G14293,G14294,G14295,G14296,G14297,G14298,G14299,G14300,
       G14301,G14302,G14303,G14304,G14305,G14306,G14307,G14308,G14309,G14310,G14311,G14312,G14313,G14314,G14315,G14316,G14317,G14318,G14319,G14320,
       G14321,G14322,G14323,G14324,G14325,G14326,G14327,G14328,G14329,G14330,G14331,G14332,G14333,G14334,G14335,G14336,G14337,G14338,G14339,G14340,
       G14341,G14342,G14343,G14344,G14345,G14346,G14347,G14348,G14349,G14350,G14351,G14352,G14353,G14354,G14355,G14356,G14357,G14358,G14359,G14360,
       G14361,G14362,G14363,G14364,G14365,G14366,G14367,G14368,G14369,G14370,G14371,G14372,G14373,G14374,G14375,G14376,G14377,G14378,G14379,G14380,
       G14381,G14382,G14383,G14384,G14385,G14386,G14387,G14388,G14389,G14390,G14391,G14392,G14393,G14394,G14395,G14396,G14397,G14398,G14399,G14400,
       G14401,G14402,G14403,G14404,G14405,G14406,G14407,G14408,G14409,G14410,G14411,G14412,G14413,G14414,G14415,G14416,G14417,G14418,G14419,G14420,
       G14421,G14422,G14423,G14424,G14425,G14426,G14427,G14428,G14429,G14430,G14431,G14432,G14433,G14434,G14435,G14436,G14437,G14438,G14439,G14440,
       G14441,G14442,G14443,G14444,G14445,G14446,G14447,G14448,G14449,G14450,G14451,G14452,G14453,G14454,G14455,G14456,G14457,G14458,G14459,G14460,
       G14461,G14462,G14463,G14464,G14465,G14466,G14467,G14468,G14469,G14470,G14471,G14472,G14473,G14474,G14475,G14476,G14477,G14478,G14479,G14480,
       G14481,G14482,G14483,G14484,G14485,G14486,G14487,G14488,G14489,G14490,G14491,G14492,G14493,G14494,G14495,G14496,G14497,G14498,G14499,G14500,
       G14501,G14502,G14503,G14504,G14505,G14506,G14507,G14508,G14509,G14510,G14511,G14512,G14513,G14514,G14515,G14516,G14517,G14518,G14519,G14520,
       G14521,G14522,G14523,G14524,G14525,G14526,G14527,G14528,G14529,G14530,G14531,G14532,G14533,G14534,G14535,G14536,G14537,G14538,G14539,G14540,
       G14541,G14542,G14543,G14544,G14545,G14546,G14547,G14548,G14549,G14550,G14551,G14552,G14553,G14554,G14555,G14556,G14557,G14558,G14559,G14560,
       G14561,G14562,G14563,G14564,G14565,G14566,G14567,G14568,G14569,G14570,G14571,G14572,G14573,G14574,G14575,G14576,G14577,G14578,G14579,G14580,
       G14581,G14582,G14583,G14584,G14585,G14586,G14587,G14588,G14589,G14590,G14591,G14592,G14593,G14594,G14595,G14596,G14597,G14598,G14599,G14600,
       G14601,G14602,G14603,G14604,G14605,G14606,G14607,G14608,G14609,G14610,G14611,G14612,G14613,G14614,G14615,G14616,G14617,G14618,G14619,G14620,
       G14621,G14622,G14623,G14624,G14625,G14626,G14627,G14628,G14629,G14630,G14631,G14632,G14633,G14634,G14635,G14636,G14637,G14638,G14639,G14640,
       G14641,G14642,G14643,G14644,G14645,G14646,G14647,G14648,G14649,G14650,G14651,G14652,G14653,G14654,G14655,G14656,G14657,G14658,G14659,G14660,
       G14661,G14662,G14663,G14664,G14665,G14666,G14667,G14668,G14669,G14670,G14671,G14672,G14673,G14674,G14675,G14676,G14677,G14678,G14679,G14680,
       G14681,G14682,G14683,G14684,G14685,G14686,G14687,G14688,G14689,G14690,G14691,G14692,G14693,G14694,G14695,G14696,G14697,G14698,G14699,G14700,
       G14701,G14702,G14703,G14704,G14705,G14706,G14707,G14708,G14709,G14710,G14711,G14712,G14713,G14714,G14715,G14716,G14717,G14718,G14719,G14720,
       G14721,G14722,G14723,G14724,G14725,G14726,G14727,G14728,G14729,G14730,G14731,G14732,G14733,G14734,G14735,G14736,G14737,G14738,G14739,G14740,
       G14741,G14742,G14743,G14744,G14745,G14746,G14747,G14748,G14749,G14750,G14751,G14752,G14753,G14754,G14755,G14756,G14757,G14758,G14759,G14760,
       G14761,G14762,G14763,G14764,G14765,G14766,G14767,G14768,G14769,G14770,G14771,G14772,G14773,G14774,G14775,G14776,G14777,G14778,G14779,G14780,
       G14781,G14782,G14783,G14784,G14785,G14786,G14787,G14788,G14789,G14790,G14791,G14792,G14793,G14794,G14795,G14796,G14797,G14798,G14799,G14800,
       G14801,G14802,G14803,G14804,G14805,G14806,G14807,G14808,G14809,G14810,G14811,G14812,G14813,G14814,G14815,G14816,G14817,G14818,G14819,G14820,
       G14821,G14822,G14823,G14824,G14825,G14826,G14827,G14828,G14829,G14830,G14831,G14832,G14833,G14834,G14835,G14836,G14837,G14838,G14839,G14840,
       G14841,G14842,G14843,G14844,G14845,G14846,G14847,G14848,G14849,G14850,G14851,G14852,G14853,G14854,G14855,G14856,G14857,G14858,G14859,G14860,
       G14861,G14862,G14863,G14864,G14865,G14866,G14867,G14868,G14869,G14870,G14871,G14872,G14873,G14874,G14875,G14876,G14877,G14878,G14879,G14880,
       G14881,G14882,G14883,G14884,G14885,G14886,G14887,G14888,G14889,G14890,G14891,G14892,G14893,G14894,G14895,G14896,G14897,G14898,G14899,G14900,
       G14901,G14902,G14903,G14904,G14905,G14906,G14907,G14908,G14909,G14910,G14911,G14912,G14913,G14914,G14915,G14916,G14917,G14918,G14919,G14920,
       G14921,G14922,G14923,G14924,G14925,G14926,G14927,G14928,G14929,G14930,G14931,G14932,G14933,G14934,G14935,G14936,G14937,G14938,G14939,G14940,
       G14941,G14942,G14943,G14944,G14945,G14946,G14947,G14948,G14949,G14950,G14951,G14952,G14953,G14954,G14955,G14956,G14957,G14958,G14959,G14960,
       G14961,G14962,G14963,G14964,G14965,G14966,G14967,G14968,G14969,G14970,G14971,G14972,G14973,G14974,G14975,G14976,G14977,G14978,G14979,G14980,
       G14981,G14982,G14983,G14984,G14985,G14986,G14987,G14988,G14989,G14990,G14991,G14992,G14993,G14994,G14995,G14996,G14997,G14998,G14999,G15000,
       G15001,G15002,G15003,G15004,G15005,G15006,G15007,G15008,G15009,G15010,G15011,G15012,G15013,G15014,G15015,G15016,G15017,G15018,G15019,G15020,
       G15021,G15022,G15023,G15024,G15025,G15026,G15027,G15028,G15029,G15030,G15031,G15032,G15033,G15034,G15035,G15036,G15037,G15038,G15039,G15040,
       G15041,G15042,G15043,G15044,G15045,G15046,G15047,G15048,G15049,G15050,G15051,G15052,G15053,G15054,G15055,G15056,G15057,G15058,G15059,G15060,
       G15061,G15062,G15063,G15064,G15065,G15066,G15067,G15068,G15069,G15070,G15071,G15072,G15073,G15074,G15075,G15076,G15077,G15078,G15079,G15080,
       G15081,G15082,G15083,G15084,G15085,G15086,G15087,G15088,G15089,G15090,G15091,G15092,G15093,G15094,G15095,G15096,G15097,G15098,G15099,G15100,
       G15101,G15102,G15103,G15104,G15105,G15106,G15107,G15108,G15109,G15110,G15111,G15112,G15113,G15114,G15115,G15116,G15117,G15118,G15119,G15120,
       G15121,G15122,G15123,G15124,G15125,G15126,G15127,G15128,G15129,G15130,G15131,G15132,G15133,G15134,G15135,G15136,G15137,G15138,G15139,G15140,
       G15141,G15142,G15143,G15144,G15145,G15146,G15147,G15148,G15149,G15150,G15151,G15152,G15153,G15154,G15155,G15156,G15157,G15158,G15159,G15160,
       G15161,G15162,G15163,G15164,G15165,G15166,G15167,G15168,G15169,G15170,G15171,G15172,G15173,G15174,G15175,G15176,G15177,G15178,G15179,G15180,
       G15181,G15182,G15183,G15184,G15185,G15186,G15187,G15188,G15189,G15190,G15191,G15192,G15193,G15194,G15195,G15196,G15197,G15198,G15199,G15200,
       G15201,G15202,G15203,G15204,G15205,G15206,G15207,G15208,G15209,G15210,G15211,G15212,G15213,G15214,G15215,G15216,G15217,G15218,G15219,G15220,
       G15221,G15222,G15223,G15224,G15225,G15226,G15227,G15228,G15229,G15230,G15231,G15232,G15233,G15234,G15235,G15236,G15237,G15238,G15239,G15240,
       G15241,G15242,G15243,G15244,G15245,G15246,G15247,G15248,G15249,G15250,G15251,G15252,G15253,G15254,G15255,G15256,G15257,G15258,G15259,G15260,
       G15261,G15262,G15263,G15264,G15265,G15266,G15267,G15268,G15269,G15270,G15271,G15272,G15273,G15274,G15275,G15276,G15277,G15278,G15279,G15280,
       G15281,G15282,G15283,G15284,G15285,G15286,G15287,G15288,G15289,G15290,G15291,G15292,G15293,G15294,G15295,G15296,G15297,G15298,G15299,G15300,
       G15301,G15302,G15303,G15304,G15305,G15306,G15307,G15308,G15309,G15310,G15311,G15312,G15313,G15314,G15315,G15316,G15317,G15318,G15319,G15320,
       G15321,G15322,G15323,G15324,G15325,G15326,G15327,G15328,G15329,G15330,G15331,G15332,G15333,G15334,G15335,G15336,G15337,G15338,G15339,G15340,
       G15341,G15342,G15343,G15344,G15345,G15346,G15347,G15348,G15349,G15350,G15351,G15352,G15353,G15354,G15355,G15356,G15357,G15358,G15359,G15360,
       G15361,G15362,G15363,G15364,G15365,G15366,G15367,G15368,G15369,G15370,G15371,G15372,G15373,G15374,G15375,G15376,G15377,G15378,G15379,G15380,
       G15381,G15382,G15383,G15384,G15385,G15386,G15387,G15388,G15389,G15390,G15391,G15392,G15393,G15394,G15395,G15396,G15397,G15398,G15399,G15400,
       G15401,G15402,G15403,G15404,G15405,G15406,G15407,G15408,G15409,G15410,G15411,G15412,G15413,G15414,G15415,G15416,G15417,G15418,G15419,G15420,
       G15421,G15422,G15423,G15424,G15425,G15426,G15427,G15428,G15429,G15430,G15431,G15432,G15433,G15434,G15435,G15436,G15437,G15438,G15439,G15440,
       G15441,G15442,G15443,G15444,G15445,G15446,G15447,G15448,G15449,G15450,G15451,G15452,G15453,G15454,G15455,G15456,G15457,G15458,G15459,G15460,
       G15461,G15462,G15463,G15464,G15465,G15466,G15467,G15468,G15469,G15470,G15471,G15472,G15473,G15474,G15475,G15476,G15477,G15478,G15479,G15480,
       G15481,G15482,G15483,G15484,G15485,G15486,G15487,G15488,G15489,G15490,G15491,G15492,G15493,G15494,G15495,G15496,G15497,G15498,G15499,G15500,
       G15501,G15502,G15503,G15504,G15505,G15506,G15507,G15508,G15509,G15510,G15511,G15512,G15513,G15514,G15515,G15516,G15517,G15518,G15519,G15520,
       G15521,G15522,G15523,G15524,G15525,G15526,G15527,G15528,G15529,G15530,G15531,G15532,G15533,G15534,G15535,G15536,G15537,G15538,G15539,G15540,
       G15541,G15542,G15543,G15544,G15545,G15546,G15547,G15548,G15549,G15550,G15551,G15552,G15553,G15554,G15555,G15556,G15557,G15558,G15559,G15560,
       G15561,G15562,G15563,G15564,G15565,G15566,G15567,G15568,G15569,G15570,G15571,G15572,G15573,G15574,G15575,G15576,G15577,G15578,G15579,G15580,
       G15581,G15582,G15583,G15584,G15585,G15586,G15587,G15588,G15589,G15590,G15591,G15592,G15593,G15594,G15595,G15596,G15597,G15598,G15599,G15600,
       G15601,G15602,G15603,G15604,G15605,G15606,G15607,G15608,G15609,G15610,G15611,G15612,G15613,G15614,G15615,G15616,G15617,G15618,G15619,G15620,
       G15621,G15622,G15623,G15624,G15625,G15626,G15627,G15628,G15629,G15630,G15631,G15632,G15633,G15634,G15635,G15636,G15637,G15638,G15639,G15640,
       G15641,G15642,G15643,G15644,G15645,G15646,G15647,G15648,G15649,G15650,G15651,G15652,G15653,G15654,G15655,G15656,G15657,G15658,G15659,G15660,
       G15661,G15662,G15663,G15664,G15665,G15666,G15667,G15668,G15669,G15670,G15671,G15672,G15673,G15674,G15675,G15676,G15677,G15678,G15679,G15680,
       G15681,G15682,G15683,G15684,G15685,G15686,G15687,G15688,G15689,G15690,G15691,G15692,G15693,G15694,G15695,G15696,G15697,G15698,G15699,G15700,
       G15701,G15702,G15703,G15704,G15705,G15706,G15707,G15708,G15709,G15710,G15711,G15712,G15713,G15714,G15715,G15716,G15717,G15718,G15719,G15720,
       G15721,G15722,G15723,G15724,G15725,G15726,G15727,G15728,G15729,G15730,G15731,G15732,G15733,G15734,G15735,G15736,G15737,G15738,G15739,G15740,
       G15741,G15742,G15743,G15744,G15745,G15746,G15747,G15748,G15749,G15750,G15751,G15752,G15753,G15754,G15755,G15756,G15757,G15758,G15759,G15760,
       G15761,G15762,G15763,G15764,G15765,G15766,G15767,G15768,G15769,G15770,G15771,G15772,G15773,G15774,G15775,G15776,G15777,G15778,G15779,G15780,
       G15781,G15782,G15783,G15784,G15785,G15786,G15787,G15788,G15789,G15790,G15791,G15792,G15793,G15794,G15795,G15796,G15797,G15798,G15799,G15800,
       G15801,G15802,G15803,G15804,G15805,G15806,G15807,G15808,G15809,G15810,G15811,G15812,G15813,G15814,G15815,G15816,G15817,G15818,G15819,G15820,
       G15821,G15822,G15823,G15824,G15825,G15826,G15827,G15828,G15829,G15830,G15831,G15832,G15833,G15834,G15835,G15836,G15837,G15838,G15839,G15840,
       G15841,G15842,G15843,G15844,G15845,G15846,G15847,G15848,G15849,G15850,G15851,G15852,G15853,G15854,G15855,G15856,G15857,G15858,G15859,G15860,
       G15861,G15862,G15863,G15864,G15865,G15866,G15867,G15868,G15869,G15870,G15871,G15872,G15873,G15874,G15875,G15876,G15877,G15878,G15879,G15880,
       G15881,G15882,G15883,G15884,G15885,G15886,G15887,G15888,G15889,G15890,G15891,G15892,G15893,G15894,G15895,G15896,G15897,G15898,G15899,G15900,
       G15901,G15902,G15903,G15904,G15905,G15906,G15907,G15908,G15909,G15910,G15911,G15912,G15913,G15914,G15915,G15916,G15917,G15918,G15919,G15920,
       G15921,G15922,G15923,G15924,G15925,G15926,G15927,G15928,G15929,G15930,G15931,G15932,G15933,G15934,G15935,G15936,G15937,G15938,G15939,G15940,
       G15941,G15942,G15943,G15944,G15945,G15946,G15947,G15948,G15949,G15950,G15951,G15952,G15953,G15954,G15955,G15956,G15957,G15958,G15959,G15960,
       G15961,G15962,G15963,G15964,G15965,G15966,G15967,G15968,G15969,G15970,G15971,G15972,G15973,G15974,G15975,G15976,G15977,G15978,G15979,G15980,
       G15981,G15982,G15983,G15984,G15985,G15986,G15987,G15988,G15989,G15990,G15991,G15992,G15993,G15994,G15995,G15996,G15997,G15998,G15999,G16000,
       G16001,G16002,G16003,G16004,G16005,G16006,G16007,G16008,G16009,G16010,G16011,G16012,G16013,G16014,G16015,G16016,G16017,G16018,G16019,G16020,
       G16021,G16022,G16023,G16024,G16025,G16026,G16027,G16028,G16029,G16030,G16031,G16032,G16033,G16034,G16035,G16036,G16037,G16038,G16039,G16040,
       G16041,G16042,G16043,G16044,G16045,G16046,G16047,G16048,G16049,G16050,G16051,G16052,G16053,G16054,G16055,G16056,G16057,G16058,G16059,G16060,
       G16061,G16062,G16063,G16064,G16065,G16066,G16067,G16068,G16069,G16070,G16071,G16072,G16073,G16074,G16075,G16076,G16077,G16078,G16079,G16080,
       G16081,G16082,G16083,G16084,G16085,G16086,G16087,G16088,G16089,G16090,G16091,G16092,G16093,G16094,G16095,G16096,G16097,G16098,G16099,G16100,
       G16101,G16102,G16103,G16104,G16105,G16106,G16107,G16108,G16109,G16110,G16111,G16112,G16113,G16114,G16115,G16116,G16117,G16118,G16119,G16120,
       G16121,G16122,G16123,G16124,G16125,G16126,G16127,G16128,G16129,G16130,G16131,G16132,G16133,G16134,G16135,G16136,G16137,G16138,G16139,G16140,
       G16141,G16142,G16143,G16144,G16145,G16146,G16147,G16148,G16149,G16150,G16151,G16152,G16153,G16154,G16155,G16156,G16157,G16158,G16159,G16160,
       G16161,G16162,G16163,G16164,G16165,G16166,G16167,G16168,G16169,G16170,G16171,G16172,G16173,G16174,G16175,G16176,G16177,G16178,G16179,G16180,
       G16181,G16182,G16183,G16184,G16185,G16186,G16187,G16188,G16189,G16190,G16191,G16192,G16193,G16194,G16195,G16196,G16197,G16198,G16199,G16200,
       G16201,G16202,G16203,G16204,G16205,G16206,G16207,G16208,G16209,G16210,G16211,G16212,G16213,G16214,G16215,G16216,G16217,G16218,G16219,G16220,
       G16221,G16222,G16223,G16224,G16225,G16226,G16227,G16228,G16229,G16230,G16231,G16232,G16233,G16234,G16235,G16236,G16237,G16238,G16239,G16240,
       G16241,G16242,G16243,G16244,G16245,G16246,G16247,G16248,G16249,G16250,G16251,G16252,G16253,G16254,G16255,G16256,G16257,G16258,G16259,G16260,
       G16261,G16262,G16263,G16264,G16265,G16266,G16267,G16268,G16269,G16270,G16271,G16272,G16273,G16274,G16275,G16276,G16277,G16278,G16279,G16280,
       G16281,G16282,G16283,G16284,G16285,G16286,G16287,G16288,G16289,G16290,G16291,G16292,G16293,G16294,G16295,G16296,G16297,G16298,G16299,G16300,
       G16301,G16302,G16303,G16304,G16305,G16306,G16307,G16308,G16309,G16310,G16311,G16312,G16313,G16314,G16315,G16316,G16317,G16318,G16319,G16320,
       G16321,G16322,G16323,G16324,G16325,G16326,G16327,G16328,G16329,G16330,G16331,G16332,G16333,G16334,G16335,G16336,G16337,G16338,G16339,G16340,
       G16341,G16342,G16343,G16344,G16345,G16346,G16347,G16348,G16349,G16350,G16351,G16352,G16353,G16354,G16355,G16356,G16357,G16358,G16359,G16360,
       G16361,G16362,G16363,G16364,G16365,G16366,G16367,G16368,G16369,G16370,G16371,G16372,G16373,G16374,G16375,G16376,G16377,G16378,G16379,G16380,
       G16381,G16382,G16383,G16384,G16385,G16386,G16387,G16388,G16389,G16390,G16391,G16392,G16393,G16394,G16395,G16396,G16397,G16398,G16399,G16400,
       G16401,G16402,G16403,G16404,G16405,G16406,G16407,G16408,G16409,G16410,G16411,G16412,G16413,G16414,G16415,G16416,G16417,G16418,G16419,G16420,
       G16421,G16422,G16423,G16424,G16425,G16426,G16427,G16428,G16429,G16430,G16431,G16432,G16433,G16434,G16435,G16436,G16437,G16438,G16439,G16440,
       G16441,G16442,G16443,G16444,G16445,G16446,G16447,G16448,G16449,G16450,G16451,G16452,G16453,G16454,G16455,G16456,G16457,G16458,G16459,G16460,
       G16461,G16462,G16463,G16464,G16465,G16466,G16467,G16468,G16469,G16470,G16471,G16472,G16473,G16474,G16475,G16476,G16477,G16478,G16479,G16480,
       G16481,G16482,G16483,G16484,G16485,G16486,G16487,G16488,G16489,G16490,G16491,G16492,G16493,G16494,G16495,G16496,G16497,G16498,G16499,G16500,
       G16501,G16502,G16503,G16504,G16505,G16506,G16507,G16508,G16509,G16510,G16511,G16512,G16513,G16514,G16515,G16516,G16517,G16518,G16519,G16520,
       G16521,G16522,G16523,G16524,G16525,G16526,G16527,G16528,G16529,G16530,G16531,G16532,G16533,G16534,G16535,G16536,G16537,G16538,G16539,G16540,
       G16541,G16542,G16543,G16544,G16545,G16546,G16547,G16548,G16549,G16550,G16551,G16552,G16553,G16554,G16555,G16556,G16557,G16558,G16559,G16560,
       G16561,G16562,G16563,G16564,G16565,G16566,G16567,G16568,G16569,G16570,G16571,G16572,G16573,G16574,G16575,G16576,G16577,G16578,G16579,G16580,
       G16581,G16582,G16583,G16584,G16585,G16586,G16587,G16588,G16589,G16590,G16591,G16592,G16593,G16594,G16595,G16596,G16597,G16598,G16599,G16600,
       G16601,G16602,G16603,G16604,G16605,G16606,G16607,G16608,G16609,G16610,G16611,G16612,G16613,G16614,G16615,G16616,G16617,G16618,G16619,G16620,
       G16621,G16622,G16623,G16624,G16625,G16626,G16627,G16628,G16629,G16630,G16631,G16632,G16633,G16634,G16635,G16636,G16637,G16638,G16639,G16640,
       G16641,G16642,G16643,G16644,G16645,G16646,G16647,G16648,G16649,G16650,G16651,G16652,G16653,G16654,G16655,G16656,G16657,G16658,G16659,G16660,
       G16661,G16662,G16663,G16664,G16665,G16666,G16667,G16668,G16669,G16670,G16671,G16672,G16673,G16674,G16675,G16676,G16677,G16678,G16679,G16680,
       G16681,G16682,G16683,G16684,G16685,G16686,G16687,G16688,G16689,G16690,G16691,G16692,G16693,G16694,G16695,G16696,G16697,G16698,G16699,G16700,
       G16701,G16702,G16703,G16704,G16705,G16706,G16707,G16708,G16709,G16710,G16711,G16712,G16713,G16714,G16715,G16716,G16717,G16718,G16719,G16720,
       G16721,G16722,G16723,G16724,G16725,G16726,G16727,G16728,G16729,G16730,G16731,G16732,G16733,G16734,G16735,G16736,G16737,G16738,G16739,G16740,
       G16741,G16742,G16743,G16744,G16745,G16746,G16747,G16748,G16749,G16750,G16751,G16752,G16753,G16754,G16755,G16756,G16757,G16758,G16759,G16760,
       G16761,G16762,G16763,G16764,G16765,G16766,G16767,G16768,G16769,G16770,G16771,G16772,G16773,G16774,G16775,G16776,G16777,G16778,G16779,G16780,
       G16781,G16782,G16783,G16784,G16785,G16786,G16787,G16788,G16789,G16790,G16791,G16792,G16793,G16794,G16795,G16796,G16797,G16798,G16799,G16800,
       G16801,G16802,G16803,G16804,G16805,G16806,G16807,G16808,G16809,G16810,G16811,G16812,G16813,G16814,G16815,G16816,G16817,G16818,G16819,G16820,
       G16821,G16822,G16823,G16824,G16825,G16826,G16827,G16828,G16829,G16830,G16831,G16832,G16833,G16834,G16835,G16836,G16837,G16838,G16839,G16840,
       G16841,G16842,G16843,G16844,G16845,G16846,G16847,G16848,G16849,G16850,G16851,G16852,G16853,G16854,G16855,G16856,G16857,G16858,G16859,G16860,
       G16861,G16862,G16863,G16864,G16865,G16866,G16867,G16868,G16869,G16870,G16871,G16872,G16873,G16874,G16875,G16876,G16877,G16878,G16879,G16880,
       G16881,G16882,G16883,G16884,G16885,G16886,G16887,G16888,G16889,G16890,G16891,G16892,G16893,G16894,G16895,G16896,G16897,G16898,G16899,G16900,
       G16901,G16902,G16903,G16904,G16905,G16906,G16907,G16908,G16909,G16910,G16911,G16912,G16913,G16914,G16915,G16916,G16917,G16918,G16919,G16920,
       G16921,G16922,G16923,G16924,G16925,G16926,G16927,G16928,G16929,G16930,G16931,G16932,G16933,G16934,G16935,G16936,G16937,G16938,G16939,G16940,
       G16941,G16942,G16943,G16944,G16945,G16946,G16947,G16948,G16949,G16950,G16951,G16952,G16953,G16954,G16955,G16956,G16957,G16958,G16959,G16960,
       G16961,G16962,G16963,G16964,G16965,G16966,G16967,G16968,G16969,G16970,G16971,G16972,G16973,G16974,G16975,G16976,G16977,G16978,G16979,G16980,
       G16981,G16982,G16983,G16984,G16985,G16986,G16987,G16988,G16989,G16990,G16991,G16992,G16993,G16994,G16995,G16996,G16997,G16998,G16999,G17000,
       G17001,G17002,G17003,G17004,G17005,G17006,G17007,G17008,G17009,G17010,G17011,G17012,G17013,G17014,G17015,G17016,G17017,G17018,G17019,G17020,
       G17021,G17022,G17023,G17024,G17025,G17026,G17027,G17028,G17029,G17030,G17031,G17032,G17033,G17034,G17035,G17036,G17037,G17038,G17039,G17040,
       G17041,G17042,G17043,G17044,G17045,G17046,G17047,G17048,G17049,G17050,G17051,G17052,G17053,G17054,G17055,G17056,G17057,G17058,G17059,G17060,
       G17061,G17062,G17063,G17064,G17065,G17066,G17067,G17068,G17069,G17070,G17071,G17072,G17073,G17074,G17075,G17076,G17077,G17078,G17079,G17080,
       G17081,G17082,G17083,G17084,G17085,G17086,G17087,G17088,G17089,G17090,G17091,G17092,G17093,G17094,G17095,G17096,G17097,G17098,G17099,G17100,
       G17101,G17102,G17103,G17104,G17105,G17106,G17107,G17108,G17109,G17110,G17111,G17112,G17113,G17114,G17115,G17116,G17117,G17118,G17119,G17120,
       G17121,G17122,G17123,G17124,G17125,G17126,G17127,G17128,G17129,G17130,G17131,G17132,G17133,G17134,G17135,G17136,G17137,G17138,G17139,G17140,
       G17141,G17142,G17143,G17144,G17145,G17146,G17147,G17148,G17149,G17150,G17151,G17152,G17153,G17154,G17155,G17156,G17157,G17158,G17159,G17160,
       G17161,G17162,G17163,G17164,G17165,G17166,G17167,G17168,G17169,G17170,G17171,G17172,G17173,G17174,G17175,G17176,G17177,G17178,G17179,G17180,
       G17181,G17182,G17183,G17184,G17185,G17186,G17187,G17188,G17189,G17190,G17191,G17192,G17193,G17194,G17195,G17196,G17197,G17198,G17199,G17200,
       G17201,G17202,G17203,G17204,G17205,G17206,G17207,G17208,G17209,G17210,G17211,G17212,G17213,G17214,G17215,G17216,G17217,G17218,G17219,G17220,
       G17221,G17222,G17223,G17224,G17225,G17226,G17227,G17228,G17229,G17230,G17231,G17232,G17233,G17234,G17235,G17236,G17237,G17238,G17239,G17240,
       G17241,G17242,G17243,G17244,G17245,G17246,G17247,G17248,G17249,G17250,G17251,G17252,G17253,G17254,G17255,G17256,G17257,G17258,G17259,G17260,
       G17261,G17262,G17263,G17264,G17265,G17266,G17267,G17268,G17269,G17270,G17271,G17272,G17273,G17274,G17275,G17276,G17277,G17278,G17279,G17280,
       G17281,G17282,G17283,G17284,G17285,G17286,G17287,G17288,G17289,G17290,G17291,G17292,G17293,G17294,G17295,G17296,G17297,G17298,G17299,G17300,
       G17301,G17302,G17303,G17304,G17305,G17306,G17307,G17308,G17309,G17310,G17311,G17312,G17313,G17314,G17315,G17316,G17317,G17318,G17319,G17320,
       G17321,G17322,G17323,G17324,G17325,G17326,G17327,G17328,G17329,G17330,G17331,G17332,G17333,G17334,G17335,G17336,G17337,G17338,G17339,G17340,
       G17341,G17342,G17343,G17344,G17345,G17346,G17347,G17348,G17349,G17350,G17351,G17352,G17353,G17354,G17355,G17356,G17357,G17358,G17359,G17360,
       G17361,G17362,G17363,G17364,G17365,G17366,G17367,G17368,G17369,G17370,G17371,G17372,G17373,G17374,G17375,G17376,G17377,G17378,G17379,G17380,
       G17381,G17382,G17383,G17384,G17385,G17386,G17387,G17388,G17389,G17390,G17391,G17392,G17393,G17394,G17395,G17396,G17397,G17398,G17399,G17400,
       G17401,G17402,G17403,G17404,G17405,G17406,G17407,G17408,G17409,G17410,G17411,G17412,G17413,G17414,G17415,G17416,G17417,G17418,G17419,G17420,
       G17421,G17422,G17423,G17424,G17425,G17426,G17427,G17428,G17429,G17430,G17431,G17432,G17433,G17434,G17435,G17436,G17437,G17438,G17439,G17440,
       G17441,G17442,G17443,G17444,G17445,G17446,G17447,G17448,G17449,G17450,G17451,G17452,G17453,G17454,G17455,G17456,G17457,G17458,G17459,G17460,
       G17461,G17462,G17463,G17464,G17465,G17466,G17467,G17468,G17469,G17470,G17471,G17472,G17473,G17474,G17475,G17476,G17477,G17478,G17479,G17480,
       G17481,G17482,G17483,G17484,G17485,G17486,G17487,G17488,G17489,G17490,G17491,G17492,G17493,G17494,G17495,G17496,G17497,G17498,G17499,G17500,
       G17501,G17502,G17503,G17504,G17505,G17506,G17507,G17508,G17509,G17510,G17511,G17512,G17513,G17514,G17515,G17516,G17517,G17518,G17519,G17520,
       G17521,G17522,G17523,G17524,G17525,G17526,G17527,G17528,G17529,G17530,G17531,G17532,G17533,G17534,G17535,G17536,G17537,G17538,G17539,G17540,
       G17541,G17542,G17543,G17544,G17545,G17546,G17547,G17548,G17549,G17550,G17551,G17552,G17553,G17554,G17555,G17556,G17557,G17558,G17559,G17560,
       G17561,G17562,G17563,G17564,G17565,G17566,G17567,G17568,G17569,G17570,G17571,G17572,G17573,G17574,G17575,G17576,G17577,G17578,G17579,G17580,
       G17581,G17582,G17583,G17584,G17585,G17586,G17587,G17588,G17589,G17590,G17591,G17592,G17593,G17594,G17595,G17596,G17597,G17598,G17599,G17600,
       G17601,G17602,G17603,G17604,G17605,G17606,G17607,G17608,G17609,G17610,G17611,G17612,G17613,G17614,G17615,G17616,G17617,G17618,G17619,G17620,
       G17621,G17622,G17623,G17624,G17625,G17626,G17627,G17628,G17629,G17630,G17631,G17632,G17633,G17634,G17635,G17636,G17637,G17638,G17639,G17640,
       G17641,G17642,G17643,G17644,G17645,G17646,G17647,G17648,G17649,G17650,G17651,G17652,G17653,G17654,G17655,G17656,G17657,G17658,G17659,G17660,
       G17661,G17662,G17663,G17664,G17665,G17666,G17667,G17668,G17669,G17670,G17671,G17672,G17673,G17674,G17675,G17676,G17677,G17678,G17679,G17680,
       G17681,G17682,G17683,G17684,G17685,G17686,G17687,G17688,G17689,G17690,G17691,G17692,G17693,G17694,G17695,G17696,G17697,G17698,G17699,G17700,
       G17701,G17702,G17703,G17704,G17705,G17706,G17707,G17708,G17709,G17710,G17711,G17712,G17713,G17714,G17715,G17716,G17717,G17718,G17719,G17720,
       G17721,G17722,G17723,G17724,G17725,G17726,G17727,G17728,G17729,G17730,G17731,G17732,G17733,G17734,G17735,G17736,G17737,G17738,G17739,G17740,
       G17741,G17742,G17743,G17744,G17745,G17746,G17747,G17748,G17749,G17750,G17751,G17752,G17753,G17754,G17755,G17756,G17757,G17758,G17759,G17760,
       G17761,G17762,G17763,G17764,G17765,G17766,G17767,G17768,G17769,G17770,G17771,G17772,G17773,G17774,G17775,G17776,G17777,G17778,G17779,G17780,
       G17781,G17782,G17783,G17784,G17785,G17786,G17787,G17788,G17789,G17790,G17791,G17792,G17793,G17794,G17795,G17796,G17797,G17798,G17799,G17800,
       G17801,G17802,G17803,G17804,G17805,G17806,G17807,G17808,G17809,G17810,G17811,G17812,G17813,G17814,G17815,G17816,G17817,G17818,G17819,G17820,
       G17821,G17822,G17823,G17824,G17825,G17826,G17827,G17828,G17829,G17830,G17831,G17832,G17833,G17834,G17835,G17836,G17837,G17838,G17839,G17840,
       G17841,G17842,G17843,G17844,G17845,G17846,G17847,G17848,G17849,G17850,G17851,G17852,G17853,G17854,G17855,G17856,G17857,G17858,G17859,G17860,
       G17861,G17862,G17863,G17864,G17865,G17866,G17867,G17868,G17869,G17870,G17871,G17872,G17873,G17874,G17875,G17876,G17877,G17878,G17879,G17880,
       G17881,G17882,G17883,G17884,G17885,G17886,G17887,G17888,G17889,G17890,G17891,G17892,G17893,G17894,G17895,G17896,G17897,G17898,G17899,G17900,
       G17901,G17902,G17903,G17904,G17905,G17906,G17907,G17908,G17909,G17910,G17911,G17912,G17913,G17914,G17915,G17916,G17917,G17918,G17919,G17920,
       G17921,G17922,G17923,G17924,G17925,G17926,G17927,G17928,G17929,G17930,G17931,G17932,G17933,G17934,G17935,G17936,G17937,G17938,G17939,G17940,
       G17941,G17942,G17943,G17944,G17945,G17946,G17947,G17948,G17949,G17950,G17951,G17952,G17953,G17954,G17955,G17956,G17957,G17958,G17959,G17960,
       G17961,G17962,G17963,G17964,G17965,G17966,G17967,G17968,G17969,G17970,G17971,G17972,G17973,G17974,G17975,G17976,G17977,G17978,G17979,G17980,
       G17981,G17982,G17983,G17984,G17985,G17986,G17987,G17988,G17989,G17990,G17991,G17992,G17993,G17994,G17995,G17996,G17997,G17998,G17999,G18000,
       G18001,G18002,G18003,G18004,G18005,G18006,G18007,G18008,G18009,G18010,G18011,G18012,G18013,G18014,G18015,G18016,G18017,G18018,G18019,G18020,
       G18021,G18022,G18023,G18024,G18025,G18026,G18027,G18028,G18029,G18030,G18031,G18032,G18033,G18034,G18035,G18036,G18037,G18038,G18039,G18040,
       G18041,G18042,G18043,G18044,G18045,G18046,G18047,G18048,G18049,G18050,G18051,G18052,G18053,G18054,G18055,G18056,G18057,G18058,G18059,G18060,
       G18061,G18062,G18063,G18064,G18065,G18066,G18067,G18068,G18069,G18070,G18071,G18072,G18073,G18074,G18075,G18076,G18077,G18078,G18079,G18080,
       G18081,G18082,G18083,G18084,G18085,G18086,G18087,G18088,G18089,G18090,G18091,G18092,G18093,G18094,G18095,G18096,G18097,G18098,G18099,G18100,
       G18101,G18102,G18103,G18104,G18105,G18106,G18107,G18108,G18109,G18110,G18111,G18112,G18113,G18114,G18115,G18116,G18117,G18118,G18119,G18120,
       G18121,G18122,G18123,G18124,G18125,G18126,G18127,G18128,G18129,G18130,G18131,G18132,G18133,G18134,G18135,G18136,G18137,G18138,G18139,G18140,
       G18141,G18142,G18143,G18144,G18145,G18146,G18147,G18148,G18149,G18150,G18151,G18152,G18153,G18154,G18155,G18156,G18157,G18158,G18159,G18160,
       G18161,G18162,G18163,G18164,G18165,G18166,G18167,G18168,G18169,G18170,G18171,G18172,G18173,G18174,G18175,G18176,G18177,G18178,G18179,G18180,
       G18181,G18182,G18183,G18184,G18185,G18186,G18187,G18188,G18189,G18190,G18191,G18192,G18193,G18194,G18195,G18196,G18197,G18198,G18199,G18200,
       G18201,G18202,G18203,G18204,G18205,G18206,G18207,G18208,G18209,G18210,G18211,G18212,G18213,G18214,G18215,G18216,G18217,G18218,G18219,G18220,
       G18221,G18222,G18223,G18224,G18225,G18226,G18227,G18228,G18229,G18230,G18231,G18232,G18233,G18234,G18235,G18236,G18237,G18238,G18239,G18240,
       G18241,G18242,G18243,G18244,G18245,G18246,G18247,G18248,G18249,G18250,G18251,G18252,G18253,G18254,G18255,G18256,G18257,G18258,G18259,G18260,
       G18261,G18262,G18263,G18264,G18265,G18266,G18267,G18268,G18269,G18270,G18271,G18272,G18273,G18274,G18275,G18276,G18277,G18278,G18279,G18280,
       G18281,G18282,G18283,G18284,G18285,G18286,G18287,G18288,G18289,G18290,G18291,G18292,G18293,G18294,G18295,G18296,G18297,G18298,G18299,G18300,
       G18301,G18302,G18303,G18304,G18305,G18306,G18307,G18308,G18309,G18310,G18311,G18312,G18313,G18314,G18315,G18316,G18317,G18318,G18319,G18320,
       G18321,G18322,G18323,G18324,G18325,G18326,G18327,G18328,G18329,G18330,G18331,G18332,G18333,G18334,G18335,G18336,G18337,G18338,G18339,G18340,
       G18341,G18342,G18343,G18344,G18345,G18346,G18347,G18348,G18349,G18350,G18351,G18352,G18353,G18354,G18355,G18356,G18357,G18358,G18359,G18360,
       G18361,G18362,G18363,G18364,G18365,G18366,G18367,G18368,G18369,G18370,G18371,G18372,G18373,G18374,G18375,G18376,G18377,G18378,G18379,G18380,
       G18381,G18382,G18383,G18384,G18385,G18386,G18387,G18388,G18389,G18390,G18391,G18392,G18393,G18394,G18395,G18396,G18397,G18398,G18399,G18400,
       G18401,G18402,G18403,G18404,G18405,G18406,G18407,G18408,G18409,G18410,G18411,G18412,G18413,G18414,G18415,G18416,G18417,G18418,G18419,G18420,
       G18421,G18422,G18423,G18424,G18425,G18426,G18427,G18428,G18429,G18430,G18431,G18432,G18433,G18434,G18435,G18436,G18437,G18438,G18439,G18440,
       G18441,G18442,G18443,G18444,G18445,G18446,G18447,G18448,G18449,G18450,G18451,G18452,G18453,G18454,G18455,G18456,G18457,G18458,G18459,G18460,
       G18461,G18462,G18463,G18464,G18465,G18466,G18467,G18468,G18469,G18470,G18471,G18472,G18473,G18474,G18475,G18476,G18477,G18478,G18479,G18480,
       G18481,G18482,G18483,G18484,G18485,G18486,G18487,G18488,G18489,G18490,G18491,G18492,G18493,G18494,G18495,G18496,G18497,G18498,G18499,G18500,
       G18501,G18502,G18503,G18504,G18505,G18506,G18507,G18508,G18509,G18510,G18511,G18512,G18513,G18514,G18515,G18516,G18517,G18518,G18519,G18520,
       G18521,G18522,G18523,G18524,G18525,G18526,G18527,G18528,G18529,G18530,G18531,G18532,G18533,G18534,G18535,G18536,G18537,G18538,G18539,G18540,
       G18541,G18542,G18543,G18544,G18545,G18546,G18547,G18548,G18549,G18550,G18551,G18552,G18553,G18554,G18555,G18556,G18557,G18558,G18559,G18560,
       G18561,G18562,G18563,G18564,G18565,G18566,G18567,G18568,G18569,G18570,G18571,G18572,G18573,G18574,G18575,G18576,G18577,G18578,G18579,G18580,
       G18581,G18582,G18583,G18584,G18585,G18586,G18587,G18588,G18589,G18590,G18591,G18592,G18593,G18594,G18595,G18596,G18597,G18598,G18599,G18600,
       G18601,G18602,G18603,G18604,G18605,G18606,G18607,G18608,G18609,G18610,G18611,G18612,G18613,G18614,G18615,G18616,G18617,G18618,G18619,G18620,
       G18621,G18622,G18623,G18624,G18625,G18626,G18627,G18628,G18629,G18630,G18631,G18632,G18633,G18634,G18635,G18636,G18637,G18638,G18639,G18640,
       G18641,G18642,G18643,G18644,G18645,G18646,G18647,G18648,G18649,G18650,G18651,G18652,G18653,G18654,G18655,G18656,G18657,G18658,G18659,G18660,
       G18661,G18662,G18663,G18664,G18665,G18666,G18667,G18668,G18669,G18670,G18671,G18672,G18673,G18674,G18675,G18676,G18677,G18678,G18679,G18680,
       G18681,G18682,G18683,G18684,G18685,G18686,G18687,G18688,G18689,G18690,G18691,G18692,G18693,G18694,G18695,G18696,G18697,G18698,G18699,G18700,
       G18701,G18702,G18703,G18704,G18705,G18706,G18707,G18708,G18709,G18710,G18711,G18712,G18713,G18714,G18715,G18716,G18717,G18718,G18719,G18720,
       G18721,G18722,G18723,G18724,G18725,G18726,G18727,G18728,G18729,G18730,G18731,G18732,G18733,G18734,G18735,G18736,G18737,G18738,G18739,G18740,
       G18741,G18742,G18743,G18744,G18745,G18746,G18747,G18748,G18749,G18750,G18751,G18752,G18753,G18754,G18755,G18756,G18757,G18758,G18759,G18760,
       G18761,G18762,G18763,G18764,G18765,G18766,G18767,G18768,G18769,G18770,G18771,G18772,G18773,G18774,G18775,G18776,G18777,G18778,G18779,G18780,
       G18781,G18782,G18783,G18784,G18785,G18786,G18787,G18788,G18789,G18790,G18791,G18792,G18793,G18794,G18795,G18796,G18797,G18798,G18799,G18800,
       G18801,G18802,G18803,G18804,G18805,G18806,G18807,G18808,G18809,G18810,G18811,G18812,G18813,G18814,G18815,G18816,G18817,G18818,G18819,G18820,
       G18821,G18822,G18823,G18824,G18825,G18826,G18827,G18828,G18829,G18830,G18831,G18832,G18833,G18834,G18835,G18836,G18837,G18838,G18839,G18840,
       G18841,G18842,G18843,G18844,G18845,G18846,G18847,G18848,G18849,G18850,G18851,G18852,G18853,G18854,G18855,G18856,G18857,G18858,G18859,G18860,
       G18861,G18862,G18863,G18864,G18865,G18866,G18867,G18868,G18869,G18870,G18871,G18872,G18873,G18874,G18875,G18876,G18877,G18878,G18879,G18880,
       G18881,G18882,G18883,G18884,G18885,G18886,G18887,G18888,G18889,G18890,G18891,G18892,G18893,G18894,G18895,G18896,G18897,G18898,G18899,G18900,
       G18901,G18902,G18903,G18904,G18905,G18906,G18907,G18908,G18909,G18910,G18911,G18912,G18913,G18914,G18915,G18916,G18917,G18918,G18919,G18920,
       G18921,G18922,G18923,G18924,G18925,G18926,G18927,G18928,G18929,G18930,G18931,G18932,G18933,G18934,G18935,G18936,G18937,G18938,G18939,G18940,
       G18941,G18942,G18943,G18944,G18945,G18946,G18947,G18948,G18949,G18950,G18951,G18952,G18953,G18954,G18955,G18956,G18957,G18958,G18959,G18960,
       G18961,G18962,G18963,G18964,G18965,G18966,G18967,G18968,G18969,G18970,G18971,G18972,G18973,G18974,G18975,G18976,G18977,G18978,G18979,G18980,
       G18981,G18982,G18983,G18984,G18985,G18986,G18987,G18988,G18989,G18990,G18991,G18992,G18993,G18994,G18995,G18996,G18997,G18998,G18999,G19000,
       G19001,G19002,G19003,G19004,G19005,G19006,G19007,G19008,G19009,G19010,G19011,G19012,G19013,G19014,G19015,G19016,G19017,G19018,G19019,G19020,
       G19021,G19022,G19023,G19024,G19025,G19026,G19027,G19028,G19029,G19030,G19031,G19032,G19033,G19034,G19035,G19036,G19037,G19038,G19039,G19040,
       G19041,G19042,G19043,G19044,G19045,G19046,G19047,G19048,G19049,G19050,G19051,G19052,G19053,G19054,G19055,G19056,G19057,G19058,G19059,G19060,
       G19061,G19062,G19063,G19064,G19065,G19066,G19067,G19068,G19069,G19070,G19071,G19072,G19073,G19074,G19075,G19076,G19077,G19078,G19079,G19080,
       G19081,G19082,G19083,G19084,G19085,G19086,G19087,G19088,G19089,G19090,G19091,G19092,G19093,G19094,G19095,G19096,G19097,G19098,G19099,G19100,
       G19101,G19102,G19103,G19104,G19105,G19106,G19107,G19108,G19109,G19110,G19111,G19112,G19113,G19114,G19115,G19116,G19117,G19118,G19119,G19120,
       G19121,G19122,G19123,G19124,G19125,G19126,G19127,G19128,G19129,G19130,G19131,G19132,G19133,G19134,G19135,G19136,G19137,G19138,G19139,G19140,
       G19141,G19142,G19143,G19144,G19145,G19146,G19147,G19148,G19149,G19150,G19151,G19152,G19153,G19154,G19155,G19156,G19157,G19158,G19159,G19160,
       G19161,G19162,G19163,G19164,G19165,G19166,G19167,G19168,G19169,G19170,G19171,G19172,G19173,G19174,G19175,G19176,G19177,G19178,G19179,G19180,
       G19181,G19182,G19183,G19184,G19185,G19186,G19187,G19188,G19189,G19190,G19191,G19192,G19193,G19194,G19195,G19196,G19197,G19198,G19199,G19200,
       G19201,G19202,G19203,G19204,G19205,G19206,G19207,G19208,G19209,G19210,G19211,G19212,G19213,G19214,G19215,G19216,G19217,G19218,G19219,G19220,
       G19221,G19222,G19223,G19224,G19225,G19226,G19227,G19228,G19229,G19230,G19231,G19232,G19233,G19234,G19235,G19236,G19237,G19238,G19239,G19240,
       G19241,G19242,G19243,G19244,G19245,G19246,G19247,G19248,G19249,G19250,G19251,G19252,G19253,G19254,G19255,G19256,G19257,G19258,G19259,G19260,
       G19261,G19262,G19263,G19264,G19265,G19266,G19267,G19268,G19269,G19270,G19271,G19272,G19273,G19274,G19275,G19276,G19277,G19278,G19279,G19280,
       G19281,G19282,G19283,G19284,G19285,G19286,G19287,G19288,G19289,G19290,G19291,G19292,G19293,G19294,G19295,G19296,G19297,G19298,G19299,G19300,
       G19301,G19302,G19303,G19304,G19305,G19306,G19307,G19308,G19309,G19310,G19311,G19312,G19313,G19314,G19315,G19316,G19317,G19318,G19319,G19320,
       G19321,G19322,G19323,G19324,G19325,G19326,G19327,G19328,G19329,G19330,G19331,G19332,G19333,G19334,G19335,G19336,G19337,G19338,G19339,G19340,
       G19341,G19342,G19343,G19344,G19345,G19346,G19347,G19348,G19349,G19350,G19351,G19352,G19353,G19354,G19355,G19356,G19357,G19358,G19359,G19360,
       G19361,G19362,G19363,G19364,G19365,G19366,G19367,G19368,G19369,G19370,G19371,G19372,G19373,G19374,G19375,G19376,G19377,G19378,G19379,G19380,
       G19381,G19382,G19383,G19384,G19385,G19386,G19387,G19388,G19389,G19390,G19391,G19392,G19393,G19394,G19395,G19396,G19397,G19398,G19399,G19400,
       G19401,G19402,G19403,G19404,G19405,G19406,G19407,G19408,G19409,G19410,G19411,G19412,G19413,G19414,G19415,G19416,G19417,G19418,G19419,G19420,
       G19421,G19422,G19423,G19424,G19425,G19426,G19427,G19428,G19429,G19430,G19431,G19432,G19433,G19434,G19435,G19436,G19437,G19438,G19439,G19440,
       G19441,G19442,G19443,G19444,G19445,G19446,G19447,G19448,G19449,G19450,G19451,G19452,G19453,G19454,G19455,G19456,G19457,G19458,G19459,G19460,
       G19461,G19462,G19463,G19464,G19465,G19466,G19467,G19468,G19469,G19470,G19471,G19472,G19473,G19474,G19475,G19476,G19477,G19478,G19479,G19480,
       G19481,G19482,G19483,G19484,G19485,G19486,G19487,G19488,G19489,G19490,G19491,G19492,G19493,G19494,G19495,G19496,G19497,G19498,G19499,G19500,
       G19501,G19502,G19503,G19504,G19505,G19506,G19507,G19508,G19509,G19510,G19511,G19512,G19513,G19514,G19515,G19516,G19517,G19518,G19519,G19520,
       G19521,G19522,G19523,G19524,G19525,G19526,G19527,G19528,G19529,G19530,G19531,G19532,G19533,G19534,G19535,G19536,G19537,G19538,G19539,G19540,
       G19541,G19542,G19543,G19544,G19545,G19546,G19547,G19548,G19549,G19550,G19551,G19552,G19553,G19554,G19555,G19556,G19557,G19558,G19559,G19560,
       G19561,G19562,G19563,G19564,G19565,G19566,G19567,G19568,G19569,G19570,G19571,G19572,G19573,G19574,G19575,G19576,G19577,G19578,G19579,G19580,
       G19581,G19582,G19583,G19584,G19585,G19586,G19587,G19588,G19589,G19590,G19591,G19592,G19593,G19594,G19595,G19596,G19597,G19598,G19599,G19600,
       G19601,G19602,G19603,G19604,G19605,G19606,G19607,G19608,G19609,G19610,G19611,G19612,G19613,G19614,G19615,G19616,G19617,G19618,G19619,G19620,
       G19621,G19622,G19623,G19624,G19625,G19626,G19627,G19628,G19629,G19630,G19631,G19632,G19633,G19634,G19635,G19636,G19637,G19638,G19639,G19640,
       G19641,G19642,G19643,G19644,G19645,G19646,G19647,G19648,G19649,G19650,G19651,G19652,G19653,G19654,G19655,G19656,G19657,G19658,G19659,G19660,
       G19661,G19662,G19663,G19664,G19665,G19666,G19667,G19668,G19669,G19670,G19671,G19672,G19673,G19674,G19675,G19676,G19677,G19678,G19679,G19680,
       G19681,G19682,G19683,G19684,G19685,G19686,G19687,G19688,G19689,G19690,G19691,G19692,G19693,G19694,G19695,G19696,G19697,G19698,G19699,G19700,
       G19701,G19702,G19703,G19704,G19705,G19706,G19707,G19708,G19709,G19710,G19711,G19712,G19713,G19714,G19715,G19716,G19717,G19718,G19719,G19720,
       G19721,G19722,G19723,G19724,G19725,G19726,G19727,G19728,G19729,G19730,G19731,G19732,G19733,G19734,G19735,G19736,G19737,G19738,G19739,G19740,
       G19741,G19742,G19743,G19744,G19745,G19746,G19747,G19748,G19749,G19750,G19751,G19752,G19753,G19754,G19755,G19756,G19757,G19758,G19759,G19760,
       G19761,G19762,G19763,G19764,G19765,G19766,G19767,G19768,G19769,G19770,G19771,G19772,G19773,G19774,G19775,G19776,G19777,G19778,G19779,G19780,
       G19781,G19782,G19783,G19784,G19785,G19786,G19787,G19788,G19789,G19790,G19791,G19792,G19793,G19794,G19795,G19796,G19797,G19798,G19799,G19800,
       G19801,G19802,G19803,G19804,G19805,G19806,G19807,G19808,G19809,G19810,G19811,G19812,G19813,G19814,G19815,G19816,G19817,G19818,G19819,G19820,
       G19821,G19822,G19823,G19824,G19825,G19826,G19827,G19828,G19829,G19830,G19831,G19832,G19833,G19834,G19835,G19836,G19837,G19838,G19839,G19840,
       G19841,G19842,G19843,G19844,G19845,G19846,G19847,G19848,G19849,G19850,G19851,G19852,G19853,G19854,G19855,G19856,G19857,G19858,G19859,G19860,
       G19861,G19862,G19863,G19864,G19865,G19866,G19867,G19868,G19869,G19870,G19871,G19872,G19873,G19874,G19875,G19876,G19877,G19878,G19879,G19880,
       G19881,G19882,G19883,G19884,G19885,G19886,G19887,G19888,G19889,G19890,G19891,G19892,G19893,G19894,G19895,G19896,G19897,G19898,G19899,G19900,
       G19901,G19902,G19903,G19904,G19905,G19906,G19907,G19908,G19909,G19910,G19911,G19912,G19913,G19914,G19915,G19916,G19917,G19918,G19919,G19920,
       G19921,G19922,G19923,G19924,G19925,G19926,G19927,G19928,G19929,G19930,G19931,G19932,G19933,G19934,G19935,G19936,G19937,G19938,G19939,G19940,
       G19941,G19942,G19943,G19944,G19945,G19946,G19947,G19948,G19949,G19950,G19951,G19952,G19953,G19954,G19955,G19956,G19957,G19958,G19959,G19960,
       G19961,G19962,G19963,G19964,G19965,G19966,G19967,G19968,G19969,G19970,G19971,G19972,G19973,G19974,G19975,G19976,G19977,G19978,G19979,G19980,
       G19981,G19982,G19983,G19984,G19985,G19986,G19987,G19988,G19989,G19990,G19991,G19992,G19993,G19994,G19995,G19996,G19997,G19998,G19999,G20000,
       G20001,G20002,G20003,G20004,G20005,G20006,G20007,G20008,G20009,G20010,G20011,G20012,G20013,G20014,G20015,G20016,G20017,G20018,G20019,G20020,
       G20021,G20022,G20023,G20024,G20025,G20026,G20027,G20028,G20029,G20030,G20031,G20032,G20033,G20034,G20035,G20036,G20037,G20038,G20039,G20040,
       G20041,G20042,G20043,G20044,G20045,G20046,G20047,G20048,G20049,G20050,G20051,G20052,G20053,G20054,G20055,G20056,G20057,G20058,G20059,G20060,
       G20061,G20062,G20063,G20064,G20065,G20066,G20067,G20068,G20069,G20070,G20071,G20072,G20073,G20074,G20075,G20076,G20077,G20078,G20079,G20080,
       G20081,G20082,G20083,G20084,G20085,G20086,G20087,G20088,G20089,G20090,G20091,G20092,G20093,G20094,G20095,G20096,G20097,G20098,G20099,G20100,
       G20101,G20102,G20103,G20104,G20105,G20106,G20107,G20108,G20109,G20110,G20111,G20112,G20113,G20114,G20115,G20116,G20117,G20118,G20119,G20120,
       G20121,G20122,G20123,G20124,G20125,G20126,G20127,G20128,G20129,G20130,G20131,G20132,G20133,G20134,G20135,G20136,G20137,G20138,G20139,G20140,
       G20141,G20142,G20143,G20144,G20145,G20146,G20147,G20148,G20149,G20150,G20151,G20152,G20153,G20154,G20155,G20156,G20157,G20158,G20159,G20160,
       G20161,G20162,G20163,G20164,G20165,G20166,G20167,G20168,G20169,G20170,G20171,G20172,G20173,G20174,G20175,G20176,G20177,G20178,G20179,G20180,
       G20181,G20182,G20183,G20184,G20185,G20186,G20187,G20188,G20189,G20190,G20191,G20192,G20193,G20194,G20195,G20196,G20197,G20198,G20199,G20200,
       G20201,G20202,G20203,G20204,G20205,G20206,G20207,G20208,G20209,G20210,G20211,G20212,G20213,G20214,G20215,G20216,G20217,G20218,G20219,G20220,
       G20221,G20222,G20223,G20224,G20225,G20226,G20227,G20228,G20229,G20230,G20231,G20232,G20233,G20234,G20235,G20236,G20237,G20238,G20239,G20240,
       G20241,G20242,G20243,G20244,G20245,G20246,G20247,G20248,G20249,G20250,G20251,G20252,G20253,G20254,G20255,G20256,G20257,G20258,G20259,G20260,
       G20261,G20262,G20263,G20264,G20265,G20266,G20267,G20268,G20269,G20270,G20271,G20272,G20273,G20274,G20275,G20276,G20277,G20278,G20279,G20280,
       G20281,G20282,G20283,G20284,G20285,G20286,G20287,G20288,G20289,G20290,G20291,G20292,G20293,G20294,G20295,G20296,G20297,G20298,G20299,G20300,
       G20301,G20302,G20303,G20304,G20305,G20306,G20307,G20308,G20309,G20310,G20311,G20312,G20313,G20314,G20315,G20316,G20317,G20318,G20319,G20320,
       G20321,G20322,G20323,G20324,G20325,G20326,G20327,G20328,G20329,G20330,G20331,G20332,G20333,G20334,G20335,G20336,G20337,G20338,G20339,G20340,
       G20341,G20342,G20343,G20344,G20345,G20346,G20347,G20348,G20349,G20350,G20351,G20352,G20353,G20354,G20355,G20356,G20357,G20358,G20359,G20360,
       G20361,G20362,G20363,G20364,G20365,G20366,G20367,G20368,G20369,G20370,G20371,G20372,G20373,G20374,G20375,G20376,G20377,G20378,G20379,G20380,
       G20381,G20382,G20383,G20384,G20385,G20386,G20387,G20388,G20389,G20390,G20391,G20392,G20393,G20394,G20395,G20396,G20397,G20398,G20399,G20400,
       G20401,G20402,G20403,G20404,G20405,G20406,G20407,G20408,G20409,G20410,G20411,G20412,G20413,G20414,G20415,G20416,G20417,G20418,G20419,G20420,
       G20421,G20422,G20423,G20424,G20425,G20426,G20427,G20428,G20429,G20430,G20431,G20432,G20433,G20434,G20435,G20436,G20437,G20438,G20439,G20440,
       G20441,G20442,G20443,G20444,G20445,G20446,G20447,G20448,G20449,G20450,G20451,G20452,G20453,G20454,G20455,G20456,G20457,G20458,G20459,G20460,
       G20461,G20462,G20463,G20464,G20465,G20466,G20467,G20468,G20469,G20470,G20471,G20472,G20473,G20474,G20475,G20476,G20477,G20478,G20479,G20480,
       G20481,G20482,G20483,G20484,G20485,G20486,G20487,G20488,G20489,G20490,G20491,G20492,G20493,G20494,G20495,G20496,G20497,G20498,G20499,G20500,
       G20501,G20502,G20503,G20504,G20505,G20506,G20507,G20508,G20509,G20510,G20511,G20512,G20513,G20514,G20515,G20516,G20517,G20518,G20519,G20520,
       G20521,G20522,G20523,G20524,G20525,G20526,G20527,G20528,G20529,G20530,G20531,G20532,G20533,G20534,G20535,G20536,G20537,G20538,G20539,G20540,
       G20541,G20542,G20543,G20544,G20545,G20546,G20547,G20548,G20549,G20550,G20551,G20552,G20553,G20554,G20555,G20556,G20557,G20558,G20559,G20560,
       G20561,G20562,G20563,G20564,G20565,G20566,G20567,G20568,G20569,G20570,G20571,G20572,G20573,G20574,G20575,G20576,G20577,G20578,G20579,G20580,
       G20581,G20582,G20583,G20584,G20585,G20586,G20587,G20588,G20589,G20590,G20591,G20592,G20593,G20594,G20595,G20596,G20597,G20598,G20599,G20600,
       G20601,G20602,G20603,G20604,G20605,G20606,G20607,G20608,G20609,G20610,G20611,G20612,G20613,G20614,G20615,G20616,G20617,G20618,G20619,G20620,
       G20621,G20622,G20623,G20624,G20625,G20626,G20627,G20628,G20629,G20630,G20631,G20632,G20633,G20634,G20635,G20636,G20637,G20638,G20639,G20640,
       G20641,G20642,G20643,G20644,G20645,G20646,G20647,G20648,G20649,G20650,G20651,G20652,G20653,G20654,G20655,G20656,G20657,G20658,G20659,G20660,
       G20661,G20662,G20663,G20664,G20665,G20666,G20667,G20668,G20669,G20670,G20671,G20672,G20673,G20674,G20675,G20676,G20677,G20678,G20679,G20680,
       G20681,G20682,G20683,G20684,G20685,G20686,G20687,G20688,G20689,G20690,G20691,G20692,G20693,G20694,G20695,G20696,G20697,G20698,G20699,G20700,
       G20701,G20702,G20703,G20704,G20705,G20706,G20707,G20708,G20709,G20710,G20711,G20712,G20713,G20714,G20715,G20716,G20717,G20718,G20719,G20720,
       G20721,G20722,G20723,G20724,G20725,G20726,G20727,G20728,G20729,G20730,G20731,G20732,G20733,G20734,G20735,G20736,G20737,G20738,G20739,G20740,
       G20741,G20742,G20743,G20744,G20745,G20746,G20747,G20748,G20749,G20750,G20751,G20752,G20753,G20754,G20755,G20756,G20757,G20758,G20759,G20760,
       G20761,G20762,G20763,G20764,G20765,G20766,G20767,G20768,G20769,G20770,G20771,G20772,G20773,G20774,G20775,G20776,G20777,G20778,G20779,G20780,
       G20781,G20782,G20783,G20784,G20785,G20786,G20787,G20788,G20789,G20790,G20791,G20792,G20793,G20794,G20795,G20796,G20797,G20798,G20799,G20800,
       G20801,G20802,G20803,G20804,G20805,G20806,G20807,G20808,G20809,G20810,G20811,G20812,G20813,G20814,G20815,G20816,G20817,G20818,G20819,G20820,
       G20821,G20822,G20823,G20824,G20825,G20826,G20827,G20828,G20829,G20830,G20831,G20832,G20833,G20834,G20835,G20836,G20837,G20838,G20839,G20840,
       G20841,G20842,G20843,G20844,G20845,G20846,G20847,G20848,G20849,G20850,G20851,G20852,G20853,G20854,G20855,G20856,G20857,G20858,G20859,G20860,
       G20861,G20862,G20863,G20864,G20865,G20866,G20867,G20868,G20869,G20870,G20871,G20872,G20873,G20874,G20875,G20876,G20877,G20878,G20879,G20880,
       G20881,G20882,G20883,G20884,G20885,G20886,G20887,G20888,G20889,G20890,G20891,G20892,G20893,G20894,G20895,G20896,G20897,G20898,G20899,G20900,
       G20901,G20902,G20903,G20904,G20905,G20906,G20907,G20908,G20909,G20910,G20911,G20912,G20913,G20914,G20915,G20916,G20917,G20918,G20919,G20920,
       G20921,G20922,G20923,G20924,G20925,G20926,G20927,G20928,G20929,G20930,G20931,G20932,G20933,G20934,G20935,G20936,G20937,G20938,G20939,G20940,
       G20941,G20942,G20943,G20944,G20945,G20946,G20947,G20948,G20949,G20950,G20951,G20952,G20953,G20954,G20955,G20956,G20957,G20958,G20959,G20960,
       G20961,G20962,G20963,G20964,G20965,G20966,G20967,G20968,G20969,G20970,G20971,G20972,G20973,G20974,G20975,G20976,G20977,G20978,G20979,G20980,
       G20981,G20982,G20983,G20984,G20985,G20986,G20987,G20988,G20989,G20990,G20991,G20992,G20993,G20994,G20995,G20996,G20997,G20998,G20999,G21000,
       G21001,G21002,G21003,G21004,G21005,G21006,G21007,G21008,G21009,G21010,G21011,G21012,G21013,G21014,G21015,G21016,G21017,G21018,G21019,G21020,
       G21021,G21022,G21023,G21024,G21025,G21026,G21027,G21028,G21029,G21030,G21031,G21032,G21033,G21034,G21035,G21036,G21037,G21038,G21039,G21040,
       G21041,G21042,G21043,G21044,G21045,G21046,G21047,G21048,G21049,G21050,G21051,G21052,G21053,G21054,G21055,G21056,G21057,G21058,G21059,G21060,
       G21061,G21062,G21063,G21064,G21065,G21066,G21067,G21068,G21069,G21070,G21071,G21072,G21073,G21074,G21075,G21076,G21077,G21078,G21079,G21080,
       G21081,G21082,G21083,G21084,G21085,G21086,G21087,G21088,G21089,G21090,G21091,G21092,G21093,G21094,G21095,G21096,G21097,G21098,G21099,G21100,
       G21101,G21102,G21103,G21104,G21105,G21106,G21107,G21108,G21109,G21110,G21111,G21112,G21113,G21114,G21115,G21116,G21117,G21118,G21119,G21120,
       G21121,G21122,G21123,G21124,G21125,G21126,G21127,G21128,G21129,G21130,G21131,G21132,G21133,G21134,G21135,G21136,G21137,G21138,G21139,G21140,
       G21141,G21142,G21143,G21144,G21145,G21146,G21147,G21148,G21149,G21150,G21151,G21152,G21153,G21154,G21155,G21156,G21157,G21158,G21159,G21160,
       G21161,G21162,G21163,G21164,G21165,G21166,G21167,G21168,G21169,G21170,G21171,G21172,G21173,G21174,G21175,G21176,G21177,G21178,G21179,G21180,
       G21181,G21182,G21183,G21184,G21185,G21186,G21187,G21188,G21189,G21190,G21191,G21192,G21193,G21194,G21195,G21196,G21197,G21198,G21199,G21200,
       G21201,G21202,G21203,G21204,G21205,G21206,G21207,G21208,G21209,G21210,G21211,G21212,G21213,G21214,G21215,G21216,G21217,G21218,G21219,G21220,
       G21221,G21222,G21223,G21224,G21225,G21226,G21227,G21228,G21229,G21230,G21231,G21232,G21233,G21234,G21235,G21236,G21237,G21238,G21239,G21240,
       G21241,G21242,G21243,G21244,G21245,G21246,G21247,G21248,G21249,G21250,G21251,G21252,G21253,G21254,G21255,G21256,G21257,G21258,G21259,G21260,
       G21261,G21262,G21263,G21264,G21265,G21266,G21267,G21268,G21269,G21270,G21271,G21272,G21273,G21274,G21275,G21276,G21277,G21278,G21279,G21280,
       G21281,G21282,G21283,G21284,G21285,G21286,G21287,G21288,G21289,G21290,G21291,G21292,G21293,G21294,G21295,G21296,G21297,G21298,G21299,G21300,
       G21301,G21302,G21303,G21304,G21305,G21306,G21307,G21308,G21309,G21310,G21311,G21312,G21313,G21314,G21315,G21316,G21317,G21318,G21319,G21320,
       G21321,G21322,G21323,G21324,G21325,G21326,G21327,G21328,G21329,G21330,G21331,G21332,G21333,G21334,G21335,G21336,G21337,G21338,G21339,G21340,
       G21341,G21342,G21343,G21344,G21345,G21346,G21347,G21348,G21349,G21350,G21351,G21352,G21353,G21354,G21355,G21356,G21357,G21358,G21359,G21360,
       G21361,G21362,G21363,G21364,G21365,G21366,G21367,G21368,G21369,G21370,G21371,G21372,G21373,G21374,G21375,G21376,G21377,G21378,G21379,G21380,
       G21381,G21382,G21383,G21384,G21385,G21386,G21387,G21388,G21389,G21390,G21391,G21392,G21393,G21394,G21395,G21396,G21397,G21398,G21399,G21400,
       G21401,G21402,G21403,G21404,G21405,G21406,G21407,G21408,G21409,G21410,G21411,G21412,G21413,G21414,G21415,G21416,G21417,G21418,G21419,G21420,
       G21421,G21422,G21423,G21424,G21425,G21426,G21427,G21428,G21429,G21430,G21431,G21432,G21433,G21434,G21435,G21436,G21437,G21438,G21439,G21440,
       G21441,G21442,G21443,G21444,G21445,G21446,G21447,G21448,G21449,G21450,G21451,G21452,G21453,G21454,G21455,G21456,G21457,G21458,G21459,G21460,
       G21461,G21462,G21463,G21464,G21465,G21466,G21467,G21468,G21469,G21470,G21471,G21472,G21473,G21474,G21475,G21476,G21477,G21478,G21479,G21480,
       G21481,G21482,G21483,G21484,G21485,G21486,G21487,G21488,G21489,G21490,G21491,G21492,G21493,G21494,G21495,G21496,G21497,G21498,G21499,G21500,
       G21501,G21502,G21503,G21504,G21505,G21506,G21507,G21508,G21509,G21510,G21511,G21512,G21513,G21514,G21515,G21516,G21517,G21518,G21519,G21520,
       G21521,G21522,G21523,G21524,G21525,G21526,G21527,G21528,G21529,G21530,G21531,G21532,G21533,G21534,G21535,G21536,G21537,G21538,G21539,G21540,
       G21541,G21542,G21543,G21544,G21545,G21546,G21547,G21548,G21549,G21550,G21551,G21552,G21553,G21554,G21555,G21556,G21557,G21558,G21559,G21560,
       G21561,G21562,G21563,G21564,G21565,G21566,G21567,G21568,G21569,G21570,G21571,G21572,G21573,G21574,G21575,G21576,G21577,G21578,G21579,G21580,
       G21581,G21582,G21583,G21584,G21585,G21586,G21587,G21588,G21589,G21590,G21591,G21592,G21593,G21594,G21595,G21596,G21597,G21598,G21599,G21600,
       G21601,G21602,G21603,G21604,G21605,G21606,G21607,G21608,G21609,G21610,G21611,G21612,G21613,G21614,G21615,G21616,G21617,G21618,G21619,G21620,
       G21621,G21622,G21623,G21624,G21625,G21626,G21627,G21628,G21629,G21630,G21631,G21632,G21633,G21634,G21635,G21636,G21637,G21638,G21639,G21640,
       G21641,G21642,G21643,G21644,G21645,G21646,G21647,G21648,G21649,G21650,G21651,G21652,G21653,G21654,G21655,G21656,G21657,G21658,G21659,G21660,
       G21661,G21662,G21663,G21664,G21665,G21666,G21667,G21668,G21669,G21670,G21671,G21672,G21673,G21674,G21675,G21676,G21677,G21678,G21679,G21680,
       G21681,G21682,G21683,G21684,G21685,G21686,G21687,G21688,G21689,G21690,G21691,G21692,G21693,G21694,G21695,G21696,G21697,G21698,G21699,G21700,
       G21701,G21702,G21703,G21704,G21705,G21706,G21707,G21708,G21709,G21710,G21711,G21712,G21713,G21714,G21715,G21716,G21717,G21718,G21719,G21720,
       G21721,G21722,G21723,G21724,G21725,G21726,G21727,G21728,G21729,G21730,G21731,G21732,G21733,G21734,G21735,G21736,G21737,G21738,G21739,G21740,
       G21741,G21742,G21743,G21744,G21745,G21746,G21747,G21748,G21749,G21750,G21751,G21752,G21753,G21754,G21755,G21756,G21757,G21758,G21759,G21760,
       G21761,G21762,G21763,G21764,G21765,G21766,G21767,G21768,G21769,G21770,G21771,G21772,G21773,G21774,G21775,G21776,G21777,G21778,G21779,G21780,
       G21781,G21782,G21783,G21784,G21785,G21786,G21787,G21788,G21789,G21790,G21791,G21792,G21793,G21794,G21795,G21796,G21797,G21798,G21799,G21800,
       G21801,G21802,G21803,G21804,G21805,G21806,G21807,G21808,G21809,G21810,G21811,G21812,G21813,G21814,G21815,G21816,G21817,G21818,G21819,G21820,
       G21821,G21822,G21823,G21824,G21825,G21826,G21827,G21828,G21829,G21830,G21831,G21832,G21833,G21834,G21835,G21836,G21837,G21838,G21839,G21840,
       G21841,G21842,G21843,G21844,G21845,G21846,G21847,G21848,G21849,G21850,G21851,G21852,G21853,G21854,G21855,G21856,G21857,G21858,G21859,G21860,
       G21861,G21862,G21863,G21864,G21865,G21866,G21867,G21868,G21869,G21870,G21871,G21872,G21873,G21874,G21875,G21876,G21877,G21878,G21879,G21880,
       G21881,G21882,G21883,G21884,G21885,G21886,G21887,G21888,G21889,G21890,G21891,G21892,G21893,G21894,G21895,G21896,G21897,G21898,G21899,G21900,
       G21901,G21902,G21903,G21904,G21905,G21906,G21907,G21908,G21909,G21910,G21911,G21912,G21913,G21914,G21915,G21916,G21917,G21918,G21919,G21920,
       G21921,G21922,G21923,G21924,G21925,G21926,G21927,G21928,G21929,G21930,G21931,G21932,G21933,G21934,G21935,G21936,G21937,G21938,G21939,G21940,
       G21941,G21942,G21943,G21944,G21945,G21946,G21947,G21948,G21949,G21950,G21951,G21952,G21953,G21954,G21955,G21956,G21957,G21958,G21959,G21960,
       G21961,G21962,G21963,G21964,G21965,G21966,G21967,G21968,G21969,G21970,G21971,G21972,G21973,G21974,G21975,G21976,G21977,G21978,G21979,G21980,
       G21981,G21982,G21983,G21984,G21985,G21986,G21987,G21988,G21989,G21990,G21991,G21992,G21993,G21994,G21995,G21996,G21997,G21998,G21999,G22000,
       G22001,G22002,G22003,G22004,G22005,G22006,G22007,G22008,G22009,G22010,G22011,G22012,G22013,G22014,G22015,G22016,G22017,G22018,G22019,G22020,
       G22021,G22022,G22023,G22024,G22025,G22026,G22027,G22028,G22029,G22030,G22031,G22032,G22033,G22034,G22035,G22036,G22037,G22038,G22039,G22040,
       G22041,G22042,G22043,G22044,G22045,G22046,G22047,G22048,G22049,G22050,G22051,G22052,G22053,G22054,G22055,G22056,G22057,G22058,G22059,G22060,
       G22061,G22062,G22063,G22064,G22065,G22066,G22067,G22068,G22069,G22070,G22071,G22072,G22073,G22074,G22075,G22076,G22077,G22078,G22079,G22080,
       G22081,G22082,G22083,G22084,G22085,G22086,G22087,G22088,G22089,G22090,G22091,G22092,G22093,G22094,G22095,G22096,G22097,G22098,G22099,G22100,
       G22101,G22102,G22103,G22104,G22105,G22106,G22107,G22108,G22109,G22110,G22111,G22112,G22113,G22114,G22115,G22116,G22117,G22118,G22119,G22120,
       G22121,G22122,G22123,G22124,G22125,G22126,G22127,G22128,G22129,G22130,G22131,G22132,G22133,G22134,G22135,G22136,G22137,G22138,G22139,G22140,
       G22141,G22142,G22143,G22144,G22145,G22146,G22147,G22148,G22149,G22150,G22151,G22152,G22153,G22154,G22155,G22156,G22157,G22158,G22159,G22160,
       G22161,G22162,G22163,G22164,G22165,G22166,G22167,G22168,G22169,G22170,G22171,G22172,G22173,G22174,G22175,G22176,G22177,G22178,G22179,G22180,
       G22181,G22182,G22183,G22184,G22185,G22186,G22187,G22188,G22189,G22190,G22191,G22192,G22193,G22194,G22195,G22196,G22197,G22198,G22199,G22200,
       G22201,G22202,G22203,G22204,G22205,G22206,G22207,G22208,G22209,G22210,G22211,G22212,G22213,G22214,G22215,G22216,G22217,G22218,G22219,G22220,
       G22221,G22222,G22223,G22224,G22225,G22226,G22227,G22228,G22229,G22230,G22231,G22232,G22233,G22234,G22235,G22236,G22237,G22238,G22239,G22240,
       G22241,G22242,G22243,G22244,G22245,G22246,G22247,G22248,G22249,G22250,G22251,G22252,G22253,G22254,G22255,G22256,G22257,G22258,G22259,G22260,
       G22261,G22262,G22263,G22264,G22265,G22266,G22267,G22268,G22269,G22270,G22271,G22272,G22273,G22274,G22275,G22276,G22277,G22278,G22279,G22280,
       G22281,G22282,G22283,G22284,G22285,G22286,G22287,G22288,G22289,G22290,G22291,G22292,G22293,G22294,G22295,G22296,G22297,G22298,G22299,G22300,
       G22301,G22302,G22303,G22304,G22305,G22306,G22307,G22308,G22309,G22310,G22311,G22312,G22313,G22314,G22315,G22316,G22317,G22318,G22319,G22320,
       G22321,G22322,G22323,G22324,G22325,G22326,G22327,G22328,G22329,G22330,G22331,G22332,G22333,G22334,G22335,G22336,G22337,G22338,G22339,G22340,
       G22341,G22342,G22343,G22344,G22345,G22346,G22347,G22348,G22349,G22350,G22351,G22352,G22353,G22354,G22355,G22356,G22357,G22358,G22359,G22360,
       G22361,G22362,G22363,G22364,G22365,G22366,G22367,G22368,G22369,G22370,G22371,G22372,G22373,G22374,G22375,G22376,G22377,G22378,G22379,G22380,
       G22381,G22382,G22383,G22384,G22385,G22386,G22387,G22388,G22389,G22390,G22391,G22392,G22393,G22394,G22395,G22396,G22397,G22398,G22399,G22400,
       G22401,G22402,G22403,G22404,G22405,G22406,G22407,G22408,G22409,G22410,G22411,G22412,G22413,G22414,G22415,G22416,G22417,G22418,G22419,G22420,
       G22421,G22422,G22423,G22424,G22425,G22426,G22427,G22428,G22429,G22430,G22431,G22432,G22433,G22434,G22435,G22436,G22437,G22438,G22439,G22440,
       G22441,G22442,G22443,G22444,G22445,G22446,G22447,G22448,G22449,G22450,G22451,G22452,G22453,G22454,G22455,G22456,G22457,G22458,G22459,G22460,
       G22461,G22462,G22463,G22464,G22465,G22466,G22467,G22468,G22469,G22470,G22471,G22472,G22473,G22474,G22475,G22476,G22477,G22478,G22479,G22480,
       G22481,G22482,G22483,G22484,G22485,G22486,G22487,G22488,G22489,G22490,G22491,G22492,G22493,G22494,G22495,G22496,G22497,G22498,G22499,G22500,
       G22501,G22502,G22503,G22504,G22505,G22506,G22507,G22508,G22509,G22510,G22511,G22512,G22513,G22514,G22515,G22516,G22517,G22518,G22519,G22520,
       G22521,G22522,G22523,G22524,G22525,G22526,G22527,G22528,G22529,G22530,G22531,G22532,G22533,G22534,G22535,G22536,G22537,G22538,G22539,G22540,
       G22541,G22542,G22543,G22544,G22545,G22546,G22547,G22548,G22549,G22550,G22551,G22552,G22553,G22554,G22555,G22556,G22557,G22558,G22559,G22560,
       G22561,G22562,G22563,G22564,G22565,G22566,G22567,G22568,G22569,G22570,G22571,G22572,G22573,G22574,G22575,G22576,G22577,G22578,G22579,G22580,
       G22581,G22582,G22583,G22584,G22585,G22586,G22587,G22588,G22589,G22590,G22591,G22592,G22593,G22594,G22595,G22596,G22597,G22598,G22599,G22600,
       G22601,G22602,G22603,G22604,G22605,G22606,G22607,G22608,G22609,G22610,G22611,G22612,G22613,G22614,G22615,G22616,G22617,G22618,G22619,G22620,
       G22621,G22622,G22623,G22624,G22625,G22626,G22627,G22628,G22629,G22630,G22631,G22632,G22633,G22634,G22635,G22636,G22637,G22638,G22639,G22640,
       G22641,G22642,G22643,G22644,G22645,G22646,G22647,G22648,G22649,G22650,G22651,G22652,G22653,G22654,G22655,G22656,G22657,G22658,G22659,G22660,
       G22661,G22662,G22663,G22664,G22665,G22666,G22667,G22668,G22669,G22670,G22671,G22672,G22673,G22674,G22675,G22676,G22677,G22678,G22679,G22680,
       G22681,G22682,G22683,G22684,G22685,G22686,G22687,G22688,G22689,G22690,G22691,G22692,G22693,G22694,G22695,G22696,G22697,G22698,G22699,G22700,
       G22701,G22702,G22703,G22704,G22705,G22706,G22707,G22708,G22709,G22710,G22711,G22712,G22713,G22714,G22715,G22716,G22717,G22718,G22719,G22720,
       G22721,G22722,G22723,G22724,G22725,G22726,G22727,G22728,G22729,G22730,G22731,G22732,G22733,G22734,G22735,G22736,G22737,G22738,G22739,G22740,
       G22741,G22742,G22743,G22744,G22745,G22746,G22747,G22748,G22749,G22750,G22751,G22752,G22753,G22754,G22755,G22756,G22757,G22758,G22759,G22760,
       G22761,G22762,G22763,G22764,G22765,G22766,G22767,G22768,G22769,G22770,G22771,G22772,G22773,G22774,G22775,G22776,G22777,G22778,G22779,G22780,
       G22781,G22782,G22783,G22784,G22785,G22786,G22787,G22788,G22789,G22790,G22791,G22792,G22793,G22794,G22795,G22796,G22797,G22798,G22799,G22800,
       G22801,G22802,G22803,G22804,G22805,G22806,G22807,G22808,G22809,G22810,G22811,G22812,G22813,G22814,G22815,G22816,G22817,G22818,G22819,G22820,
       G22821,G22822,G22823,G22824,G22825,G22826,G22827,G22828,G22829,G22830,G22831,G22832,G22833,G22834,G22835,G22836,G22837,G22838,G22839,G22840,
       G22841,G22842,G22843,G22844,G22845,G22846,G22847,G22848,G22849,G22850,G22851,G22852,G22853,G22854,G22855,G22856,G22857,G22858,G22859,G22860,
       G22861,G22862,G22863,G22864,G22865,G22866,G22867,G22868,G22869,G22870,G22871,G22872,G22873,G22874,G22875,G22876,G22877,G22878,G22879,G22880,
       G22881,G22882,G22883,G22884,G22885,G22886,G22887,G22888,G22889,G22890,G22891,G22892,G22893,G22894,G22895,G22896,G22897,G22898,G22899,G22900,
       G22901,G22902,G22903,G22904,G22905,G22906,G22907,G22908,G22909,G22910,G22911,G22912,G22913,G22914,G22915,G22916,G22917,G22918,G22919,G22920,
       G22921,G22922,G22923,G22924,G22925,G22926,G22927,G22928,G22929,G22930,G22931,G22932,G22933,G22934,G22935,G22936,G22937,G22938,G22939,G22940,
       G22941,G22942,G22943,G22944,G22945,G22946,G22947,G22948,G22949,G22950,G22951,G22952,G22953,G22954,G22955,G22956,G22957,G22958,G22959,G22960,
       G22961,G22962,G22963,G22964,G22965,G22966,G22967,G22968,G22969,G22970,G22971,G22972,G22973,G22974,G22975,G22976,G22977,G22978,G22979,G22980,
       G22981,G22982,G22983,G22984,G22985,G22986,G22987,G22988,G22989,G22990,G22991,G22992,G22993,G22994,G22995,G22996,G22997,G22998,G22999,G23000,
       G23001,G23002,G23003,G23004,G23005,G23006,G23007,G23008,G23009,G23010,G23011,G23012,G23013,G23014,G23015,G23016,G23017,G23018,G23019,G23020,
       G23021,G23022,G23023,G23024,G23025,G23026,G23027,G23028,G23029,G23030,G23031,G23032,G23033,G23034,G23035,G23036,G23037,G23038,G23039,G23040,
       G23041,G23042,G23043,G23044,G23045,G23046,G23047,G23048,G23049,G23050,G23051,G23052,G23053,G23054,G23055,G23056,G23057,G23058,G23059,G23060,
       G23061,G23062,G23063,G23064,G23065,G23066,G23067,G23068,G23069,G23070,G23071,G23072,G23073,G23074,G23075,G23076,G23077,G23078,G23079,G23080,
       G23081,G23082,G23083,G23084,G23085,G23086,G23087,G23088,G23089,G23090,G23091,G23092,G23093,G23094,G23095,G23096,G23097,G23098,G23099,G23100,
       G23101,G23102,G23103,G23104,G23105,G23106,G23107,G23108,G23109,G23110,G23111,G23112,G23113,G23114,G23115,G23116,G23117,G23118,G23119,G23120,
       G23121,G23122,G23123,G23124,G23125,G23126,G23127,G23128,G23129,G23130,G23131,G23132,G23133,G23134,G23135,G23136,G23137,G23138,G23139,G23140,
       G23141,G23142,G23143,G23144,G23145,G23146,G23147,G23148,G23149,G23150,G23151,G23152,G23153,G23154,G23155,G23156,G23157,G23158,G23159,G23160,
       G23161,G23162,G23163,G23164,G23165,G23166,G23167,G23168,G23169,G23170,G23171,G23172,G23173,G23174,G23175,G23176,G23177,G23178,G23179,G23180,
       G23181,G23182,G23183,G23184,G23185,G23186,G23187,G23188,G23189,G23190,G23191,G23192,G23193,G23194,G23195,G23196,G23197,G23198,G23199,G23200,
       G23201,G23202,G23203,G23204,G23205,G23206,G23207,G23208,G23209,G23210,G23211,G23212,G23213,G23214,G23215,G23216,G23217,G23218,G23219,G23220,
       G23221,G23222,G23223,G23224,G23225,G23226,G23227,G23228,G23229,G23230,G23231,G23232,G23233,G23234,G23235,G23236,G23237,G23238,G23239,G23240,
       G23241,G23242,G23243,G23244,G23245,G23246,G23247,G23248,G23249,G23250,G23251,G23252,G23253,G23254,G23255,G23256,G23257,G23258,G23259,G23260,
       G23261,G23262,G23263,G23264,G23265,G23266,G23267,G23268,G23269,G23270,G23271,G23272,G23273,G23274,G23275,G23276,G23277,G23278,G23279,G23280,
       G23281,G23282,G23283,G23284,G23285,G23286,G23287,G23288,G23289,G23290,G23291,G23292,G23293,G23294,G23295,G23296,G23297,G23298,G23299,G23300,
       G23301,G23302,G23303,G23304,G23305,G23306,G23307,G23308,G23309,G23310,G23311,G23312,G23313,G23314,G23315,G23316,G23317,G23318,G23319,G23320,
       G23321,G23322,G23323,G23324,G23325,G23326,G23327,G23328,G23329,G23330,G23331,G23332,G23333,G23334,G23335,G23336,G23337,G23338,G23339,G23340,
       G23341,G23342,G23343,G23344,G23345,G23346,G23347,G23348,G23349,G23350,G23351,G23352,G23353,G23354,G23355,G23356,G23357,G23358,G23359,G23360,
       G23361,G23362,G23363,G23364,G23365,G23366,G23367,G23368,G23369,G23370,G23371,G23372,G23373,G23374,G23375,G23376,G23377,G23378,G23379,G23380,
       G23381,G23382,G23383,G23384,G23385,G23386,G23387,G23388,G23389,G23390,G23391,G23392,G23393,G23394,G23395,G23396,G23397,G23398,G23399,G23400,
       G23401,G23402,G23403,G23404,G23405,G23406,G23407,G23408,G23409,G23410,G23411,G23412,G23413,G23414,G23415,G23416,G23417,G23418,G23419,G23420,
       G23421,G23422,G23423,G23424,G23425,G23426,G23427,G23428,G23429,G23430,G23431,G23432,G23433,G23434,G23435,G23436,G23437,G23438,G23439,G23440,
       G23441,G23442,G23443,G23444,G23445,G23446,G23447,G23448,G23449,G23450,G23451,G23452,G23453,G23454,G23455,G23456,G23457,G23458,G23459,G23460,
       G23461,G23462,G23463,G23464,G23465,G23466,G23467,G23468,G23469,G23470,G23471,G23472,G23473,G23474,G23475,G23476,G23477,G23478,G23479,G23480,
       G23481,G23482,G23483,G23484,G23485,G23486,G23487,G23488,G23489,G23490,G23491,G23492,G23493,G23494,G23495,G23496,G23497,G23498,G23499,G23500,
       G23501,G23502,G23503,G23504,G23505,G23506,G23507,G23508,G23509,G23510,G23511,G23512,G23513,G23514,G23515,G23516,G23517,G23518,G23519,G23520,
       G23521,G23522,G23523,G23524,G23525,G23526,G23527,G23528,G23529,G23530,G23531,G23532,G23533,G23534,G23535,G23536,G23537,G23538,G23539,G23540,
       G23541,G23542,G23543,G23544,G23545,G23546,G23547,G23548,G23549,G23550,G23551,G23552,G23553,G23554,G23555,G23556,G23557,G23558,G23559,G23560,
       G23561,G23562,G23563,G23564,G23565,G23566,G23567,G23568,G23569,G23570,G23571,G23572,G23573,G23574,G23575,G23576,G23577,G23578,G23579,G23580,
       G23581,G23582,G23583,G23584,G23585,G23586,G23587,G23588,G23589,G23590,G23591,G23592,G23593,G23594,G23595,G23596,G23597,G23598,G23599,G23600,
       G23601,G23602,G23603,G23604,G23605,G23606,G23607,G23608,G23609,G23610,G23611,G23612,G23613,G23614,G23615,G23616,G23617,G23618,G23619,G23620,
       G23621,G23622,G23623,G23624,G23625,G23626,G23627,G23628,G23629,G23630,G23631,G23632,G23633,G23634,G23635,G23636,G23637,G23638,G23639,G23640,
       G23641,G23642,G23643,G23644,G23645,G23646,G23647,G23648,G23649,G23650,G23651,G23652,G23653,G23654,G23655,G23656,G23657,G23658,G23659,G23660,
       G23661,G23662,G23663,G23664,G23665,G23666,G23667,G23668,G23669,G23670,G23671,G23672,G23673,G23674,G23675,G23676,G23677,G23678,G23679,G23680,
       G23681,G23682,G23683,G23684,G23685,G23686,G23687,G23688,G23689,G23690,G23691,G23692,G23693,G23694,G23695,G23696,G23697,G23698,G23699,G23700,
       G23701,G23702,G23703,G23704,G23705,G23706,G23707,G23708,G23709,G23710,G23711,G23712,G23713,G23714,G23715,G23716,G23717,G23718,G23719,G23720,
       G23721,G23722,G23723,G23724,G23725,G23726,G23727,G23728,G23729,G23730,G23731,G23732,G23733,G23734,G23735,G23736,G23737,G23738,G23739,G23740,
       G23741,G23742,G23743,G23744,G23745,G23746,G23747,G23748,G23749,G23750,G23751,G23752,G23753,G23754,G23755,G23756,G23757,G23758,G23759,G23760,
       G23761,G23762,G23763,G23764,G23765,G23766,G23767,G23768,G23769,G23770,G23771,G23772,G23773,G23774,G23775,G23776,G23777,G23778,G23779,G23780,
       G23781,G23782,G23783,G23784,G23785,G23786,G23787,G23788,G23789,G23790,G23791,G23792,G23793,G23794,G23795,G23796,G23797,G23798,G23799,G23800,
       G23801,G23802,G23803,G23804,G23805,G23806,G23807,G23808,G23809,G23810,G23811,G23812,G23813,G23814,G23815,G23816,G23817,G23818,G23819,G23820,
       G23821,G23822,G23823,G23824,G23825,G23826,G23827,G23828,G23829,G23830,G23831,G23832,G23833,G23834,G23835,G23836,G23837,G23838,G23839,G23840,
       G23841,G23842,G23843,G23844,G23845,G23846,G23847,G23848,G23849,G23850,G23851,G23852,G23853,G23854,G23855,G23856,G23857,G23858,G23859,G23860,
       G23861,G23862,G23863,G23864,G23865,G23866,G23867,G23868,G23869,G23870,G23871,G23872,G23873,G23874,G23875,G23876,G23877,G23878,G23879,G23880,
       G23881,G23882,G23883,G23884,G23885,G23886,G23887,G23888,G23889,G23890,G23891,G23892,G23893,G23894,G23895,G23896,G23897,G23898,G23899,G23900,
       G23901,G23902,G23903,G23904,G23905,G23906,G23907,G23908,G23909,G23910,G23911,G23912,G23913,G23914,G23915,G23916,G23917,G23918,G23919,G23920,
       G23921,G23922,G23923,G23924,G23925,G23926,G23927,G23928,G23929,G23930,G23931,G23932,G23933,G23934,G23935,G23936,G23937,G23938,G23939,G23940,
       G23941,G23942,G23943,G23944,G23945,G23946,G23947,G23948,G23949,G23950,G23951,G23952,G23953,G23954,G23955,G23956,G23957,G23958,G23959,G23960,
       G23961,G23962,G23963,G23964,G23965,G23966,G23967,G23968,G23969,G23970,G23971,G23972,G23973,G23974,G23975,G23976,G23977,G23978,G23979,G23980,
       G23981,G23982,G23983,G23984,G23985,G23986,G23987,G23988,G23989,G23990,G23991,G23992,G23993,G23994,G23995,G23996,G23997,G23998,G23999,G24000,
       G24001,G24002,G24003,G24004,G24005,G24006,G24007,G24008,G24009,G24010,G24011,G24012,G24013,G24014,G24015,G24016,G24017,G24018,G24019,G24020,
       G24021,G24022,G24023,G24024,G24025,G24026,G24027,G24028,G24029,G24030,G24031,G24032,G24033,G24034,G24035,G24036,G24037,G24038,G24039,G24040,
       G24041,G24042,G24043,G24044,G24045,G24046,G24047,G24048,G24049,G24050,G24051,G24052,G24053,G24054,G24055,G24056,G24057,G24058,G24059,G24060,
       G24061,G24062,G24063,G24064,G24065,G24066,G24067,G24068,G24069,G24070,G24071,G24072,G24073,G24074,G24075,G24076,G24077,G24078,G24079,G24080,
       G24081,G24082,G24083,G24084,G24085,G24086,G24087,G24088,G24089,G24090,G24091,G24092,G24093,G24094,G24095,G24096,G24097,G24098,G24099,G24100,
       G24101,G24102,G24103,G24104,G24105,G24106,G24107,G24108,G24109,G24110,G24111,G24112,G24113,G24114,G24115,G24116,G24117,G24118,G24119,G24120,
       G24121,G24122,G24123,G24124,G24125,G24126,G24127,G24128,G24129,G24130,G24131,G24132,G24133,G24134,G24135,G24136,G24137,G24138,G24139,G24140,
       G24141,G24142,G24143,G24144,G24145,G24146,G24147,G24148,G24149,G24150,G24151,G24152,G24153,G24154,G24155,G24156,G24157,G24158,G24159,G24160,
       G24161,G24162,G24163,G24164,G24165,G24166,G24167,G24168,G24169,G24170,G24171,G24172,G24173,G24174,G24175,G24176,G24177,G24178,G24179,G24180,
       G24181,G24182,G24183,G24184,G24185,G24186,G24187,G24188,G24189,G24190,G24191,G24192,G24193,G24194,G24195,G24196,G24197,G24198,G24199,G24200,
       G24201,G24202,G24203,G24204,G24205,G24206,G24207,G24208,G24209,G24210,G24211,G24212,G24213,G24214,G24215,G24216,G24217,G24218,G24219,G24220,
       G24221,G24222,G24223,G24224,G24225,G24226,G24227,G24228,G24229,G24230,G24231,G24232,G24233,G24234,G24235,G24236,G24237,G24238,G24239,G24240,
       G24241,G24242,G24243,G24244,G24245,G24246,G24247,G24248,G24249,G24250,G24251,G24252,G24253,G24254,G24255,G24256,G24257,G24258,G24259,G24260,
       G24261,G24262,G24263,G24264,G24265,G24266,G24267,G24268,G24269,G24270,G24271,G24272,G24273,G24274,G24275,G24276,G24277,G24278,G24279,G24280,
       G24281,G24282,G24283,G24284,G24285,G24286,G24287,G24288,G24289,G24290,G24291,G24292,G24293,G24294,G24295,G24296,G24297,G24298,G24299,G24300,
       G24301,G24302,G24303,G24304,G24305,G24306,G24307,G24308,G24309,G24310,G24311,G24312,G24313,G24314,G24315,G24316,G24317,G24318,G24319,G24320,
       G24321,G24322,G24323,G24324,G24325,G24326,G24327,G24328,G24329,G24330,G24331,G24332,G24333,G24334,G24335,G24336,G24337,G24338,G24339,G24340,
       G24341,G24342,G24343,G24344,G24345,G24346,G24347,G24348,G24349,G24350,G24351,G24352,G24353,G24354,G24355,G24356,G24357,G24358,G24359,G24360,
       G24361,G24362,G24363,G24364,G24365,G24366,G24367,G24368,G24369,G24370,G24371,G24372,G24373,G24374,G24375,G24376,G24377,G24378,G24379,G24380,
       G24381,G24382,G24383,G24384,G24385,G24386,G24387,G24388,G24389,G24390,G24391,G24392,G24393,G24394,G24395,G24396,G24397,G24398,G24399,G24400,
       G24401,G24402,G24403,G24404,G24405,G24406,G24407,G24408,G24409,G24410,G24411,G24412,G24413,G24414,G24415,G24416,G24417,G24418,G24419,G24420,
       G24421,G24422,G24423,G24424,G24425,G24426,G24427,G24428,G24429,G24430,G24431,G24432,G24433,G24434,G24435,G24436,G24437,G24438,G24439,G24440,
       G24441,G24442,G24443,G24444,G24445,G24446,G24447,G24448,G24449,G24450,G24451,G24452,G24453,G24454,G24455,G24456,G24457,G24458,G24459,G24460,
       G24461,G24462,G24463,G24464,G24465,G24466,G24467,G24468,G24469,G24470,G24471,G24472,G24473,G24474,G24475,G24476,G24477,G24478,G24479,G24480,
       G24481,G24482,G24483,G24484,G24485,G24486,G24487,G24488,G24489,G24490,G24491,G24492,G24493,G24494,G24495,G24496,G24497,G24498,G24499,G24500,
       G24501,G24502,G24503,G24504,G24505,G24506,G24507,G24508,G24509,G24510,G24511,G24512,G24513,G24514,G24515,G24516,G24517,G24518,G24519,G24520,
       G24521,G24522,G24523,G24524,G24525,G24526,G24527,G24528,G24529,G24530,G24531,G24532,G24533,G24534,G24535,G24536,G24537,G24538,G24539,G24540,
       G24541,G24542,G24543,G24544,G24545,G24546,G24547,G24548,G24549,G24550,G24551,G24552,G24553,G24554,G24555,G24556,G24557,G24558,G24559,G24560,
       G24561,G24562,G24563,G24564,G24565,G24566,G24567,G24568,G24569,G24570,G24571,G24572,G24573,G24574,G24575,G24576,G24577,G24578,G24579,G24580,
       G24581,G24582,G24583,G24584,G24585,G24586,G24587,G24588,G24589,G24590,G24591,G24592,G24593,G24594,G24595,G24596,G24597,G24598,G24599,G24600,
       G24601,G24602,G24603,G24604,G24605,G24606,G24607,G24608,G24609,G24610,G24611,G24612,G24613,G24614,G24615,G24616,G24617,G24618,G24619,G24620,
       G24621,G24622,G24623,G24624,G24625,G24626,G24627,G24628,G24629,G24630,G24631,G24632,G24633,G24634,G24635,G24636,G24637,G24638,G24639,G24640,
       G24641,G24642,G24643,G24644,G24645,G24646,G24647,G24648,G24649,G24650,G24651,G24652,G24653,G24654,G24655,G24656,G24657,G24658,G24659,G24660,
       G24661,G24662,G24663,G24664,G24665,G24666,G24667,G24668,G24669,G24670,G24671,G24672,G24673,G24674,G24675,G24676,G24677,G24678,G24679,G24680,
       G24681,G24682,G24683,G24684,G24685,G24686,G24687,G24688,G24689,G24690,G24691,G24692,G24693,G24694,G24695,G24696,G24697,G24698,G24699,G24700,
       G24701,G24702,G24703,G24704,G24705,G24706,G24707,G24708,G24709,G24710,G24711,G24712,G24713,G24714,G24715,G24716,G24717,G24718,G24719,G24720,
       G24721,G24722,G24723,G24724,G24725,G24726,G24727,G24728,G24729,G24730,G24731,G24732,G24733,G24734,G24735,G24736,G24737,G24738,G24739,G24740,
       G24741,G24742,G24743,G24744,G24745,G24746,G24747,G24748,G24749,G24750,G24751,G24752,G24753,G24754,G24755,G24756,G24757,G24758,G24759,G24760,
       G24761,G24762,G24763,G24764,G24765,G24766,G24767,G24768,G24769,G24770,G24771,G24772,G24773,G24774,G24775,G24776,G24777,G24778,G24779,G24780,
       G24781,G24782,G24783,G24784,G24785,G24786,G24787,G24788,G24789,G24790,G24791,G24792,G24793,G24794,G24795,G24796,G24797,G24798,G24799,G24800,
       G24801,G24802,G24803,G24804,G24805,G24806,G24807,G24808,G24809,G24810,G24811,G24812,G24813,G24814,G24815,G24816,G24817,G24818,G24819,G24820,
       G24821,G24822,G24823,G24824,G24825,G24826,G24827,G24828,G24829,G24830,G24831,G24832,G24833,G24834,G24835,G24836,G24837,G24838,G24839,G24840,
       G24841,G24842,G24843,G24844,G24845,G24846,G24847,G24848,G24849,G24850,G24851,G24852,G24853,G24854,G24855,G24856,G24857,G24858,G24859,G24860,
       G24861,G24862,G24863,G24864,G24865,G24866,G24867,G24868,G24869,G24870,G24871,G24872,G24873,G24874,G24875,G24876,G24877,G24878,G24879,G24880,
       G24881,G24882,G24883,G24884,G24885,G24886,G24887,G24888,G24889,G24890,G24891,G24892,G24893,G24894,G24895,G24896,G24897,G24898,G24899,G24900,
       G24901,G24902,G24903,G24904,G24905,G24906,G24907,G24908,G24909,G24910,G24911,G24912,G24913,G24914,G24915,G24916,G24917,G24918,G24919,G24920,
       G24921,G24922,G24923,G24924,G24925,G24926,G24927,G24928,G24929,G24930,G24931,G24932,G24933,G24934,G24935,G24936,G24937,G24938,G24939,G24940,
       G24941,G24942,G24943,G24944,G24945,G24946,G24947,G24948,G24949,G24950,G24951,G24952,G24953,G24954,G24955,G24956,G24957,G24958,G24959,G24960,
       G24961,G24962,G24963,G24964,G24965,G24966,G24967,G24968,G24969,G24970,G24971,G24972,G24973,G24974,G24975,G24976,G24977,G24978,G24979,G24980,
       G24981,G24982,G24983,G24984,G24985,G24986,G24987,G24988,G24989,G24990,G24991,G24992,G24993,G24994,G24995,G24996,G24997,G24998,G24999,G25000,
       G25001,G25002,G25003,G25004,G25005,G25006,G25007,G25008,G25009,G25010,G25011,G25012,G25013,G25014,G25015,G25016,G25017,G25018,G25019,G25020,
       G25021,G25022,G25023,G25024,G25025,G25026,G25027,G25028,G25029,G25030,G25031,G25032,G25033,G25034,G25035,G25036,G25037,G25038,G25039,G25040,
       G25041,G25042,G25043,G25044,G25045,G25046,G25047,G25048,G25049,G25050,G25051,G25052,G25053,G25054,G25055,G25056,G25057,G25058,G25059,G25060,
       G25061,G25062,G25063,G25064,G25065,G25066,G25067,G25068,G25069,G25070,G25071,G25072,G25073,G25074,G25075,G25076,G25077,G25078,G25079,G25080,
       G25081,G25082,G25083,G25084,G25085,G25086,G25087,G25088,G25089,G25090,G25091,G25092,G25093,G25094,G25095,G25096,G25097,G25098,G25099,G25100,
       G25101,G25102,G25103,G25104,G25105,G25106,G25107,G25108,G25109,G25110,G25111,G25112,G25113,G25114,G25115,G25116,G25117,G25118,G25119,G25120,
       G25121,G25122,G25123,G25124,G25125,G25126,G25127,G25128,G25129,G25130,G25131,G25132,G25133,G25134,G25135,G25136,G25137,G25138,G25139,G25140,
       G25141,G25142,G25143,G25144,G25145,G25146,G25147,G25148,G25149,G25150,G25151,G25152,G25153,G25154,G25155,G25156,G25157,G25158,G25159,G25160,
       G25161,G25162,G25163,G25164,G25165,G25166,G25167,G25168,G25169,G25170,G25171,G25172,G25173,G25174,G25175,G25176,G25177,G25178,G25179,G25180,
       G25181,G25182,G25183,G25184,G25185,G25186,G25187,G25188,G25189,G25190,G25191,G25192,G25193,G25194,G25195,G25196,G25197,G25198,G25199,G25200,
       G25201,G25202,G25203,G25204,G25205,G25206,G25207,G25208,G25209,G25210,G25211,G25212,G25213,G25214,G25215,G25216,G25217,G25218,G25219,G25220,
       G25221,G25222,G25223,G25224,G25225,G25226,G25227,G25228,G25229,G25230,G25231,G25232,G25233,G25234,G25235,G25236,G25237,G25238,G25239,G25240,
       G25241,G25242,G25243,G25244,G25245,G25246,G25247,G25248,G25249,G25250,G25251,G25252,G25253,G25254,G25255,G25256,G25257,G25258,G25259,G25260,
       G25261,G25262,G25263,G25264,G25265,G25266,G25267,G25268,G25269,G25270,G25271,G25272,G25273,G25274,G25275,G25276,G25277,G25278,G25279,G25280,
       G25281,G25282,G25283,G25284,G25285,G25286,G25287,G25288,G25289,G25290,G25291,G25292,G25293,G25294,G25295,G25296,G25297,G25298,G25299,G25300,
       G25301,G25302,G25303,G25304,G25305,G25306,G25307,G25308,G25309,G25310,G25311,G25312,G25313,G25314,G25315,G25316,G25317,G25318,G25319,G25320,
       G25321,G25322,G25323,G25324,G25325,G25326,G25327,G25328,G25329,G25330,G25331,G25332,G25333,G25334,G25335,G25336,G25337,G25338,G25339,G25340,
       G25341,G25342,G25343,G25344,G25345,G25346,G25347,G25348,G25349,G25350,G25351,G25352,G25353,G25354,G25355,G25356,G25357,G25358,G25359,G25360,
       G25361,G25362,G25363,G25364,G25365,G25366,G25367,G25368,G25369,G25370,G25371,G25372,G25373,G25374,G25375,G25376,G25377,G25378,G25379,G25380,
       G25381,G25382,G25383,G25384,G25385,G25386,G25387,G25388,G25389,G25390,G25391,G25392,G25393,G25394,G25395,G25396,G25397,G25398,G25399,G25400,
       G25401,G25402,G25403,G25404,G25405,G25406,G25407,G25408,G25409,G25410,G25411,G25412,G25413,G25414,G25415,G25416,G25417,G25418,G25419,G25420,
       G25421,G25422,G25423,G25424,G25425,G25426,G25427,G25428,G25429,G25430,G25431,G25432,G25433,G25434,G25435,G25436,G25437,G25438,G25439,G25440,
       G25441,G25442,G25443,G25444,G25445,G25446,G25447,G25448,G25449,G25450,G25451,G25452,G25453,G25454,G25455,G25456,G25457,G25458,G25459,G25460,
       G25461,G25462,G25463,G25464,G25465,G25466,G25467,G25468,G25469,G25470,G25471,G25472,G25473,G25474,G25475,G25476,G25477,G25478,G25479,G25480,
       G25481,G25482,G25483,G25484,G25485,G25486,G25487,G25488,G25489,G25490,G25491,G25492,G25493,G25494,G25495,G25496,G25497,G25498,G25499,G25500,
       G25501,G25502,G25503,G25504,G25505,G25506,G25507,G25508,G25509,G25510,G25511,G25512,G25513,G25514,G25515,G25516,G25517,G25518,G25519,G25520,
       G25521,G25522,G25523,G25524,G25525,G25526,G25527,G25528,G25529,G25530,G25531,G25532,G25533,G25534,G25535,G25536,G25537,G25538,G25539,G25540,
       G25541,G25542,G25543,G25544,G25545,G25546,G25547,G25548,G25549,G25550,G25551,G25552,G25553,G25554,G25555,G25556,G25557,G25558,G25559,G25560,
       G25561,G25562,G25563,G25564,G25565,G25566,G25567,G25568,G25569,G25570,G25571,G25572,G25573,G25574,G25575,G25576,G25577,G25578,G25579,G25580,
       G25581,G25582,G25583,G25584,G25585,G25586,G25587,G25588,G25589,G25590,G25591,G25592,G25593,G25594,G25595,G25596,G25597,G25598,G25599,G25600,
       G25601,G25602,G25603,G25604,G25605,G25606,G25607,G25608,G25609,G25610,G25611,G25612,G25613,G25614,G25615,G25616,G25617,G25618,G25619,G25620,
       G25621,G25622,G25623,G25624,G25625,G25626,G25627,G25628,G25629,G25630,G25631,G25632,G25633,G25634,G25635,G25636,G25637,G25638,G25639,G25640,
       G25641,G25642,G25643,G25644,G25645,G25646,G25647,G25648,G25649,G25650,G25651,G25652,G25653,G25654,G25655,G25656,G25657,G25658,G25659,G25660,
       G25661,G25662,G25663,G25664,G25665,G25666,G25667,G25668,G25669,G25670,G25671,G25672,G25673,G25674,G25675,G25676,G25677,G25678,G25679,G25680,
       G25681,G25682,G25683,G25684,G25685,G25686,G25687,G25688,G25689,G25690,G25691,G25692,G25693,G25694,G25695,G25696,G25697,G25698,G25699,G25700,
       G25701,G25702,G25703,G25704,G25705,G25706,G25707,G25708,G25709,G25710,G25711,G25712,G25713,G25714,G25715,G25716,G25717,G25718,G25719,G25720,
       G25721,G25722,G25723,G25724,G25725,G25726,G25727,G25728,G25729,G25730,G25731,G25732,G25733,G25734,G25735,G25736,G25737,G25738,G25739,G25740,
       G25741,G25742,G25743,G25744,G25745,G25746,G25747,G25748,G25749,G25750,G25751,G25752,G25753,G25754,G25755,G25756,G25757,G25758,G25759,G25760,
       G25761,G25762,G25763,G25764,G25765,G25766,G25767,G25768,G25769,G25770,G25771,G25772,G25773,G25774,G25775,G25776,G25777,G25778,G25779,G25780,
       G25781,G25782,G25783,G25784,G25785,G25786,G25787,G25788,G25789,G25790,G25791,G25792,G25793,G25794,G25795,G25796,G25797,G25798,G25799,G25800,
       G25801,G25802,G25803,G25804,G25805,G25806,G25807,G25808,G25809,G25810,G25811,G25812,G25813,G25814,G25815,G25816,G25817,G25818,G25819,G25820,
       G25821,G25822,G25823,G25824,G25825,G25826,G25827,G25828,G25829,G25830,G25831,G25832,G25833,G25834,G25835,G25836,G25837,G25838,G25839,G25840,
       G25841,G25842,G25843,G25844,G25845,G25846,G25847,G25848,G25849,G25850,G25851,G25852,G25853,G25854,G25855,G25856,G25857,G25858,G25859,G25860,
       G25861,G25862,G25863,G25864,G25865,G25866,G25867,G25868,G25869,G25870,G25871,G25872,G25873,G25874,G25875,G25876,G25877,G25878,G25879,G25880,
       G25881,G25882,G25883,G25884,G25885,G25886,G25887,G25888,G25889,G25890,G25891,G25892,G25893,G25894,G25895,G25896,G25897,G25898,G25899,G25900,
       G25901,G25902,G25903,G25904,G25905,G25906,G25907,G25908,G25909,G25910,G25911,G25912,G25913,G25914,G25915,G25916,G25917,G25918,G25919,G25920,
       G25921,G25922,G25923,G25924,G25925,G25926,G25927,G25928,G25929,G25930,G25931,G25932,G25933,G25934,G25935,G25936,G25937,G25938,G25939,G25940,
       G25941,G25942,G25943,G25944,G25945,G25946,G25947,G25948,G25949,G25950,G25951,G25952,G25953,G25954,G25955,G25956,G25957,G25958,G25959,G25960,
       G25961,G25962,G25963,G25964,G25965,G25966,G25967,G25968,G25969,G25970,G25971,G25972,G25973,G25974,G25975,G25976,G25977,G25978,G25979,G25980,
       G25981,G25982,G25983,G25984,G25985,G25986,G25987,G25988,G25989,G25990,G25991,G25992,G25993,G25994,G25995,G25996,G25997,G25998,G25999,G26000,
       G26001,G26002,G26003,G26004,G26005,G26006,G26007,G26008,G26009,G26010,G26011,G26012,G26013,G26014,G26015,G26016,G26017,G26018,G26019,G26020,
       G26021,G26022,G26023,G26024,G26025,G26026,G26027,G26028,G26029,G26030,G26031,G26032,G26033,G26034,G26035,G26036,G26037,G26038,G26039,G26040,
       G26041,G26042,G26043,G26044,G26045,G26046,G26047,G26048,G26049,G26050,G26051,G26052,G26053,G26054,G26055,G26056,G26057,G26058,G26059,G26060,
       G26061,G26062,G26063,G26064,G26065,G26066,G26067,G26068,G26069,G26070,G26071,G26072,G26073,G26074,G26075,G26076,G26077,G26078,G26079,G26080,
       G26081,G26082,G26083,G26084,G26085,G26086,G26087,G26088,G26089,G26090,G26091,G26092,G26093,G26094,G26095,G26096,G26097,G26098,G26099,G26100,
       G26101,G26102,G26103,G26104,G26105,G26106,G26107,G26108,G26109,G26110,G26111,G26112,G26113,G26114,G26115,G26116,G26117,G26118,G26119,G26120,
       G26121,G26122,G26123,G26124,G26125,G26126,G26127,G26128,G26129,G26130,G26131,G26132,G26133,G26134,G26135,G26136,G26137,G26138,G26139,G26140,
       G26141,G26142,G26143,G26144,G26145,G26146,G26147,G26148,G26149,G26150,G26151,G26152,G26153,G26154,G26155,G26156,G26157,G26158,G26159,G26160,
       G26161,G26162,G26163,G26164,G26165,G26166,G26167,G26168,G26169,G26170,G26171,G26172,G26173,G26174,G26175,G26176,G26177,G26178,G26179,G26180,
       G26181,G26182,G26183,G26184,G26185,G26186,G26187,G26188,G26189,G26190,G26191,G26192,G26193,G26194,G26195,G26196,G26197,G26198,G26199,G26200,
       G26201,G26202,G26203,G26204,G26205,G26206,G26207,G26208,G26209,G26210,G26211,G26212,G26213,G26214,G26215,G26216,G26217,G26218,G26219,G26220,
       G26221,G26222,G26223,G26224,G26225,G26226,G26227,G26228,G26229,G26230,G26231,G26232,G26233,G26234,G26235,G26236,G26237,G26238,G26239,G26240,
       G26241,G26242,G26243,G26244,G26245,G26246,G26247,G26248,G26249,G26250,G26251,G26252,G26253,G26254,G26255,G26256,G26257,G26258,G26259,G26260,
       G26261,G26262,G26263,G26264,G26265,G26266,G26267,G26268,G26269,G26270,G26271,G26272,G26273,G26274,G26275,G26276,G26277,G26278,G26279,G26280,
       G26281,G26282,G26283,G26284,G26285,G26286,G26287,G26288,G26289,G26290,G26291,G26292,G26293,G26294,G26295,G26296,G26297,G26298,G26299,G26300,
       G26301,G26302,G26303,G26304,G26305,G26306,G26307,G26308,G26309,G26310,G26311,G26312,G26313,G26314,G26315,G26316,G26317,G26318,G26319,G26320,
       G26321,G26322,G26323,G26324,G26325,G26326,G26327,G26328,G26329,G26330,G26331,G26332,G26333,G26334,G26335,G26336,G26337,G26338,G26339,G26340,
       G26341,G26342,G26343,G26344,G26345,G26346,G26347,G26348,G26349,G26350,G26351,G26352,G26353,G26354,G26355,G26356,G26357,G26358,G26359,G26360,
       G26361,G26362,G26363,G26364,G26365,G26366,G26367,G26368,G26369,G26370,G26371,G26372,G26373,G26374,G26375,G26376,G26377,G26378,G26379,G26380,
       G26381,G26382,G26383,G26384,G26385,G26386,G26387,G26388,G26389,G26390,G26391,G26392,G26393,G26394,G26395,G26396,G26397,G26398,G26399,G26400,
       G26401,G26402,G26403,G26404,G26405,G26406,G26407,G26408,G26409,G26410,G26411,G26412,G26413,G26414,G26415,G26416,G26417,G26418,G26419,G26420,
       G26421,G26422,G26423,G26424,G26425,G26426,G26427,G26428,G26429,G26430,G26431,G26432,G26433,G26434,G26435,G26436,G26437,G26438,G26439,G26440,
       G26441,G26442,G26443,G26444,G26445,G26446,G26447,G26448,G26449,G26450,G26451,G26452,G26453,G26454,G26455,G26456,G26457,G26458,G26459,G26460,
       G26461,G26462,G26463,G26464,G26465,G26466,G26467,G26468,G26469,G26470,G26471,G26472,G26473,G26474,G26475,G26476,G26477,G26478,G26479,G26480,
       G26481,G26482,G26483,G26484,G26485,G26486,G26487,G26488,G26489,G26490,G26491,G26492,G26493,G26494,G26495,G26496,G26497,G26498,G26499,G26500,
       G26501,G26502,G26503,G26504,G26505,G26506,G26507,G26508,G26509,G26510,G26511,G26512,G26513,G26514,G26515,G26516,G26517,G26518,G26519,G26520,
       G26521,G26522,G26523,G26524,G26525,G26526,G26527,G26528,G26529,G26530,G26531,G26532,G26533,G26534,G26535,G26536,G26537,G26538,G26539,G26540,
       G26541,G26542,G26543,G26544,G26545,G26546,G26547,G26548,G26549,G26550,G26551,G26552,G26553,G26554,G26555,G26556,G26557,G26558,G26559,G26560,
       G26561,G26562,G26563,G26564,G26565,G26566,G26567,G26568,G26569,G26570,G26571,G26572,G26573,G26574,G26575,G26576,G26577,G26578,G26579,G26580,
       G26581,G26582,G26583,G26584,G26585,G26586,G26587,G26588,G26589,G26590,G26591,G26592,G26593,G26594,G26595,G26596,G26597,G26598,G26599,G26600,
       G26601,G26602,G26603,G26604,G26605,G26606,G26607,G26608,G26609,G26610,G26611,G26612,G26613,G26614,G26615,G26616,G26617,G26618,G26619,G26620,
       G26621,G26622,G26623,G26624,G26625,G26626,G26627,G26628,G26629,G26630,G26631,G26632,G26633,G26634,G26635,G26636,G26637,G26638,G26639,G26640,
       G26641,G26642,G26643,G26644,G26645,G26646,G26647,G26648,G26649,G26650,G26651,G26652,G26653,G26654,G26655,G26656,G26657,G26658,G26659,G26660,
       G26661,G26662,G26663,G26664,G26665,G26666,G26667,G26668,G26669,G26670,G26671,G26672,G26673,G26674,G26675,G26676,G26677,G26678,G26679,G26680,
       G26681,G26682,G26683,G26684,G26685,G26686,G26687,G26688,G26689,G26690,G26691,G26692,G26693,G26694,G26695,G26696,G26697,G26698,G26699,G26700,
       G26701,G26702,G26703,G26704,G26705,G26706,G26707,G26708,G26709,G26710,G26711,G26712,G26713,G26714,G26715,G26716,G26717,G26718,G26719,G26720,
       G26721,G26722,G26723,G26724,G26725,G26726,G26727,G26728,G26729,G26730,G26731,G26732,G26733,G26734,G26735,G26736,G26737,G26738,G26739,G26740,
       G26741,G26742,G26743,G26744,G26745,G26746,G26747,G26748,G26749,G26750,G26751,G26752,G26753,G26754,G26755,G26756,G26757,G26758,G26759,G26760,
       G26761,G26762,G26763,G26764,G26765,G26766,G26767,G26768,G26769,G26770,G26771,G26772,G26773,G26774,G26775,G26776,G26777,G26778,G26779,G26780,
       G26781,G26782,G26783,G26784,G26785,G26786,G26787,G26788,G26789,G26790,G26791,G26792,G26793,G26794,G26795,G26796,G26797,G26798,G26799,G26800,
       G26801,G26802,G26803,G26804,G26805,G26806,G26807,G26808,G26809,G26810,G26811,G26812,G26813,G26814,G26815,G26816,G26817,G26818,G26819,G26820,
       G26821,G26822,G26823,G26824,G26825,G26826,G26827,G26828,G26829,G26830,G26831,G26832,G26833,G26834,G26835,G26836,G26837,G26838,G26839,G26840,
       G26841,G26842,G26843,G26844,G26845,G26846,G26847,G26848,G26849,G26850,G26851,G26852,G26853,G26854,G26855,G26856,G26857,G26858,G26859,G26860,
       G26861,G26862,G26863,G26864,G26865,G26866,G26867,G26868,G26869,G26870,G26871,G26872,G26873,G26874,G26875,G26876,G26877,G26878,G26879,G26880,
       G26881,G26882,G26883,G26884,G26885,G26886,G26887,G26888,G26889,G26890,G26891,G26892,G26893,G26894,G26895,G26896,G26897,G26898,G26899,G26900,
       G26901,G26902,G26903,G26904,G26905,G26906,G26907,G26908,G26909,G26910,G26911,G26912,G26913,G26914,G26915,G26916,G26917,G26918,G26919,G26920,
       G26921,G26922,G26923,G26924,G26925,G26926,G26927,G26928,G26929,G26930,G26931,G26932,G26933,G26934,G26935,G26936,G26937,G26938,G26939,G26940,
       G26941,G26942,G26943,G26944,G26945,G26946,G26947,G26948,G26949,G26950,G26951,G26952,G26953,G26954,G26955,G26956,G26957,G26958,G26959,G26960,
       G26961,G26962,G26963,G26964,G26965,G26966,G26967,G26968,G26969,G26970,G26971,G26972,G26973,G26974,G26975,G26976,G26977,G26978,G26979,G26980,
       G26981,G26982,G26983,G26984,G26985,G26986,G26987,G26988,G26989,G26990,G26991,G26992,G26993,G26994,G26995,G26996,G26997,G26998,G26999,G27000,
       G27001,G27002,G27003,G27004,G27005,G27006,G27007,G27008,G27009,G27010,G27011,G27012,G27013,G27014,G27015,G27016,G27017,G27018,G27019,G27020,
       G27021,G27022,G27023,G27024,G27025,G27026,G27027,G27028,G27029,G27030,G27031,G27032,G27033,G27034,G27035,G27036,G27037,G27038,G27039,G27040,
       G27041,G27042,G27043,G27044,G27045,G27046,G27047,G27048,G27049,G27050,G27051,G27052,G27053,G27054,G27055,G27056,G27057,G27058,G27059,G27060,
       G27061,G27062,G27063,G27064,G27065,G27066,G27067,G27068,G27069,G27070,G27071,G27072,G27073,G27074,G27075,G27076,G27077,G27078,G27079,G27080,
       G27081,G27082,G27083,G27084,G27085,G27086,G27087,G27088,G27089,G27090,G27091,G27092,G27093,G27094,G27095,G27096,G27097,G27098,G27099,G27100,
       G27101,G27102,G27103,G27104,G27105,G27106,G27107,G27108,G27109,G27110,G27111,G27112,G27113,G27114,G27115,G27116,G27117,G27118,G27119,G27120,
       G27121,G27122,G27123,G27124,G27125,G27126,G27127,G27128,G27129,G27130,G27131,G27132,G27133,G27134,G27135,G27136,G27137,G27138,G27139,G27140,
       G27141,G27142,G27143,G27144,G27145,G27146,G27147,G27148,G27149,G27150,G27151,G27152,G27153,G27154,G27155,G27156,G27157,G27158,G27159,G27160,
       G27161,G27162,G27163,G27164,G27165,G27166,G27167,G27168,G27169,G27170,G27171,G27172,G27173,G27174,G27175,G27176,G27177,G27178,G27179,G27180,
       G27181,G27182,G27183,G27184,G27185,G27186,G27187,G27188,G27189,G27190,G27191,G27192,G27193,G27194,G27195,G27196,G27197,G27198,G27199,G27200,
       G27201,G27202,G27203,G27204,G27205,G27206,G27207,G27208,G27209,G27210,G27211,G27212,G27213,G27214,G27215,G27216,G27217,G27218,G27219,G27220,
       G27221,G27222,G27223,G27224,G27225,G27226,G27227,G27228,G27229,G27230,G27231,G27232,G27233,G27234,G27235,G27236,G27237,G27238,G27239,G27240,
       G27241,G27242,G27243,G27244,G27245,G27246,G27247,G27248,G27249,G27250,G27251,G27252,G27253,G27254,G27255,G27256,G27257,G27258,G27259,G27260,
       G27261,G27262,G27263,G27264,G27265,G27266,G27267,G27268,G27269,G27270,G27271,G27272,G27273,G27274,G27275,G27276,G27277,G27278,G27279,G27280,
       G27281,G27282,G27283,G27284,G27285,G27286,G27287,G27288,G27289,G27290,G27291,G27292,G27293,G27294,G27295,G27296,G27297,G27298,G27299,G27300,
       G27301,G27302,G27303,G27304,G27305,G27306,G27307,G27308,G27309,G27310,G27311,G27312,G27313,G27314,G27315,G27316,G27317,G27318,G27319,G27320,
       G27321,G27322,G27323,G27324,G27325,G27326,G27327,G27328,G27329,G27330,G27331,G27332,G27333,G27334,G27335,G27336,G27337,G27338,G27339,G27340,
       G27341,G27342,G27343,G27344,G27345,G27346,G27347,G27348,G27349,G27350,G27351,G27352,G27353,G27354,G27355,G27356,G27357,G27358,G27359,G27360,
       G27361,G27362,G27363,G27364,G27365,G27366,G27367,G27368,G27369,G27370,G27371,G27372,G27373,G27374,G27375,G27376,G27377,G27378,G27379,G27380,
       G27381,G27382,G27383,G27384,G27385,G27386,G27387,G27388,G27389,G27390,G27391,G27392,G27393,G27394,G27395,G27396,G27397,G27398,G27399,G27400,
       G27401,G27402,G27403,G27404,G27405,G27406,G27407,G27408,G27409,G27410,G27411,G27412,G27413,G27414,G27415,G27416,G27417,G27418,G27419,G27420,
       G27421,G27422,G27423,G27424,G27425,G27426,G27427,G27428,G27429,G27430,G27431,G27432,G27433,G27434,G27435,G27436,G27437,G27438,G27439,G27440,
       G27441,G27442,G27443,G27444,G27445,G27446,G27447,G27448,G27449,G27450,G27451,G27452,G27453,G27454,G27455,G27456,G27457,G27458,G27459,G27460,
       G27461,G27462,G27463,G27464,G27465,G27466,G27467,G27468,G27469,G27470,G27471,G27472,G27473,G27474,G27475,G27476,G27477,G27478,G27479,G27480,
       G27481,G27482,G27483,G27484,G27485,G27486,G27487,G27488,G27489,G27490,G27491,G27492,G27493,G27494,G27495,G27496,G27497,G27498,G27499,G27500,
       G27501,G27502,G27503,G27504,G27505,G27506,G27507,G27508,G27509,G27510,G27511,G27512,G27513,G27514,G27515,G27516,G27517,G27518,G27519,G27520,
       G27521,G27522,G27523,G27524,G27525,G27526,G27527,G27528,G27529,G27530,G27531,G27532,G27533,G27534,G27535,G27536,G27537,G27538,G27539,G27540,
       G27541,G27542,G27543,G27544,G27545,G27546,G27547,G27548,G27549,G27550,G27551,G27552,G27553,G27554,G27555,G27556,G27557,G27558,G27559,G27560,
       G27561,G27562,G27563,G27564,G27565,G27566,G27567,G27568,G27569,G27570,G27571,G27572,G27573,G27574,G27575,G27576,G27577,G27578,G27579,G27580,
       G27581,G27582,G27583,G27584,G27585,G27586,G27587,G27588,G27589,G27590,G27591,G27592,G27593,G27594,G27595,G27596,G27597,G27598,G27599,G27600,
       G27601,G27602,G27603,G27604,G27605,G27606,G27607,G27608,G27609,G27610,G27611,G27612,G27613,G27614,G27615,G27616,G27617,G27618,G27619,G27620,
       G27621,G27622,G27623,G27624,G27625,G27626,G27627,G27628,G27629,G27630,G27631,G27632,G27633,G27634,G27635,G27636,G27637,G27638,G27639,G27640,
       G27641,G27642,G27643,G27644,G27645,G27646,G27647,G27648,G27649,G27650,G27651,G27652,G27653,G27654,G27655,G27656,G27657,G27658,G27659,G27660,
       G27661,G27662,G27663,G27664,G27665,G27666,G27667,G27668,G27669,G27670,G27671,G27672,G27673,G27674,G27675,G27676,G27677,G27678,G27679,G27680,
       G27681,G27682,G27683,G27684,G27685,G27686,G27687,G27688,G27689,G27690,G27691,G27692,G27693,G27694,G27695,G27696,G27697,G27698,G27699,G27700,
       G27701,G27702,G27703,G27704,G27705,G27706,G27707,G27708,G27709,G27710,G27711,G27712,G27713,G27714,G27715,G27716,G27717,G27718,G27719,G27720,
       G27721,G27722,G27723,G27724,G27725,G27726,G27727,G27728,G27729,G27730,G27731,G27732,G27733,G27734,G27735,G27736,G27737,G27738,G27739,G27740,
       G27741,G27742,G27743,G27744,G27745,G27746,G27747,G27748,G27749,G27750,G27751,G27752,G27753,G27754,G27755,G27756,G27757,G27758,G27759,G27760,
       G27761,G27762,G27763,G27764,G27765,G27766,G27767,G27768,G27769,G27770,G27771,G27772,G27773,G27774,G27775,G27776,G27777,G27778,G27779,G27780,
       G27781,G27782,G27783,G27784,G27785,G27786,G27787,G27788,G27789,G27790,G27791,G27792,G27793,G27794,G27795,G27796,G27797,G27798,G27799,G27800,
       G27801,G27802,G27803,G27804,G27805,G27806,G27807,G27808,G27809,G27810,G27811,G27812,G27813,G27814,G27815,G27816,G27817,G27818,G27819,G27820,
       G27821,G27822,G27823,G27824,G27825,G27826,G27827,G27828,G27829,G27830,G27831,G27832,G27833,G27834,G27835,G27836,G27837,G27838,G27839,G27840,
       G27841,G27842,G27843,G27844,G27845,G27846,G27847,G27848,G27849,G27850,G27851,G27852,G27853,G27854,G27855,G27856,G27857,G27858,G27859,G27860,
       G27861,G27862,G27863,G27864,G27865,G27866,G27867,G27868,G27869,G27870,G27871,G27872,G27873,G27874,G27875,G27876,G27877,G27878,G27879,G27880,
       G27881,G27882,G27883,G27884,G27885,G27886,G27887,G27888,G27889,G27890,G27891,G27892,G27893,G27894,G27895,G27896,G27897,G27898,G27899,G27900,
       G27901,G27902,G27903,G27904,G27905,G27906,G27907,G27908,G27909,G27910,G27911,G27912,G27913,G27914,G27915,G27916,G27917,G27918,G27919,G27920,
       G27921,G27922,G27923,G27924,G27925,G27926,G27927,G27928,G27929,G27930,G27931,G27932,G27933,G27934,G27935,G27936,G27937,G27938,G27939,G27940,
       G27941,G27942,G27943,G27944,G27945,G27946,G27947,G27948,G27949,G27950,G27951,G27952,G27953,G27954,G27955,G27956,G27957,G27958,G27959,G27960,
       G27961,G27962,G27963,G27964,G27965,G27966,G27967,G27968,G27969,G27970,G27971,G27972,G27973,G27974,G27975,G27976,G27977,G27978,G27979,G27980,
       G27981,G27982,G27983,G27984,G27985,G27986,G27987,G27988,G27989,G27990,G27991,G27992,G27993,G27994,G27995,G27996,G27997,G27998,G27999,G28000,
       G28001,G28002,G28003,G28004,G28005,G28006,G28007,G28008,G28009,G28010,G28011,G28012,G28013,G28014,G28015,G28016,G28017,G28018,G28019,G28020,
       G28021,G28022,G28023,G28024,G28025,G28026,G28027,G28028,G28029,G28030,G28031,G28032,G28033,G28034,G28035,G28036,G28037,G28038,G28039,G28040,
       G28041,G28042,G28043,G28044,G28045,G28046,G28047,G28048,G28049,G28050,G28051,G28052,G28053,G28054,G28055,G28056,G28057,G28058,G28059,G28060,
       G28061,G28062,G28063,G28064,G28065,G28066,G28067,G28068,G28069,G28070,G28071,G28072,G28073,G28074,G28075,G28076,G28077,G28078,G28079,G28080,
       G28081,G28082,G28083,G28084,G28085,G28086,G28087,G28088,G28089,G28090,G28091,G28092,G28093,G28094,G28095,G28096,G28097,G28098,G28099,G28100,
       G28101,G28102,G28103,G28104,G28105,G28106,G28107,G28108,G28109,G28110,G28111,G28112,G28113,G28114,G28115,G28116,G28117,G28118,G28119,G28120,
       G28121,G28122,G28123,G28124,G28125,G28126,G28127,G28128,G28129,G28130,G28131,G28132,G28133,G28134,G28135,G28136,G28137,G28138,G28139,G28140,
       G28141,G28142,G28143,G28144,G28145,G28146,G28147,G28148,G28149,G28150,G28151,G28152,G28153,G28154,G28155,G28156,G28157,G28158,G28159,G28160,
       G28161,G28162,G28163,G28164,G28165,G28166,G28167,G28168,G28169,G28170,G28171,G28172,G28173,G28174,G28175,G28176,G28177,G28178,G28179,G28180,
       G28181,G28182,G28183,G28184,G28185,G28186,G28187,G28188,G28189,G28190,G28191,G28192,G28193,G28194,G28195,G28196,G28197,G28198,G28199,G28200,
       G28201,G28202,G28203,G28204,G28205,G28206,G28207,G28208,G28209,G28210,G28211,G28212,G28213,G28214,G28215,G28216,G28217,G28218,G28219,G28220,
       G28221,G28222,G28223,G28224,G28225,G28226,G28227,G28228,G28229,G28230,G28231,G28232,G28233,G28234,G28235,G28236,G28237,G28238,G28239,G28240,
       G28241,G28242,G28243,G28244,G28245,G28246,G28247,G28248,G28249,G28250,G28251,G28252,G28253,G28254,G28255,G28256,G28257,G28258,G28259,G28260,
       G28261,G28262,G28263,G28264,G28265,G28266,G28267,G28268,G28269,G28270,G28271,G28272,G28273,G28274,G28275,G28276,G28277,G28278,G28279,G28280,
       G28281,G28282,G28283,G28284,G28285,G28286,G28287,G28288,G28289,G28290,G28291,G28292,G28293,G28294,G28295,G28296,G28297,G28298,G28299,G28300,
       G28301,G28302,G28303,G28304,G28305,G28306,G28307,G28308,G28309,G28310,G28311,G28312,G28313,G28314,G28315,G28316,G28317,G28318,G28319,G28320,
       G28321,G28322,G28323,G28324,G28325,G28326,G28327,G28328,G28329,G28330,G28331,G28332,G28333,G28334,G28335,G28336,G28337,G28338,G28339,G28340,
       G28341,G28342,G28343,G28344,G28345,G28346,G28347,G28348,G28349,G28350,G28351,G28352,G28353,G28354,G28355,G28356,G28357,G28358,G28359,G28360,
       G28361,G28362,G28363,G28364,G28365,G28366,G28367,G28368,G28369,G28370,G28371,G28372,G28373,G28374,G28375,G28376,G28377,G28378,G28379,G28380,
       G28381,G28382,G28383,G28384,G28385,G28386,G28387,G28388,G28389,G28390,G28391,G28392,G28393,G28394,G28395,G28396,G28397,G28398,G28399,G28400,
       G28401,G28402,G28403,G28404,G28405,G28406,G28407,G28408,G28409,G28410,G28411,G28412,G28413,G28414,G28415,G28416,G28417,G28418,G28419,G28420,
       G28421,G28422,G28423,G28424,G28425,G28426,G28427,G28428,G28429,G28430,G28431,G28432,G28433,G28434,G28435,G28436,G28437,G28438,G28439,G28440,
       G28441,G28442,G28443,G28444,G28445,G28446,G28447,G28448,G28449,G28450,G28451,G28452,G28453,G28454,G28455,G28456,G28457,G28458,G28459,G28460,
       G28461,G28462,G28463,G28464,G28465,G28466,G28467,G28468,G28469,G28470,G28471,G28472,G28473,G28474,G28475,G28476,G28477,G28478,G28479,G28480,
       G28481,G28482,G28483,G28484,G28485,G28486,G28487,G28488,G28489,G28490,G28491,G28492,G28493,G28494,G28495,G28496,G28497,G28498,G28499,G28500,
       G28501,G28502,G28503,G28504,G28505,G28506,G28507,G28508,G28509,G28510,G28511,G28512,G28513,G28514,G28515,G28516,G28517,G28518,G28519,G28520,
       G28521,G28522,G28523,G28524,G28525,G28526,G28527,G28528,G28529,G28530,G28531,G28532,G28533,G28534,G28535,G28536,G28537,G28538,G28539,G28540,
       G28541,G28542,G28543,G28544,G28545,G28546,G28547,G28548,G28549,G28550,G28551,G28552,G28553,G28554,G28555,G28556,G28557,G28558,G28559,G28560,
       G28561,G28562,G28563,G28564,G28565,G28566,G28567,G28568,G28569,G28570,G28571,G28572,G28573,G28574,G28575,G28576,G28577,G28578,G28579,G28580,
       G28581,G28582,G28583,G28584,G28585,G28586,G28587,G28588,G28589,G28590,G28591,G28592,G28593,G28594,G28595,G28596,G28597,G28598,G28599,G28600,
       G28601,G28602,G28603,G28604,G28605,G28606,G28607,G28608,G28609,G28610,G28611,G28612,G28613,G28614,G28615,G28616,G28617,G28618,G28619,G28620,
       G28621,G28622,G28623,G28624,G28625,G28626,G28627,G28628,G28629,G28630,G28631,G28632,G28633,G28634,G28635,G28636,G28637,G28638,G28639,G28640,
       G28641,G28642,G28643,G28644,G28645,G28646,G28647,G28648,G28649,G28650,G28651,G28652,G28653,G28654,G28655,G28656,G28657,G28658,G28659,G28660,
       G28661,G28662,G28663,G28664,G28665,G28666,G28667,G28668,G28669,G28670,G28671,G28672,G28673,G28674,G28675,G28676,G28677,G28678,G28679,G28680,
       G28681,G28682,G28683,G28684,G28685,G28686,G28687,G28688,G28689,G28690,G28691,G28692,G28693,G28694,G28695,G28696,G28697,G28698,G28699,G28700,
       G28701,G28702,G28703,G28704,G28705,G28706,G28707,G28708,G28709,G28710,G28711,G28712,G28713,G28714,G28715,G28716,G28717,G28718,G28719,G28720,
       G28721,G28722,G28723,G28724,G28725,G28726,G28727,G28728,G28729,G28730,G28731,G28732,G28733,G28734,G28735,G28736,G28737,G28738,G28739,G28740,
       G28741,G28742,G28743,G28744,G28745,G28746,G28747,G28748,G28749,G28750,G28751,G28752,G28753,G28754,G28755,G28756,G28757,G28758,G28759,G28760,
       G28761,G28762,G28763,G28764,G28765,G28766,G28767,G28768,G28769,G28770,G28771,G28772,G28773,G28774,G28775,G28776,G28777,G28778,G28779,G28780,
       G28781,G28782,G28783,G28784,G28785,G28786,G28787,G28788,G28789,G28790,G28791,G28792,G28793,G28794,G28795,G28796,G28797,G28798,G28799,G28800,
       G28801,G28802,G28803,G28804,G28805,G28806,G28807,G28808,G28809,G28810,G28811,G28812,G28813,G28814,G28815,G28816,G28817,G28818,G28819,G28820,
       G28821,G28822,G28823,G28824,G28825,G28826,G28827,G28828,G28829,G28830,G28831,G28832,G28833,G28834,G28835,G28836,G28837,G28838,G28839,G28840,
       G28841,G28842,G28843,G28844,G28845,G28846,G28847,G28848,G28849,G28850,G28851,G28852,G28853,G28854,G28855,G28856,G28857,G28858,G28859,G28860,
       G28861,G28862,G28863,G28864,G28865,G28866,G28867,G28868,G28869,G28870,G28871,G28872,G28873,G28874,G28875,G28876,G28877,G28878,G28879,G28880,
       G28881,G28882,G28883,G28884,G28885,G28886,G28887,G28888,G28889,G28890,G28891,G28892,G28893,G28894,G28895,G28896,G28897,G28898,G28899,G28900,
       G28901,G28902,G28903,G28904,G28905,G28906,G28907,G28908,G28909,G28910,G28911,G28912,G28913,G28914,G28915,G28916,G28917,G28918,G28919,G28920,
       G28921,G28922,G28923,G28924,G28925,G28926,G28927,G28928,G28929,G28930,G28931,G28932,G28933,G28934,G28935,G28936,G28937,G28938,G28939,G28940,
       G28941,G28942,G28943,G28944,G28945,G28946,G28947,G28948,G28949,G28950,G28951,G28952,G28953,G28954,G28955,G28956,G28957,G28958,G28959,G28960,
       G28961,G28962,G28963,G28964,G28965,G28966,G28967,G28968,G28969,G28970,G28971,G28972,G28973,G28974,G28975,G28976,G28977,G28978,G28979,G28980,
       G28981,G28982,G28983,G28984,G28985,G28986,G28987,G28988,G28989,G28990,G28991,G28992,G28993,G28994,G28995,G28996,G28997,G28998,G28999,G29000,
       G29001,G29002,G29003,G29004,G29005,G29006,G29007,G29008,G29009,G29010,G29011,G29012,G29013,G29014,G29015,G29016,G29017,G29018,G29019,G29020,
       G29021,G29022,G29023,G29024,G29025,G29026,G29027,G29028,G29029,G29030,G29031,G29032,G29033,G29034,G29035,G29036,G29037,G29038,G29039,G29040,
       G29041,G29042,G29043,G29044,G29045,G29046,G29047,G29048,G29049,G29050,G29051,G29052,G29053,G29054,G29055,G29056,G29057,G29058,G29059,G29060,
       G29061,G29062,G29063,G29064,G29065,G29066,G29067,G29068,G29069,G29070,G29071,G29072,G29073,G29074,G29075,G29076,G29077,G29078,G29079,G29080,
       G29081,G29082,G29083,G29084,G29085,G29086,G29087,G29088,G29089,G29090,G29091,G29092,G29093,G29094,G29095,G29096,G29097,G29098,G29099,G29100,
       G29101,G29102,G29103,G29104,G29105,G29106,G29107,G29108,G29109,G29110,G29111,G29112,G29113,G29114,G29115,G29116,G29117,G29118,G29119,G29120,
       G29121,G29122,G29123,G29124,G29125,G29126,G29127,G29128,G29129,G29130,G29131,G29132,G29133,G29134,G29135,G29136,G29137,G29138,G29139,G29140,
       G29141,G29142,G29143,G29144,G29145,G29146,G29147,G29148,G29149,G29150,G29151,G29152,G29153,G29154,G29155,G29156,G29157,G29158,G29159,G29160,
       G29161,G29162,G29163,G29164,G29165,G29166,G29167,G29168,G29169,G29170,G29171,G29172,G29173,G29174,G29175,G29176,G29177,G29178,G29179,G29180,
       G29181,G29182,G29183,G29184,G29185,G29186,G29187,G29188,G29189,G29190,G29191,G29192,G29193,G29194,G29195,G29196,G29197,G29198,G29199,G29200,
       G29201,G29202,G29203,G29204,G29205,G29206,G29207,G29208,G29209,G29210,G29211,G29212,G29213,G29214,G29215,G29216,G29217,G29218,G29219,G29220,
       G29221,G29222,G29223,G29224,G29225,G29226,G29227,G29228,G29229,G29230,G29231,G29232,G29233,G29234,G29235,G29236,G29237,G29238,G29239,G29240,
       G29241,G29242,G29243,G29244,G29245,G29246,G29247,G29248,G29249,G29250,G29251,G29252,G29253,G29254,G29255,G29256,G29257,G29258,G29259,G29260,
       G29261,G29262,G29263,G29264,G29265,G29266,G29267,G29268,G29269,G29270,G29271,G29272,G29273,G29274,G29275,G29276,G29277,G29278,G29279,G29280,
       G29281,G29282,G29283,G29284,G29285,G29286,G29287,G29288,G29289,G29290,G29291,G29292,G29293,G29294,G29295,G29296,G29297,G29298,G29299,G29300,
       G29301,G29302,G29303,G29304,G29305,G29306,G29307,G29308,G29309,G29310,G29311,G29312,G29313,G29314,G29315,G29316,G29317,G29318,G29319,G29320,
       G29321,G29322,G29323,G29324,G29325,G29326,G29327,G29328,G29329,G29330,G29331,G29332,G29333,G29334,G29335,G29336,G29337,G29338,G29339,G29340,
       G29341,G29342,G29343,G29344,G29345,G29346,G29347,G29348,G29349,G29350,G29351,G29352,G29353,G29354,G29355,G29356,G29357,G29358,G29359,G29360,
       G29361,G29362,G29363,G29364,G29365,G29366,G29367,G29368,G29369,G29370,G29371,G29372,G29373,G29374,G29375,G29376,G29377,G29378,G29379,G29380,
       G29381,G29382,G29383,G29384,G29385,G29386,G29387,G29388,G29389,G29390,G29391,G29392,G29393,G29394,G29395,G29396,G29397,G29398,G29399,G29400,
       G29401,G29402,G29403,G29404,G29405,G29406,G29407,G29408,G29409,G29410,G29411,G29412,G29413,G29414,G29415,G29416,G29417,G29418,G29419,G29420,
       G29421,G29422,G29423,G29424,G29425,G29426,G29427,G29428,G29429,G29430,G29431,G29432,G29433,G29434,G29435,G29436,G29437,G29438,G29439,G29440,
       G29441,G29442,G29443,G29444,G29445,G29446,G29447,G29448,G29449,G29450,G29451,G29452,G29453,G29454,G29455,G29456,G29457,G29458,G29459,G29460,
       G29461,G29462,G29463,G29464,G29465,G29466,G29467,G29468,G29469,G29470,G29471,G29472,G29473,G29474,G29475,G29476,G29477,G29478,G29479,G29480,
       G29481,G29482,G29483,G29484,G29485,G29486,G29487,G29488,G29489,G29490,G29491,G29492,G29493,G29494,G29495,G29496,G29497,G29498,G29499,G29500,
       G29501,G29502,G29503,G29504,G29505,G29506,G29507,G29508,G29509,G29510,G29511,G29512,G29513,G29514,G29515,G29516,G29517,G29518,G29519,G29520,
       G29521,G29522,G29523,G29524,G29525,G29526,G29527,G29528,G29529,G29530,G29531,G29532,G29533,G29534,G29535,G29536,G29537,G29538,G29539,G29540,
       G29541,G29542,G29543,G29544,G29545,G29546,G29547,G29548,G29549,G29550,G29551,G29552,G29553,G29554,G29555,G29556,G29557,G29558,G29559,G29560,
       G29561,G29562,G29563,G29564,G29565,G29566,G29567,G29568,G29569,G29570,G29571,G29572,G29573,G29574,G29575,G29576,G29577,G29578,G29579,G29580,
       G29581,G29582,G29583,G29584,G29585,G29586,G29587,G29588,G29589,G29590,G29591,G29592,G29593,G29594,G29595,G29596,G29597,G29598,G29599,G29600,
       G29601,G29602,G29603,G29604,G29605,G29606,G29607,G29608,G29609,G29610,G29611,G29612,G29613,G29614,G29615,G29616,G29617,G29618,G29619,G29620,
       G29621,G29622,G29623,G29624,G29625,G29626,G29627,G29628,G29629,G29630,G29631,G29632,G29633,G29634,G29635,G29636,G29637,G29638,G29639,G29640,
       G29641,G29642,G29643,G29644,G29645,G29646,G29647,G29648,G29649,G29650,G29651,G29652,G29653,G29654,G29655,G29656,G29657,G29658,G29659,G29660,
       G29661,G29662,G29663,G29664,G29665,G29666,G29667,G29668,G29669,G29670,G29671,G29672,G29673,G29674,G29675,G29676,G29677,G29678,G29679,G29680,
       G29681,G29682,G29683,G29684,G29685,G29686,G29687,G29688,G29689,G29690,G29691,G29692,G29693,G29694,G29695,G29696,G29697,G29698,G29699,G29700,
       G29701,G29702,G29703,G29704,G29705,G29706,G29707,G29708,G29709,G29710,G29711,G29712,G29713,G29714,G29715,G29716,G29717,G29718,G29719,G29720,
       G29721,G29722,G29723,G29724,G29725,G29726,G29727,G29728,G29729,G29730,G29731,G29732,G29733,G29734,G29735,G29736,G29737,G29738,G29739,G29740,
       G29741,G29742,G29743,G29744,G29745,G29746,G29747,G29748,G29749,G29750,G29751,G29752,G29753,G29754,G29755,G29756,G29757,G29758,G29759,G29760,
       G29761,G29762,G29763,G29764,G29765,G29766,G29767,G29768,G29769,G29770,G29771,G29772,G29773,G29774,G29775,G29776,G29777,G29778,G29779,G29780,
       G29781,G29782,G29783,G29784,G29785,G29786,G29787,G29788,G29789,G29790,G29791,G29792,G29793,G29794,G29795,G29796,G29797,G29798,G29799,G29800,
       G29801,G29802,G29803,G29804,G29805,G29806,G29807,G29808,G29809,G29810,G29811,G29812,G29813,G29814,G29815,G29816,G29817,G29818,G29819,G29820,
       G29821,G29822,G29823,G29824,G29825,G29826,G29827,G29828,G29829,G29830,G29831,G29832,G29833,G29834,G29835,G29836,G29837,G29838,G29839,G29840,
       G29841,G29842,G29843,G29844,G29845,G29846,G29847,G29848,G29849,G29850,G29851,G29852,G29853,G29854,G29855,G29856,G29857,G29858,G29859,G29860,
       G29861,G29862,G29863,G29864,G29865,G29866,G29867,G29868,G29869,G29870,G29871,G29872,G29873,G29874,G29875,G29876,G29877,G29878,G29879,G29880,
       G29881,G29882,G29883,G29884,G29885,G29886,G29887,G29888,G29889,G29890,G29891,G29892,G29893,G29894,G29895,G29896,G29897,G29898,G29899,G29900,
       G29901,G29902,G29903,G29904,G29905,G29906,G29907,G29908,G29909,G29910,G29911,G29912,G29913,G29914,G29915,G29916,G29917,G29918,G29919,G29920,
       G29921,G29922,G29923,G29924,G29925,G29926,G29927,G29928,G29929,G29930,G29931,G29932,G29933,G29934,G29935,G29936,G29937,G29938,G29939,G29940,
       G29941,G29942,G29943,G29944,G29945,G29946,G29947,G29948,G29949,G29950,G29951,G29952,G29953,G29954,G29955,G29956,G29957,G29958,G29959,G29960,
       G29961,G29962,G29963,G29964,G29965,G29966,G29967,G29968,G29969,G29970,G29971,G29972,G29973,G29974,G29975,G29976,G29977,G29978,G29979,G29980,
       G29981,G29982,G29983,G29984,G29985,G29986,G29987,G29988,G29989,G29990,G29991,G29992,G29993,G29994,G29995,G29996,G29997,G29998,G29999,G30000,
       G30001,G30002,G30003,G30004,G30005,G30006,G30007,G30008,G30009,G30010,G30011,G30012,G30013,G30014,G30015,G30016,G30017,G30018,G30019,G30020,
       G30021,G30022,G30023,G30024,G30025,G30026,G30027,G30028,G30029,G30030,G30031,G30032,G30033,G30034,G30035,G30036,G30037,G30038,G30039,G30040,
       G30041,G30042,G30043,G30044,G30045,G30046,G30047,G30048,G30049,G30050,G30051,G30052,G30053,G30054,G30055,G30056,G30057,G30058,G30059,G30060,
       G30061,G30062,G30063,G30064,G30065,G30066,G30067,G30068,G30069,G30070,G30071,G30072,G30073,G30074,G30075,G30076,G30077,G30078,G30079,G30080,
       G30081,G30082,G30083,G30084,G30085,G30086,G30087,G30088,G30089,G30090,G30091,G30092,G30093,G30094,G30095,G30096,G30097,G30098,G30099,G30100,
       G30101,G30102,G30103,G30104,G30105,G30106,G30107,G30108,G30109,G30110,G30111,G30112,G30113,G30114,G30115,G30116,G30117,G30118,G30119,G30120,
       G30121,G30122,G30123,G30124,G30125,G30126,G30127,G30128,G30129,G30130,G30131,G30132,G30133,G30134,G30135,G30136,G30137,G30138,G30139,G30140,
       G30141,G30142,G30143,G30144,G30145,G30146,G30147,G30148,G30149,G30150,G30151,G30152,G30153,G30154,G30155,G30156,G30157,G30158,G30159,G30160,
       G30161,G30162,G30163,G30164,G30165,G30166,G30167,G30168,G30169,G30170,G30171,G30172,G30173,G30174,G30175,G30176,G30177,G30178,G30179,G30180,
       G30181,G30182,G30183,G30184,G30185,G30186,G30187,G30188,G30189,G30190,G30191,G30192,G30193,G30194,G30195,G30196,G30197,G30198,G30199,G30200,
       G30201,G30202,G30203,G30204,G30205,G30206,G30207,G30208,G30209,G30210,G30211,G30212,G30213,G30214,G30215,G30216,G30217,G30218,G30219,G30220,
       G30221,G30222,G30223,G30224,G30225,G30226,G30227,G30228,G30229,G30230,G30231,G30232,G30233,G30234,G30235,G30236,G30237,G30238,G30239,G30240,
       G30241,G30242,G30243,G30244,G30245,G30246,G30247,G30248,G30249,G30250,G30251,G30252,G30253,G30254,G30255,G30256,G30257,G30258,G30259,G30260,
       G30261,G30262,G30263,G30264,G30265,G30266,G30267,G30268,G30269,G30270,G30271,G30272,G30273,G30274,G30275,G30276,G30277,G30278,G30279,G30280,
       G30281,G30282,G30283,G30284,G30285,G30286,G30287,G30288,G30289,G30290,G30291,G30292,G30293,G30294,G30295,G30296,G30297,G30298,G30299,G30300,
       G30301,G30302,G30303,G30304,G30305,G30306,G30307,G30308,G30309,G30310,G30311,G30312,G30313,G30314,G30315,G30316,G30317,G30318,G30319,G30320,
       G30321,G30322,G30323,G30324,G30325,G30326,G30327,G30328,G30329,G30330,G30331,G30332,G30333,G30334,G30335,G30336,G30337,G30338,G30339,G30340,
       G30341,G30342,G30343,G30344,G30345,G30346,G30347,G30348,G30349,G30350,G30351,G30352,G30353,G30354,G30355,G30356,G30357,G30358,G30359,G30360,
       G30361,G30362,G30363,G30364,G30365,G30366,G30367,G30368,G30369,G30370,G30371,G30372,G30373,G30374,G30375,G30376,G30377,G30378,G30379,G30380,
       G30381,G30382,G30383,G30384,G30385,G30386,G30387,G30388,G30389,G30390,G30391,G30392,G30393,G30394,G30395,G30396,G30397,G30398,G30399,G30400,
       G30401,G30402,G30403,G30404,G30405,G30406,G30407,G30408,G30409,G30410,G30411,G30412,G30413,G30414,G30415,G30416,G30417,G30418,G30419,G30420,
       G30421,G30422,G30423,G30424,G30425,G30426,G30427,G30428,G30429,G30430,G30431,G30432,G30433,G30434,G30435,G30436,G30437,G30438,G30439,G30440,
       G30441,G30442,G30443,G30444,G30445,G30446,G30447,G30448,G30449,G30450,G30451,G30452,G30453,G30454,G30455,G30456,G30457,G30458,G30459,G30460,
       G30461,G30462,G30463,G30464,G30465,G30466,G30467,G30468,G30469,G30470,G30471,G30472,G30473,G30474,G30475,G30476,G30477,G30478,G30479,G30480,
       G30481,G30482,G30483,G30484,G30485,G30486,G30487,G30488,G30489,G30490,G30491,G30492,G30493,G30494,G30495,G30496,G30497,G30498,G30499,G30500,
       G30501,G30502,G30503,G30504,G30505,G30506,G30507,G30508,G30509,G30510,G30511,G30512,G30513,G30514,G30515,G30516,G30517,G30518,G30519,G30520,
       G30521,G30522,G30523,G30524,G30525,G30526,G30527,G30528,G30529,G30530,G30531,G30532,G30533,G30534,G30535,G30536,G30537,G30538,G30539,G30540,
       G30541,G30542,G30543,G30544,G30545,G30546,G30547,G30548,G30549,G30550,G30551,G30552,G30553,G30554,G30555,G30556,G30557,G30558,G30559,G30560,
       G30561,G30562,G30563,G30564,G30565,G30566,G30567,G30568,G30569,G30570,G30571,G30572,G30573,G30574,G30575,G30576,G30577,G30578,G30579,G30580,
       G30581,G30582,G30583,G30584,G30585,G30586,G30587,G30588,G30589,G30590,G30591,G30592,G30593,G30594,G30595,G30596,G30597,G30598,G30599,G30600,
       G30601,G30602,G30603,G30604,G30605,G30606,G30607,G30608,G30609,G30610,G30611,G30612,G30613,G30614,G30615,G30616,G30617,G30618,G30619,G30620,
       G30621,G30622,G30623,G30624,G30625,G30626,G30627,G30628,G30629,G30630,G30631,G30632,G30633,G30634,G30635,G30636,G30637,G30638,G30639,G30640,
       G30641,G30642,G30643,G30644,G30645,G30646,G30647,G30648,G30649,G30650,G30651,G30652,G30653,G30654,G30655,G30656,G30657,G30658,G30659,G30660,
       G30661,G30662,G30663,G30664,G30665,G30666,G30667,G30668,G30669,G30670,G30671,G30672,G30673,G30674,G30675,G30676,G30677,G30678,G30679,G30680,
       G30681,G30682,G30683,G30684,G30685,G30686,G30687,G30688,G30689,G30690,G30691,G30692,G30693,G30694,G30695,G30696,G30697,G30698,G30699,G30700,
       G30701,G30702,G30703,G30704,G30705,G30706,G30707,G30708,G30709,G30710,G30711,G30712,G30713,G30714,G30715,G30716,G30717,G30718,G30719,G30720,
       G30721,G30722,G30723,G30724,G30725,G30726,G30727,G30728,G30729,G30730,G30731,G30732,G30733,G30734,G30735,G30736,G30737,G30738,G30739,G30740,
       G30741,G30742,G30743,G30744,G30745,G30746,G30747,G30748,G30749,G30750,G30751,G30752,G30753,G30754,G30755,G30756,G30757,G30758,G30759,G30760,
       G30761,G30762,G30763,G30764,G30765,G30766,G30767,G30768,G30769,G30770,G30771,G30772,G30773,G30774,G30775,G30776,G30777,G30778,G30779,G30780,
       G30781,G30782,G30783,G30784,G30785,G30786,G30787,G30788,G30789,G30790,G30791,G30792,G30793,G30794,G30795,G30796,G30797,G30798,G30799,G30800,
       G30801,G30802,G30803,G30804,G30805,G30806,G30807,G30808,G30809,G30810,G30811,G30812,G30813,G30814,G30815,G30816,G30817,G30818,G30819,G30820,
       G30821,G30822,G30823,G30824,G30825,G30826,G30827,G30828,G30829,G30830,G30831,G30832,G30833,G30834,G30835,G30836,G30837,G30838,G30839,G30840,
       G30841,G30842,G30843,G30844,G30845,G30846,G30847,G30848,G30849,G30850,G30851,G30852,G30853,G30854,G30855,G30856,G30857,G30858,G30859,G30860,
       G30861,G30862,G30863,G30864,G30865,G30866,G30867,G30868,G30869,G30870,G30871,G30872,G30873,G30874,G30875,G30876,G30877,G30878,G30879,G30880,
       G30881,G30882,G30883,G30884,G30885,G30886,G30887,G30888,G30889,G30890,G30891,G30892,G30893,G30894,G30895,G30896,G30897,G30898,G30899,G30900,
       G30901,G30902,G30903,G30904,G30905,G30906,G30907,G30908,G30909,G30910,G30911,G30912,G30913,G30914,G30915,G30916,G30917,G30918,G30919,G30920,
       G30921,G30922,G30923,G30924,G30925,G30926,G30927,G30928,G30929,G30930,G30931,G30932,G30933,G30934,G30935,G30936,G30937,G30938,G30939,G30940,
       G30941,G30942,G30943,G30944,G30945,G30946,G30947,G30948,G30949,G30950,G30951,G30952,G30953,G30954,G30955,G30956,G30957,G30958,G30959,G30960,
       G30961,G30962,G30963,G30964,G30965,G30966,G30967,G30968,G30969,G30970,G30971,G30972,G30973,G30974,G30975,G30976,G30977,G30978,G30979,G30980,
       G30981,G30982,G30983,G30984,G30985,G30986,G30987,G30988,G30989,G30990,G30991,G30992,G30993,G30994,G30995,G30996,G30997,G30998,G30999,G31000,
       G31001,G31002,G31003,G31004,G31005,G31006,G31007,G31008,G31009,G31010,G31011,G31012,G31013,G31014,G31015,G31016,G31017,G31018,G31019,G31020,
       G31021,G31022,G31023,G31024,G31025,G31026,G31027,G31028,G31029,G31030,G31031,G31032,G31033,G31034,G31035,G31036,G31037,G31038,G31039,G31040,
       G31041,G31042,G31043,G31044,G31045,G31046,G31047,G31048,G31049,G31050,G31051,G31052,G31053,G31054,G31055,G31056,G31057,G31058,G31059,G31060,
       G31061,G31062,G31063,G31064,G31065,G31066,G31067,G31068,G31069,G31070,G31071,G31072,G31073,G31074,G31075,G31076,G31077,G31078,G31079,G31080,
       G31081,G31082,G31083,G31084,G31085,G31086,G31087,G31088,G31089,G31090,G31091,G31092,G31093,G31094,G31095,G31096,G31097,G31098,G31099,G31100,
       G31101,G31102,G31103,G31104,G31105,G31106,G31107,G31108,G31109,G31110,G31111,G31112,G31113,G31114,G31115,G31116,G31117,G31118,G31119,G31120,
       G31121,G31122,G31123,G31124,G31125,G31126,G31127,G31128,G31129,G31130,G31131,G31132,G31133,G31134,G31135,G31136,G31137,G31138,G31139,G31140,
       G31141,G31142,G31143,G31144,G31145,G31146,G31147,G31148,G31149,G31150,G31151,G31152,G31153,G31154,G31155,G31156,G31157,G31158,G31159,G31160,
       G31161,G31162,G31163,G31164,G31165,G31166,G31167,G31168,G31169,G31170,G31171,G31172,G31173,G31174,G31175,G31176,G31177,G31178,G31179,G31180,
       G31181,G31182,G31183,G31184,G31185,G31186,G31187,G31188,G31189,G31190,G31191,G31192,G31193,G31194,G31195,G31196,G31197,G31198,G31199,G31200,
       G31201,G31202,G31203,G31204,G31205,G31206,G31207,G31208,G31209,G31210,G31211,G31212,G31213,G31214,G31215,G31216,G31217,G31218,G31219,G31220,
       G31221,G31222,G31223,G31224,G31225,G31226,G31227,G31228,G31229,G31230,G31231,G31232,G31233,G31234,G31235,G31236,G31237,G31238,G31239,G31240,
       G31241,G31242,G31243,G31244,G31245,G31246,G31247,G31248,G31249,G31250,G31251,G31252,G31253,G31254,G31255,G31256,G31257,G31258,G31259,G31260,
       G31261,G31262,G31263,G31264,G31265,G31266,G31267,G31268,G31269,G31270,G31271,G31272,G31273,G31274,G31275,G31276,G31277,G31278,G31279,G31280,
       G31281,G31282,G31283,G31284,G31285,G31286,G31287,G31288,G31289,G31290,G31291,G31292,G31293,G31294,G31295,G31296,G31297,G31298,G31299,G31300,
       G31301,G31302,G31303,G31304,G31305,G31306,G31307,G31308,G31309,G31310,G31311,G31312,G31313,G31314,G31315,G31316,G31317,G31318,G31319,G31320,
       G31321,G31322,G31323,G31324,G31325,G31326,G31327,G31328,G31329,G31330,G31331,G31332,G31333,G31334,G31335,G31336,G31337,G31338,G31339,G31340,
       G31341,G31342,G31343,G31344,G31345,G31346,G31347,G31348,G31349,G31350,G31351,G31352,G31353,G31354,G31355,G31356,G31357,G31358,G31359,G31360,
       G31361,G31362,G31363,G31364,G31365,G31366,G31367,G31368,G31369,G31370,G31371,G31372,G31373,G31374,G31375,G31376,G31377,G31378,G31379,G31380,
       G31381,G31382,G31383,G31384,G31385,G31386,G31387,G31388,G31389,G31390,G31391,G31392,G31393,G31394,G31395,G31396,G31397,G31398,G31399,G31400,
       G31401,G31402,G31403,G31404,G31405,G31406,G31407,G31408,G31409,G31410,G31411,G31412,G31413,G31414,G31415,G31416,G31417,G31418,G31419,G31420,
       G31421,G31422,G31423,G31424,G31425,G31426,G31427,G31428,G31429,G31430,G31431,G31432,G31433,G31434,G31435,G31436,G31437,G31438,G31439,G31440,
       G31441,G31442,G31443,G31444,G31445,G31446,G31447,G31448,G31449,G31450,G31451,G31452,G31453,G31454,G31455,G31456,G31457,G31458,G31459,G31460,
       G31461,G31462,G31463,G31464,G31465,G31466,G31467,G31468,G31469,G31470,G31471,G31472,G31473,G31474,G31475,G31476,G31477,G31478,G31479,G31480,
       G31481,G31482,G31483,G31484,G31485,G31486,G31487,G31488,G31489,G31490,G31491,G31492,G31493,G31494,G31495,G31496,G31497,G31498,G31499,G31500,
       G31501,G31502,G31503,G31504,G31505,G31506,G31507,G31508,G31509,G31510,G31511,G31512,G31513,G31514,G31515,G31516,G31517,G31518,G31519,G31520,
       G31521,G31522,G31523,G31524,G31525,G31526,G31527,G31528,G31529,G31530,G31531,G31532,G31533,G31534,G31535,G31536,G31537,G31538,G31539,G31540,
       G31541,G31542,G31543,G31544,G31545,G31546,G31547,G31548,G31549,G31550,G31551,G31552,G31553,G31554,G31555,G31556,G31557,G31558,G31559,G31560,
       G31561,G31562,G31563,G31564,G31565,G31566,G31567,G31568,G31569,G31570,G31571,G31572,G31573,G31574,G31575,G31576,G31577,G31578,G31579,G31580,
       G31581,G31582,G31583,G31584,G31585,G31586,G31587,G31588,G31589,G31590,G31591,G31592,G31593,G31594,G31595,G31596,G31597,G31598,G31599,G31600,
       G31601,G31602,G31603,G31604,G31605,G31606,G31607,G31608,G31609,G31610,G31611,G31612,G31613,G31614,G31615,G31616,G31617,G31618,G31619,G31620,
       G31621,G31622,G31623,G31624,G31625,G31626,G31627,G31628,G31629,G31630,G31631,G31632,G31633,G31634,G31635,G31636,G31637,G31638,G31639,G31640,
       G31641,G31642,G31643,G31644,G31645,G31646,G31647,G31648,G31649,G31650,G31651,G31652,G31653,G31654,G31655,G31656,G31657,G31658,G31659,G31660,
       G31661,G31662,G31663,G31664,G31665,G31666,G31667,G31668,G31669,G31670,G31671,G31672,G31673,G31674,G31675,G31676,G31677,G31678,G31679,G31680,
       G31681,G31682,G31683,G31684,G31685,G31686,G31687,G31688,G31689,G31690,G31691,G31692,G31693,G31694,G31695,G31696,G31697,G31698,G31699,G31700,
       G31701,G31702,G31703,G31704,G31705,G31706,G31707,G31708,G31709,G31710,G31711,G31712,G31713,G31714,G31715,G31716,G31717,G31718,G31719,G31720,
       G31721,G31722,G31723,G31724,G31725,G31726,G31727,G31728,G31729,G31730,G31731,G31732,G31733,G31734,G31735,G31736,G31737,G31738,G31739,G31740,
       G31741,G31742,G31743,G31744,G31745,G31746,G31747,G31748,G31749,G31750,G31751,G31752,G31753,G31754,G31755,G31756,G31757,G31758,G31759,G31760,
       G31761,G31762,G31763,G31764,G31765,G31766,G31767,G31768,G31769,G31770,G31771,G31772,G31773,G31774,G31775,G31776,G31777,G31778,G31779,G31780,
       G31781,G31782,G31783,G31784,G31785,G31786,G31787,G31788,G31789,G31790,G31791,G31792,G31793,G31794,G31795,G31796,G31797,G31798,G31799,G31800,
       G31801,G31802,G31803,G31804,G31805,G31806,G31807,G31808,G31809,G31810,G31811,G31812,G31813,G31814,G31815,G31816,G31817,G31818,G31819,G31820,
       G31821,G31822,G31823,G31824,G31825,G31826,G31827,G31828,G31829,G31830,G31831,G31832,G31833,G31834,G31835,G31836,G31837,G31838,G31839,G31840,
       G31841,G31842,G31843,G31844,G31845,G31846,G31847,G31848,G31849,G31850,G31851,G31852,G31853,G31854,G31855,G31856,G31857,G31858,G31859,G31860,
       G31861,G31862,G31863,G31864,G31865,G31866,G31867,G31868,G31869,G31870,G31871,G31872,G31873,G31874,G31875,G31876,G31877,G31878,G31879,G31880,
       G31881,G31882,G31883,G31884,G31885,G31886,G31887,G31888,G31889,G31890,G31891,G31892,G31893,G31894,G31895,G31896,G31897,G31898,G31899,G31900,
       G31901,G31902,G31903,G31904,G31905,G31906,G31907,G31908,G31909,G31910,G31911,G31912,G31913,G31914,G31915,G31916,G31917,G31918,G31919,G31920,
       G31921,G31922,G31923,G31924,G31925,G31926,G31927,G31928,G31929,G31930,G31931,G31932,G31933,G31934,G31935,G31936,G31937,G31938,G31939,G31940,
       G31941,G31942,G31943,G31944,G31945,G31946,G31947,G31948,G31949,G31950,G31951,G31952,G31953,G31954,G31955,G31956,G31957,G31958,G31959,G31960,
       G31961,G31962,G31963,G31964,G31965,G31966,G31967,G31968,G31969,G31970,G31971,G31972,G31973,G31974,G31975,G31976,G31977,G31978,G31979,G31980,
       G31981,G31982,G31983,G31984,G31985,G31986,G31987,G31988,G31989,G31990,G31991,G31992,G31993,G31994,G31995,G31996,G31997,G31998,G31999,G32000,
       G32001,G32002,G32003,G32004,G32005,G32006,G32007,G32008,G32009,G32010,G32011,G32012,G32013,G32014,G32015,G32016,G32017,G32018,G32019,G32020,
       G32021,G32022,G32023,G32024,G32025,G32026,G32027,G32028,G32029,G32030,G32031,G32032,G32033,G32034,G32035,G32036,G32037,G32038,G32039,G32040,
       G32041,G32042,G32043,G32044,G32045,G32046,G32047,G32048,G32049,G32050,G32051,G32052,G32053,G32054,G32055,G32056,G32057,G32058,G32059,G32060,
       G32061,G32062,G32063,G32064,G32065,G32066,G32067,G32068,G32069,G32070,G32071,G32072,G32073,G32074,G32075,G32076,G32077,G32078,G32079,G32080,
       G32081,G32082,G32083,G32084,G32085,G32086,G32087,G32088,G32089,G32090,G32091,G32092,G32093,G32094,G32095,G32096,G32097,G32098,G32099,G32100,
       G32101,G32102,G32103,G32104,G32105,G32106,G32107,G32108,G32109,G32110,G32111,G32112,G32113,G32114,G32115,G32116,G32117,G32118,G32119,G32120,
       G32121,G32122,G32123,G32124,G32125,G32126,G32127,G32128,G32129,G32130,G32131,G32132,G32133,G32134,G32135,G32136,G32137,G32138,G32139,G32140,
       G32141,G32142,G32143,G32144,G32145,G32146,G32147,G32148,G32149,G32150,G32151,G32152,G32153,G32154,G32155,G32156,G32157,G32158,G32159,G32160,
       G32161,G32162,G32163,G32164,G32165,G32166,G32167,G32168,G32169,G32170,G32171,G32172,G32173,G32174,G32175,G32176,G32177,G32178,G32179,G32180,
       G32181,G32182,G32183,G32184,G32185,G32186,G32187,G32188,G32189,G32190,G32191,G32192,G32193,G32194,G32195,G32196,G32197,G32198,G32199,G32200,
       G32201,G32202,G32203,G32204,G32205,G32206,G32207,G32208,G32209,G32210,G32211,G32212,G32213,G32214,G32215,G32216,G32217,G32218,G32219,G32220,
       G32221,G32222,G32223,G32224,G32225,G32226,G32227,G32228,G32229,G32230,G32231,G32232,G32233,G32234,G32235,G32236,G32237,G32238,G32239,G32240,
       G32241,G32242,G32243,G32244,G32245,G32246,G32247,G32248,G32249,G32250,G32251,G32252,G32253,G32254,G32255,G32256,G32257,G32258,G32259,G32260,
       G32261,G32262,G32263,G32264,G32265,G32266,G32267,G32268,G32269,G32270,G32271,G32272,G32273,G32274,G32275,G32276,G32277,G32278,G32279,G32280,
       G32281,G32282,G32283,G32284,G32285,G32286,G32287,G32288,G32289,G32290,G32291,G32292,G32293,G32294,G32295,G32296,G32297,G32298,G32299,G32300,
       G32301,G32302,G32303,G32304,G32305,G32306,G32307,G32308,G32309,G32310,G32311,G32312,G32313,G32314,G32315,G32316,G32317,G32318,G32319,G32320,
       G32321,G32322,G32323,G32324,G32325,G32326,G32327,G32328,G32329,G32330,G32331,G32332,G32333,G32334,G32335,G32336,G32337,G32338,G32339,G32340,
       G32341,G32342,G32343,G32344,G32345,G32346,G32347,G32348,G32349,G32350,G32351,G32352,G32353,G32354,G32355,G32356,G32357,G32358,G32359,G32360,
       G32361,G32362,G32363,G32364,G32365,G32366,G32367,G32368,G32369,G32370,G32371,G32372,G32373,G32374,G32375,G32376,G32377,G32378,G32379,G32380,
       G32381,G32382,G32383,G32384,G32385,G32386,G32387,G32388,G32389,G32390,G32391,G32392,G32393,G32394,G32395,G32396,G32397,G32398,G32399,G32400,
       G32401,G32402,G32403,G32404,G32405,G32406,G32407,G32408,G32409,G32410,G32411,G32412,G32413,G32414,G32415,G32416,G32417,G32418,G32419,G32420,
       G32421,G32422,G32423,G32424,G32425,G32426,G32427,G32428,G32429,G32430,G32431,G32432,G32433,G32434,G32435,G32436,G32437,G32438,G32439,G32440,
       G32441,G32442,G32443,G32444,G32445,G32446,G32447,G32448,G32449,G32450,G32451,G32452,G32453,G32454,G32455,G32456,G32457,G32458,G32459,G32460,
       G32461,G32462,G32463,G32464,G32465,G32466,G32467,G32468,G32469,G32470,G32471,G32472,G32473,G32474,G32475,G32476,G32477,G32478,G32479,G32480,
       G32481,G32482,G32483,G32484,G32485,G32486,G32487,G32488,G32489,G32490,G32491,G32492,G32493,G32494,G32495,G32496,G32497,G32498,G32499,G32500,
       G32501,G32502,G32503,G32504,G32505,G32506,G32507,G32508,G32509,G32510,G32511,G32512,G32513,G32514,G32515,G32516,G32517,G32518,G32519,G32520,
       G32521,G32522,G32523,G32524,G32525,G32526,G32527,G32528,G32529,G32530,G32531,G32532,G32533,G32534,G32535,G32536,G32537,G32538,G32539,G32540,
       G32541,G32542,G32543,G32544,G32545,G32546,G32547,G32548,G32549,G32550,G32551,G32552,G32553,G32554,G32555,G32556,G32557,G32558,G32559,G32560,
       G32561,G32562,G32563,G32564,G32565,G32566,G32567,G32568,G32569,G32570,G32571,G32572,G32573,G32574,G32575,G32576,G32577,G32578,G32579,G32580,
       G32581,G32582,G32583,G32584,G32585,G32586,G32587,G32588,G32589,G32590,G32591,G32592,G32593,G32594,G32595,G32596,G32597,G32598,G32599,G32600,
       G32601,G32602,G32603,G32604,G32605,G32606,G32607,G32608,G32609,G32610,G32611,G32612,G32613,G32614,G32615,G32616,G32617,G32618,G32619,G32620,
       G32621,G32622,G32623,G32624,G32625,G32626,G32627,G32628,G32629,G32630,G32631,G32632,G32633,G32634,G32635,G32636,G32637,G32638,G32639,G32640,
       G32641,G32642,G32643,G32644,G32645,G32646,G32647,G32648,G32649,G32650,G32651,G32652,G32653,G32654,G32655,G32656,G32657,G32658,G32659,G32660,
       G32661,G32662,G32663,G32664,G32665,G32666,G32667,G32668,G32669,G32670,G32671,G32672,G32673,G32674,G32675,G32676,G32677,G32678,G32679,G32680,
       G32681,G32682,G32683,G32684,G32685,G32686,G32687,G32688,G32689,G32690,G32691,G32692,G32693,G32694,G32695,G32696,G32697,G32698,G32699,G32700,
       G32701,G32702,G32703,G32704,G32705,G32706,G32707,G32708,G32709,G32710,G32711,G32712,G32713,G32714,G32715,G32716,G32717,G32718,G32719,G32720,
       G32721,G32722,G32723,G32724,G32725,G32726,G32727,G32728,G32729,G32730,G32731,G32732,G32733,G32734,G32735,G32736,G32737,G32738,G32739,G32740,
       G32741,G32742,G32743,G32744,G32745,G32746,G32747,G32748,G32749,G32750,G32751,G32752,G32753,G32754,G32755,G32756,G32757,G32758,G32759,G32760,
       G32761,G32762,G32763,G32764,G32765,G32766,G32767,G32768,G32769,G32770,G32771,G32772,G32773,G32774,G32775,G32776,G32777,G32778,G32779,G32780,
       G32781,G32782,G32783,G32784,G32785,G32786,G32787,G32788,G32789,G32790,G32791,G32792,G32793,G32794,G32795,G32796,G32797,G32798,G32799,G32800,
       G32801,G32802,G32803,G32804,G32805,G32806,G32807,G32808,G32809,G32810,G32811,G32812,G32813,G32814,G32815,G32816,G32817,G32818,G32819,G32820,
       G32821,G32822,G32823,G32824,G32825,G32826,G32827,G32828,G32829,G32830,G32831,G32832,G32833,G32834,G32835,G32836,G32837,G32838,G32839,G32840,
       G32841,G32842,G32843,G32844,G32845,G32846,G32847,G32848,G32849,G32850,G32851,G32852,G32853,G32854,G32855,G32856,G32857,G32858,G32859,G32860,
       G32861,G32862,G32863,G32864,G32865,G32866,G32867,G32868,G32869,G32870,G32871,G32872,G32873,G32874,G32875,G32876,G32877,G32878,G32879,G32880,
       G32881,G32882,G32883,G32884,G32885,G32886,G32887,G32888,G32889,G32890,G32891,G32892,G32893,G32894,G32895,G32896,G32897,G32898,G32899,G32900,
       G32901,G32902,G32903,G32904,G32905,G32906,G32907,G32908,G32909,G32910,G32911,G32912,G32913,G32914,G32915,G32916,G32917,G32918,G32919,G32920,
       G32921,G32922,G32923,G32924,G32925,G32926,G32927,G32928,G32929,G32930,G32931,G32932,G32933,G32934,G32935,G32936,G32937,G32938,G32939,G32940,
       G32941,G32942,G32943,G32944,G32945,G32946,G32947,G32948,G32949,G32950,G32951,G32952,G32953,G32954,G32955,G32956,G32957,G32958,G32959,G32960,
       G32961,G32962,G32963,G32964,G32965,G32966,G32967,G32968,G32969,G32970,G32971,G32972,G32973,G32974,G32975,G32976,G32977,G32978,G32979,G32980,
       G32981,G32982,G32983,G32984,G32985,G32986,G32987,G32988,G32989,G32990,G32991,G32992,G32993,G32994,G32995,G32996,G32997,G32998,G32999,G33000,
       G33001,G33002,G33003,G33004,G33005,G33006,G33007,G33008,G33009,G33010,G33011,G33012,G33013,G33014,G33015,G33016,G33017,G33018,G33019,G33020,
       G33021,G33022,G33023,G33024,G33025,G33026,G33027,G33028,G33029,G33030,G33031,G33032,G33033,G33034,G33035,G33036,G33037,G33038,G33039,G33040,
       G33041,G33042,G33043,G33044,G33045,G33046,G33047,G33048,G33049,G33050,G33051,G33052,G33053,G33054,G33055,G33056,G33057,G33058,G33059,G33060,
       G33061,G33062,G33063,G33064,G33065,G33066,G33067,G33068,G33069,G33070,G33071,G33072,G33073,G33074,G33075,G33076,G33077,G33078,G33079,G33080,
       G33081,G33082,G33083,G33084,G33085,G33086,G33087,G33088,G33089,G33090,G33091,G33092,G33093,G33094,G33095,G33096,G33097,G33098,G33099,G33100,
       G33101,G33102,G33103,G33104,G33105,G33106,G33107,G33108,G33109,G33110,G33111,G33112,G33113,G33114,G33115,G33116,G33117,G33118,G33119,G33120,
       G33121,G33122,G33123,G33124,G33125,G33126,G33127,G33128,G33129,G33130,G33131,G33132,G33133,G33134,G33135,G33136,G33137,G33138,G33139,G33140,
       G33141,G33142,G33143,G33144,G33145,G33146,G33147,G33148,G33149,G33150,G33151,G33152,G33153,G33154,G33155,G33156,G33157,G33158,G33159,G33160,
       G33161,G33162,G33163,G33164,G33165,G33166,G33167,G33168,G33169,G33170,G33171,G33172,G33173,G33174,G33175,G33176,G33177,G33178,G33179,G33180,
       G33181,G33182,G33183,G33184,G33185,G33186,G33187,G33188,G33189,G33190,G33191,G33192,G33193,G33194,G33195,G33196,G33197,G33198,G33199,G33200,
       G33201,G33202,G33203,G33204,G33205,G33206,G33207,G33208,G33209,G33210,G33211,G33212,G33213,G33214,G33215,G33216,G33217,G33218,G33219,G33220,
       G33221,G33222,G33223,G33224,G33225,G33226,G33227,G33228,G33229,G33230,G33231,G33232,G33233,G33234,G33235,G33236,G33237,G33238,G33239,G33240,
       G33241,G33242,G33243,G33244,G33245,G33246,G33247,G33248,G33249,G33250,G33251,G33252,G33253,G33254,G33255,G33256,G33257,G33258,G33259,G33260,
       G33261,G33262,G33263,G33264,G33265,G33266,G33267,G33268,G33269,G33270,G33271,G33272,G33273,G33274,G33275,G33276,G33277,G33278,G33279,G33280,
       G33281,G33282,G33283,G33284,G33285,G33286,G33287,G33288,G33289,G33290,G33291,G33292,G33293,G33294,G33295,G33296,G33297,G33298,G33299,G33300,
       G33301,G33302,G33303,G33304,G33305,G33306,G33307,G33308,G33309,G33310,G33311,G33312,G33313,G33314,G33315,G33316,G33317,G33318,G33319,G33320,
       G33321,G33322,G33323,G33324,G33325,G33326,G33327,G33328,G33329,G33330,G33331,G33332,G33333,G33334,G33335,G33336,G33337,G33338,G33339,G33340,
       G33341,G33342,G33343,G33344,G33345,G33346,G33347,G33348,G33349,G33350,G33351,G33352,G33353,G33354,G33355,G33356,G33357,G33358,G33359,G33360,
       G33361,G33362,G33363,G33364,G33365,G33366,G33367,G33368,G33369,G33370,G33371,G33372,G33373,G33374,G33375,G33376,G33377,G33378,G33379,G33380,
       G33381,G33382,G33383,G33384,G33385,G33386,G33387,G33388,G33389,G33390,G33391,G33392,G33393,G33394,G33395,G33396,G33397,G33398,G33399,G33400,
       G33401,G33402,G33403,G33404,G33405,G33406,G33407,G33408,G33409,G33410,G33411,G33412,G33413,G33414,G33415,G33416,G33417,G33418,G33419,G33420,
       G33421,G33422,G33423,G33424,G33425,G33426,G33427,G33428,G33429,G33430,G33431,G33432,G33433,G33434,G33435,G33436,G33437,G33438,G33439,G33440,
       G33441,G33442,G33443,G33444,G33445,G33446,G33447,G33448,G33449,G33450,G33451,G33452,G33453,G33454,G33455,G33456,G33457,G33458,G33459,G33460,
       G33461,G33462,G33463,G33464,G33465,G33466,G33467,G33468,G33469,G33470,G33471,G33472,G33473,G33474,G33475,G33476,G33477,G33478,G33479,G33480,
       G33481,G33482,G33483,G33484,G33485,G33486,G33487,G33488,G33489,G33490,G33491,G33492,G33493,G33494,G33495,G33496,G33497,G33498,G33499,G33500,
       G33501,G33502,G33503,G33504,G33505,G33506,G33507,G33508,G33509,G33510,G33511,G33512,G33513,G33514,G33515,G33516,G33517,G33518,G33519,G33520,
       G33521,G33522,G33523,G33524,G33525,G33526,G33527,G33528,G33529,G33530,G33531,G33532,G33533,G33534,G33535,G33536,G33537,G33538,G33539,G33540,
       G33541,G33542,G33543,G33544,G33545,G33546,G33547,G33548,G33549,G33550,G33551,G33552,G33553,G33554,G33555,G33556,G33557,G33558,G33559,G33560,
       G33561,G33562,G33563,G33564,G33565,G33566,G33567,G33568,G33569,G33570,G33571,G33572,G33573,G33574,G33575,G33576,G33577,G33578,G33579,G33580,
       G33581,G33582,G33583,G33584,G33585,G33586,G33587,G33588,G33589,G33590,G33591,G33592,G33593,G33594,G33595,G33596,G33597,G33598,G33599,G33600,
       G33601,G33602,G33603,G33604,G33605,G33606,G33607,G33608,G33609,G33610,G33611,G33612,G33613,G33614,G33615,G33616,G33617,G33618,G33619,G33620,
       G33621,G33622,G33623,G33624,G33625,G33626,G33627,G33628,G33629,G33630,G33631,G33632,G33633,G33634,G33635,G33636,G33637,G33638,G33639,G33640,
       G33641,G33642,G33643,G33644,G33645,G33646,G33647,G33648,G33649,G33650,G33651,G33652,G33653,G33654,G33655,G33656,G33657,G33658,G33659,G33660,
       G33661,G33662,G33663,G33664,G33665,G33666,G33667,G33668,G33669,G33670,G33671,G33672,G33673,G33674,G33675,G33676,G33677,G33678,G33679,G33680,
       G33681,G33682,G33683,G33684,G33685,G33686,G33687,G33688,G33689,G33690,G33691,G33692,G33693,G33694,G33695,G33696,G33697,G33698,G33699,G33700,
       G33701,G33702,G33703,G33704,G33705,G33706,G33707,G33708,G33709,G33710,G33711,G33712,G33713,G33714,G33715,G33716,G33717,G33718,G33719,G33720,
       G33721,G33722,G33723,G33724,G33725,G33726,G33727,G33728,G33729,G33730,G33731,G33732,G33733,G33734,G33735,G33736,G33737,G33738,G33739,G33740,
       G33741,G33742,G33743,G33744,G33745,G33746,G33747,G33748,G33749,G33750,G33751,G33752,G33753,G33754,G33755,G33756,G33757,G33758,G33759,G33760,
       G33761,G33762,G33763,G33764,G33765,G33766,G33767,G33768,G33769,G33770,G33771,G33772,G33773,G33774,G33775,G33776,G33777,G33778,G33779,G33780,
       G33781,G33782,G33783,G33784,G33785,G33786,G33787,G33788,G33789,G33790,G33791,G33792,G33793,G33794,G33795,G33796,G33797,G33798,G33799,G33800,
       G33801,G33802,G33803,G33804,G33805,G33806,G33807,G33808,G33809,G33810,G33811,G33812,G33813,G33814,G33815,G33816,G33817,G33818,G33819,G33820,
       G33821,G33822,G33823,G33824,G33825,G33826,G33827,G33828,G33829,G33830,G33831,G33832,G33833,G33834,G33835,G33836,G33837,G33838,G33839,G33840,
       G33841,G33842,G33843,G33844,G33845,G33846,G33847,G33848,G33849,G33850,G33851,G33852,G33853,G33854,G33855,G33856,G33857,G33858,G33859,G33860,
       G33861,G33862,G33863,G33864,G33865,G33866,G33867,G33868,G33869,G33870,G33871,G33872,G33873,G33874,G33875,G33876,G33877,G33878,G33879,G33880,
       G33881,G33882,G33883,G33884,G33885,G33886,G33887,G33888,G33889,G33890,G33891,G33892,G33893,G33894,G33895,G33896,G33897,G33898,G33899,G33900,
       G33901,G33902,G33903,G33904,G33905,G33906,G33907,G33908,G33909,G33910,G33911,G33912,G33913,G33914,G33915,G33916,G33917,G33918,G33919,G33920,
       G33921,G33922,G33923,G33924,G33925,G33926,G33927,G33928,G33929,G33930,G33931,G33932,G33933,G33934,G33935,G33936,G33937,G33938,G33939,G33940,
       G33941,G33942,G33943,G33944,G33945,G33946,G33947,G33948,G33949,G33950,G33951,G33952,G33953,G33954,G33955,G33956,G33957,G33958,G33959,G33960,
       G33961,G33962,G33963,G33964,G33965,G33966,G33967,G33968,G33969,G33970,G33971,G33972,G33973,G33974,G33975,G33976,G33977,G33978,G33979,G33980,
       G33981,G33982,G33983,G33984,G33985,G33986,G33987,G33988,G33989,G33990,G33991,G33992,G33993,G33994,G33995,G33996,G33997,G33998,G33999,G34000,
       G34001,G34002,G34003,G34004,G34005,G34006,G34007,G34008,G34009,G34010,G34011,G34012,G34013,G34014,G34015,G34016,G34017,G34018,G34019,G34020,
       G34021,G34022,G34023,G34024,G34025,G34026,G34027,G34028,G34029,G34030,G34031,G34032,G34033,G34034,G34035,G34036,G34037,G34038,G34039,G34040,
       G34041,G34042,G34043,G34044,G34045,G34046,G34047,G34048,G34049,G34050,G34051,G34052,G34053,G34054,G34055,G34056,G34057,G34058,G34059,G34060,
       G34061,G34062,G34063,G34064,G34065,G34066,G34067,G34068,G34069,G34070,G34071,G34072,G34073,G34074,G34075,G34076,G34077,G34078,G34079,G34080,
       G34081,G34082,G34083,G34084,G34085,G34086,G34087,G34088,G34089,G34090,G34091,G34092,G34093,G34094,G34095,G34096,G34097,G34098,G34099,G34100,
       G34101,G34102,G34103,G34104,G34105,G34106,G34107,G34108,G34109,G34110,G34111,G34112,G34113,G34114,G34115,G34116,G34117,G34118,G34119,G34120,
       G34121,G34122,G34123,G34124,G34125,G34126,G34127,G34128,G34129,G34130,G34131,G34132,G34133,G34134,G34135,G34136,G34137,G34138,G34139,G34140,
       G34141,G34142,G34143,G34144,G34145,G34146,G34147,G34148,G34149,G34150,G34151,G34152,G34153,G34154,G34155,G34156,G34157,G34158,G34159,G34160,
       G34161,G34162,G34163,G34164,G34165,G34166,G34167,G34168,G34169,G34170,G34171,G34172,G34173,G34174,G34175,G34176,G34177,G34178,G34179,G34180,
       G34181,G34182,G34183,G34184,G34185,G34186,G34187,G34188,G34189,G34190,G34191,G34192,G34193,G34194,G34195,G34196,G34197,G34198,G34199,G34200,
       G34201,G34202,G34203,G34204,G34205,G34206,G34207,G34208,G34209,G34210,G34211,G34212,G34213,G34214,G34215,G34216,G34217,G34218,G34219,G34220,
       G34221,G34222,G34223,G34224,G34225,G34226,G34227,G34228,G34229,G34230,G34231,G34232,G34233,G34234,G34235,G34236,G34237,G34238,G34239,G34240,
       G34241,G34242,G34243,G34244,G34245,G34246,G34247,G34248,G34249,G34250,G34251,G34252,G34253,G34254,G34255,G34256,G34257,G34258,G34259,G34260,
       G34261,G34262,G34263,G34264,G34265,G34266,G34267,G34268,G34269,G34270,G34271,G34272,G34273,G34274,G34275,G34276,G34277,G34278,G34279,G34280,
       G34281,G34282,G34283,G34284,G34285,G34286,G34287,G34288,G34289,G34290,G34291,G34292,G34293,G34294,G34295,G34296,G34297,G34298,G34299,G34300,
       G34301,G34302,G34303,G34304,G34305,G34306,G34307,G34308,G34309,G34310,G34311,G34312,G34313,G34314,G34315,G34316,G34317,G34318,G34319,G34320,
       G34321,G34322,G34323,G34324,G34325,G34326,G34327,G34328,G34329,G34330,G34331,G34332,G34333,G34334,G34335,G34336,G34337,G34338,G34339,G34340,
       G34341,G34342,G34343,G34344,G34345,G34346,G34347,G34348,G34349,G34350,G34351,G34352,G34353,G34354,G34355,G34356,G34357,G34358,G34359,G34360,
       G34361,G34362,G34363,G34364,G34365,G34366,G34367,G34368,G34369,G34370,G34371,G34372,G34373,G34374,G34375,G34376,G34377,G34378,G34379,G34380,
       G34381,G34382,G34383,G34384,G34385,G34386,G34387,G34388,G34389,G34390,G34391,G34392,G34393,G34394,G34395,G34396,G34397,G34398,G34399,G34400,
       G34401,G34402,G34403,G34404,G34405,G34406,G34407,G34408,G34409,G34410,G34411,G34412,G34413,G34414,G34415,G34416,G34417,G34418,G34419,G34420,
       G34421,G34422,G34423,G34424,G34425,G34426,G34427,G34428,G34429,G34430,G34431,G34432,G34433,G34434,G34435,G34436,G34437,G34438,G34439,G34440,
       G34441,G34442,G34443,G34444,G34445,G34446,G34447,G34448,G34449,G34450,G34451,G34452,G34453,G34454,G34455,G34456,G34457,G34458,G34459,G34460,
       G34461,G34462,G34463,G34464,G34465,G34466,G34467,G34468,G34469,G34470,G34471,G34472,G34473,G34474,G34475,G34476,G34477,G34478,G34479,G34480,
       G34481,G34482,G34483,G34484,G34485,G34486,G34487,G34488,G34489,G34490,G34491,G34492,G34493,G34494,G34495,G34496,G34497,G34498,G34499,G34500,
       G34501,G34502,G34503,G34504,G34505,G34506,G34507,G34508,G34509,G34510,G34511,G34512,G34513,G34514,G34515,G34516,G34517,G34518,G34519,G34520,
       G34521,G34522,G34523,G34524,G34525,G34526,G34527,G34528,G34529,G34530,G34531,G34532,G34533,G34534,G34535,G34536,G34537,G34538,G34539,G34540,
       G34541,G34542,G34543,G34544,G34545,G34546,G34547,G34548,G34549,G34550,G34551,G34552,G34553,G34554,G34555,G34556,G34557,G34558,G34559,G34560,
       G34561,G34562,G34563,G34564,G34565,G34566,G34567,G34568,G34569,G34570,G34571,G34572,G34573,G34574,G34575,G34576,G34577,G34578,G34579,G34580,
       G34581,G34582,G34583,G34584,G34585,G34586,G34587,G34588,G34589,G34590,G34591,G34592,G34593,G34594,G34595,G34596,G34597,G34598,G34599,G34600,
       G34601,G34602,G34603,G34604,G34605,G34606,G34607,G34608,G34609,G34610,G34611,G34612,G34613,G34614,G34615,G34616,G34617,G34618,G34619,G34620,
       G34621,G34622,G34623,G34624,G34625,G34626,G34627,G34628,G34629,G34630,G34631,G34632,G34633,G34634,G34635,G34636,G34637,G34638,G34639,G34640,
       G34641,G34642,G34643,G34644,G34645,G34646,G34647,G34648,G34649,G34650,G34651,G34652,G34653,G34654,G34655,G34656,G34657,G34658,G34659,G34660,
       G34661,G34662,G34663,G34664,G34665,G34666,G34667,G34668,G34669,G34670,G34671,G34672,G34673,G34674,G34675,G34676,G34677,G34678,G34679,G34680,
       G34681,G34682,G34683,G34684,G34685,G34686,G34687,G34688,G34689,G34690,G34691,G34692,G34693,G34694,G34695,G34696,G34697,G34698,G34699,G34700,
       G34701,G34702,G34703,G34704,G34705,G34706,G34707,G34708,G34709,G34710,G34711,G34712,G34713,G34714,G34715,G34716,G34717,G34718,G34719,G34720,
       G34721,G34722,G34723,G34724,G34725,G34726,G34727,G34728,G34729,G34730,G34731,G34732,G34733,G34734,G34735,G34736,G34737,G34738,G34739,G34740,
       G34741,G34742,G34743,G34744,G34745,G34746,G34747,G34748,G34749,G34750,G34751,G34752,G34753,G34754,G34755,G34756,G34757,G34758,G34759,G34760,
       G34761,G34762,G34763,G34764,G34765,G34766,G34767,G34768,G34769,G34770,G34771,G34772,G34773,G34774,G34775,G34776,G34777,G34778,G34779,G34780,
       G34781,G34782,G34783,G34784,G34785,G34786,G34787,G34788,G34789,G34790,G34791,G34792,G34793,G34794,G34795,G34796,G34797,G34798,G34799,G34800,
       G34801,G34802,G34803,G34804,G34805,G34806,G34807,G34808,G34809,G34810,G34811,G34812,G34813,G34814,G34815,G34816,G34817,G34818,G34819,G34820,
       G34821,G34822,G34823,G34824,G34825,G34826,G34827,G34828,G34829,G34830,G34831,G34832,G34833,G34834,G34835,G34836,G34837,G34838,G34839,G34840,
       G34841,G34842,G34843,G34844,G34845,G34846,G34847,G34848,G34849,G34850,G34851,G34852,G34853,G34854,G34855,G34856,G34857,G34858,G34859,G34860,
       G34861,G34862,G34863,G34864,G34865,G34866,G34867,G34868,G34869,G34870,G34871,G34872,G34873,G34874,G34875,G34876,G34877,G34878,G34879,G34880,
       G34881,G34882,G34883,G34884,G34885,G34886,G34887,G34888,G34889,G34890,G34891,G34892,G34893,G34894,G34895,G34896,G34897,G34898,G34899,G34900,
       G34901,G34902,G34903,G34904,G34905,G34906,G34907,G34908,G34909,G34910,G34911,G34912,G34913,G34914,G34915,G34916,G34917,G34918,G34919,G34920,
       G34921,G34922,G34923,G34924,G34925,G34926,G34927,G34928,G34929,G34930,G34931,G34932,G34933,G34934,G34935,G34936,G34937,G34938,G34939,G34940,
       G34941,G34942,G34943,G34944,G34945,G34946,G34947,G34948,G34949,G34950,G34951,G34952,G34953,G34954,G34955,G34956,G34957,G34958,G34959,G34960,
       G34961,G34962,G34963,G34964,G34965,G34966,G34967,G34968,G34969,G34970,G34971,G34972,G34973,G34974,G34975,G34976,G34977,G34978,G34979,G34980,
       G34981,G34982,G34983,G34984,G34985,G34986,G34987,G34988,G34989,G34990,G34991,G34992,G34993,G34994,G34995,G34996,G34997,G34998,G34999,G35000,
       G35001,G35002,G35003,G35004,G35005,G35006,G35007,G35008,G35009,G35010,G35011,G35012,G35013,G35014,G35015,G35016,G35017,G35018,G35019,G35020,
       G35021,G35022,G35023,G35024,G35025,G35026,G35027,G35028,G35029,G35030,G35031,G35032,G35033,G35034,G35035,G35036,G35037,G35038,G35039,G35040,
       G35041,G35042,G35043,G35044,G35045,G35046,G35047,G35048,G35049,G35050,G35051,G35052,G35053,G35054,G35055,G35056,G35057,G35058,G35059,G35060,
       G35061,G35062,G35063,G35064,G35065,G35066,G35067,G35068,G35069,G35070,G35071,G35072,G35073,G35074,G35075,G35076,G35077,G35078,G35079,G35080,
       G35081,G35082,G35083,G35084,G35085,G35086,G35087,G35088,G35089,G35090,G35091,G35092,G35093,G35094,G35095,G35096,G35097,G35098,G35099,G35100,
       G35101,G35102,G35103,G35104,G35105,G35106,G35107,G35108,G35109,G35110,G35111,G35112,G35113,G35114,G35115,G35116,G35117,G35118,G35119,G35120,
       G35121,G35122,G35123,G35124,G35125,G35126,G35127,G35128,G35129,G35130,G35131,G35132,G35133,G35134,G35135,G35136,G35137,G35138,G35139,G35140,
       G35141,G35142,G35143,G35144,G35145,G35146,G35147,G35148,G35149,G35150,G35151,G35152,G35153,G35154,G35155,G35156,G35157,G35158,G35159,G35160,
       G35161,G35162,G35163,G35164,G35165,G35166,G35167,G35168,G35169,G35170,G35171,G35172,G35173,G35174,G35175,G35176,G35177,G35178,G35179,G35180,
       G35181,G35182,G35183,G35184,G35185,G35186,G35187,G35188,G35189,G35190,G35191,G35192,G35193,G35194,G35195,G35196,G35197,G35198,G35199,G35200,
       G35201,G35202,G35203,G35204,G35205,G35206,G35207,G35208,G35209,G35210,G35211,G35212,G35213,G35214,G35215,G35216,G35217,G35218,G35219,G35220,
       G35221,G35222,G35223,G35224,G35225,G35226,G35227,G35228,G35229,G35230,G35231,G35232,G35233,G35234,G35235,G35236,G35237,G35238,G35239,G35240,
       G35241,G35242,G35243,G35244,G35245,G35246,G35247,G35248,G35249,G35250,G35251,G35252,G35253,G35254,G35255,G35256,G35257,G35258,G35259,G35260,
       G35261,G35262,G35263,G35264,G35265,G35266,G35267,G35268,G35269,G35270,G35271,G35272,G35273,G35274,G35275,G35276,G35277,G35278,G35279,G35280,
       G35281,G35282,G35283,G35284,G35285,G35286,G35287,G35288,G35289,G35290,G35291,G35292,G35293,G35294,G35295,G35296,G35297,G35298,G35299,G35300,
       G35301,G35302,G35303,G35304,G35305,G35306,G35307,G35308,G35309,G35310,G35311,G35312,G35313,G35314,G35315,G35316,G35317,G35318,G35319,G35320,
       G35321,G35322,G35323,G35324,G35325,G35326,G35327,G35328,G35329,G35330,G35331,G35332,G35333,G35334,G35335,G35336,G35337,G35338,G35339,G35340,
       G35341,G35342,G35343,G35344,G35345,G35346,G35347,G35348,G35349,G35350,G35351,G35352,G35353,G35354,G35355,G35356,G35357,G35358,G35359,G35360,
       G35361,G35362,G35363,G35364,G35365,G35366,G35367,G35368,G35369,G35370,G35371,G35372,G35373,G35374,G35375,G35376,G35377,G35378,G35379,G35380,
       G35381,G35382,G35383,G35384,G35385,G35386,G35387,G35388,G35389,G35390,G35391,G35392,G35393,G35394,G35395,G35396,G35397,G35398,G35399,G35400,
       G35401,G35402,G35403,G35404,G35405,G35406,G35407,G35408,G35409,G35410,G35411,G35412,G35413,G35414,G35415,G35416,G35417,G35418,G35419,G35420,
       G35421,G35422,G35423,G35424,G35425,G35426,G35427,G35428,G35429,G35430,G35431,G35432,G35433,G35434,G35435,G35436,G35437,G35438,G35439,G35440,
       G35441,G35442,G35443,G35444,G35445,G35446,G35447,G35448,G35449,G35450,G35451,G35452,G35453,G35454,G35455,G35456,G35457,G35458,G35459,G35460,
       G35461,G35462,G35463,G35464,G35465,G35466,G35467,G35468,G35469,G35470,G35471,G35472,G35473,G35474,G35475,G35476,G35477,G35478,G35479,G35480,
       G35481,G35482,G35483,G35484,G35485,G35486,G35487,G35488,G35489,G35490,G35491,G35492,G35493,G35494,G35495,G35496,G35497,G35498,G35499,G35500,
       G35501,G35502,G35503,G35504,G35505,G35506,G35507,G35508,G35509,G35510,G35511,G35512,G35513,G35514,G35515,G35516,G35517,G35518,G35519,G35520,
       G35521,G35522,G35523,G35524,G35525,G35526,G35527,G35528,G35529,G35530,G35531,G35532,G35533,G35534,G35535,G35536,G35537,G35538,G35539,G35540,
       G35541,G35542,G35543,G35544,G35545,G35546,G35547,G35548,G35549,G35550,G35551,G35552,G35553,G35554,G35555,G35556,G35557,G35558,G35559,G35560,
       G35561,G35562,G35563,G35564,G35565,G35566,G35567,G35568,G35569,G35570,G35571,G35572,G35573,G35574,G35575,G35576,G35577,G35578,G35579,G35580,
       G35581,G35582,G35583,G35584,G35585,G35586,G35587,G35588,G35589,G35590,G35591,G35592,G35593,G35594,G35595,G35596,G35597,G35598,G35599,G35600,
       G35601,G35602,G35603,G35604,G35605,G35606,G35607,G35608,G35609,G35610,G35611,G35612,G35613,G35614,G35615,G35616,G35617,G35618,G35619,G35620,
       G35621,G35622,G35623,G35624,G35625,G35626,G35627,G35628,G35629,G35630,G35631,G35632,G35633,G35634,G35635,G35636,G35637,G35638,G35639,G35640,
       G35641,G35642,G35643,G35644,G35645,G35646,G35647,G35648,G35649,G35650,G35651,G35652,G35653,G35654,G35655,G35656,G35657,G35658,G35659,G35660,
       G35661,G35662,G35663,G35664,G35665,G35666,G35667,G35668,G35669,G35670,G35671,G35672,G35673,G35674,G35675,G35676,G35677,G35678,G35679,G35680,
       G35681,G35682,G35683,G35684,G35685,G35686,G35687,G35688,G35689,G35690,G35691,G35692,G35693,G35694,G35695,G35696,G35697,G35698,G35699,G35700,
       G35701,G35702,G35703,G35704,G35705,G35706,G35707,G35708,G35709,G35710,G35711,G35712,G35713,G35714,G35715,G35716,G35717,G35718,G35719,G35720,
       G35721,G35722,G35723,G35724,G35725,G35726,G35727,G35728,G35729,G35730,G35731,G35732,G35733,G35734,G35735,G35736,G35737,G35738,G35739,G35740,
       G35741,G35742,G35743,G35744,G35745,G35746,G35747,G35748,G35749,G35750,G35751,G35752,G35753,G35754,G35755,G35756,G35757,G35758,G35759,G35760,
       G35761,G35762,G35763,G35764,G35765,G35766,G35767,G35768,G35769,G35770,G35771,G35772,G35773,G35774,G35775,G35776,G35777,G35778,G35779,G35780,
       G35781,G35782,G35783,G35784,G35785,G35786,G35787,G35788,G35789,G35790,G35791,G35792,G35793,G35794,G35795,G35796,G35797,G35798,G35799,G35800,
       G35801,G35802,G35803,G35804,G35805,G35806,G35807,G35808,G35809,G35810,G35811,G35812,G35813,G35814,G35815,G35816,G35817,G35818,G35819,G35820,
       G35821,G35822,G35823,G35824,G35825,G35826,G35827,G35828,G35829,G35830,G35831,G35832,G35833,G35834,G35835,G35836,G35837,G35838,G35839,G35840,
       G35841,G35842,G35843,G35844,G35845,G35846,G35847,G35848,G35849,G35850,G35851,G35852,G35853,G35854,G35855,G35856,G35857,G35858,G35859,G35860,
       G35861,G35862,G35863,G35864,G35865,G35866,G35867,G35868,G35869,G35870,G35871,G35872,G35873,G35874,G35875,G35876,G35877,G35878,G35879,G35880,
       G35881,G35882,G35883,G35884,G35885,G35886,G35887,G35888,G35889,G35890,G35891,G35892,G35893,G35894,G35895,G35896,G35897,G35898,G35899,G35900,
       G35901,G35902,G35903,G35904,G35905,G35906,G35907,G35908,G35909,G35910,G35911,G35912,G35913,G35914,G35915,G35916,G35917,G35918,G35919,G35920,
       G35921,G35922,G35923,G35924,G35925,G35926,G35927,G35928,G35929,G35930,G35931,G35932,G35933,G35934,G35935,G35936,G35937,G35938,G35939,G35940,
       G35941,G35942,G35943,G35944,G35945,G35946,G35947,G35948,G35949,G35950,G35951,G35952,G35953,G35954,G35955,G35956,G35957,G35958,G35959,G35960,
       G35961,G35962,G35963,G35964,G35965,G35966,G35967,G35968,G35969,G35970,G35971,G35972,G35973,G35974,G35975,G35976,G35977,G35978,G35979,G35980,
       G35981,G35982,G35983,G35984,G35985,G35986,G35987,G35988,G35989,G35990,G35991,G35992,G35993,G35994,G35995,G35996,G35997,G35998,G35999,G36000,
       G36001,G36002,G36003,G36004,G36005,G36006,G36007,G36008,G36009,G36010,G36011,G36012,G36013,G36014,G36015,G36016,G36017,G36018,G36019,G36020,
       G36021,G36022,G36023,G36024,G36025,G36026,G36027,G36028,G36029,G36030,G36031,G36032,G36033,G36034,G36035,G36036,G36037,G36038,G36039,G36040,
       G36041,G36042,G36043,G36044,G36045,G36046,G36047,G36048,G36049,G36050,G36051,G36052,G36053,G36054,G36055,G36056,G36057,G36058,G36059,G36060,
       G36061,G36062,G36063,G36064,G36065,G36066,G36067,G36068,G36069,G36070,G36071,G36072,G36073,G36074,G36075,G36076,G36077,G36078,G36079,G36080,
       G36081,G36082,G36083,G36084,G36085,G36086,G36087,G36088,G36089,G36090,G36091,G36092,G36093,G36094,G36095,G36096,G36097,G36098,G36099,G36100,
       G36101,G36102,G36103,G36104,G36105,G36106,G36107,G36108,G36109,G36110,G36111,G36112,G36113,G36114,G36115,G36116,G36117,G36118,G36119,G36120,
       G36121,G36122,G36123,G36124,G36125,G36126,G36127,G36128,G36129,G36130,G36131,G36132,G36133,G36134,G36135,G36136,G36137,G36138,G36139,G36140,
       G36141,G36142,G36143,G36144,G36145,G36146,G36147,G36148,G36149,G36150,G36151,G36152,G36153,G36154,G36155,G36156,G36157,G36158,G36159,G36160,
       G36161,G36162,G36163,G36164,G36165,G36166,G36167,G36168,G36169,G36170,G36171,G36172,G36173,G36174,G36175,G36176,G36177,G36178,G36179,G36180,
       G36181,G36182,G36183,G36184,G36185,G36186,G36187,G36188,G36189,G36190,G36191,G36192,G36193,G36194,G36195,G36196,G36197,G36198,G36199,G36200,
       G36201,G36202,G36203,G36204,G36205,G36206,G36207,G36208,G36209,G36210,G36211,G36212,G36213,G36214,G36215,G36216,G36217,G36218,G36219,G36220,
       G36221,G36222,G36223,G36224,G36225,G36226,G36227,G36228,G36229,G36230,G36231,G36232,G36233,G36234,G36235,G36236,G36237,G36238,G36239,G36240,
       G36241,G36242,G36243,G36244,G36245,G36246,G36247,G36248,G36249,G36250,G36251,G36252,G36253,G36254,G36255,G36256,G36257,G36258,G36259,G36260,
       G36261,G36262,G36263,G36264,G36265,G36266,G36267,G36268,G36269,G36270,G36271,G36272,G36273,G36274,G36275,G36276,G36277,G36278,G36279,G36280,
       G36281,G36282,G36283,G36284,G36285,G36286,G36287,G36288,G36289,G36290,G36291,G36292,G36293,G36294,G36295,G36296,G36297,G36298,G36299,G36300,
       G36301,G36302,G36303,G36304,G36305,G36306,G36307,G36308,G36309,G36310,G36311,G36312,G36313,G36314,G36315,G36316,G36317,G36318,G36319,G36320,
       G36321,G36322,G36323,G36324,G36325,G36326,G36327,G36328,G36329,G36330,G36331,G36332,G36333,G36334,G36335,G36336,G36337,G36338,G36339,G36340,
       G36341,G36342,G36343,G36344,G36345,G36346,G36347,G36348,G36349,G36350,G36351,G36352,G36353,G36354,G36355,G36356,G36357,G36358,G36359,G36360,
       G36361,G36362,G36363,G36364,G36365,G36366,G36367,G36368,G36369,G36370,G36371,G36372,G36373,G36374,G36375,G36376,G36377,G36378,G36379,G36380,
       G36381,G36382,G36383,G36384,G36385,G36386,G36387,G36388,G36389,G36390,G36391,G36392,G36393,G36394,G36395,G36396,G36397,G36398,G36399,G36400,
       G36401,G36402,G36403,G36404,G36405,G36406,G36407,G36408,G36409,G36410,G36411,G36412,G36413,G36414,G36415,G36416,G36417,G36418,G36419,G36420,
       G36421,G36422,G36423,G36424,G36425,G36426,G36427,G36428,G36429,G36430,G36431,G36432,G36433,G36434,G36435,G36436,G36437,G36438,G36439,G36440,
       G36441,G36442,G36443,G36444,G36445,G36446,G36447,G36448,G36449,G36450,G36451,G36452,G36453,G36454,G36455,G36456,G36457,G36458,G36459,G36460,
       G36461,G36462,G36463,G36464,G36465,G36466,G36467,G36468,G36469,G36470,G36471,G36472,G36473,G36474,G36475,G36476,G36477,G36478,G36479,G36480,
       G36481,G36482,G36483,G36484,G36485,G36486,G36487,G36488,G36489,G36490,G36491,G36492,G36493,G36494,G36495,G36496,G36497,G36498,G36499,G36500,
       G36501,G36502,G36503,G36504,G36505,G36506,G36507,G36508,G36509,G36510,G36511,G36512,G36513,G36514,G36515,G36516,G36517,G36518,G36519,G36520,
       G36521,G36522,G36523,G36524,G36525,G36526,G36527,G36528,G36529,G36530,G36531,G36532,G36533,G36534,G36535,G36536,G36537,G36538,G36539,G36540,
       G36541,G36542,G36543,G36544,G36545,G36546,G36547,G36548,G36549,G36550,G36551,G36552,G36553,G36554,G36555,G36556,G36557,G36558,G36559,G36560,
       G36561,G36562,G36563,G36564,G36565,G36566,G36567,G36568,G36569,G36570,G36571,G36572,G36573,G36574,G36575,G36576,G36577,G36578,G36579,G36580,
       G36581,G36582,G36583,G36584,G36585,G36586,G36587,G36588,G36589,G36590,G36591,G36592,G36593,G36594,G36595,G36596,G36597,G36598,G36599,G36600,
       G36601,G36602,G36603,G36604,G36605,G36606,G36607,G36608,G36609,G36610,G36611,G36612,G36613,G36614,G36615,G36616,G36617,G36618,G36619,G36620,
       G36621,G36622,G36623,G36624,G36625,G36626,G36627,G36628,G36629,G36630,G36631,G36632,G36633,G36634,G36635,G36636,G36637,G36638,G36639,G36640,
       G36641,G36642,G36643,G36644,G36645,G36646,G36647,G36648,G36649,G36650,G36651,G36652,G36653,G36654,G36655,G36656,G36657,G36658,G36659,G36660,
       G36661,G36662,G36663,G36664,G36665,G36666,G36667,G36668,G36669,G36670,G36671,G36672,G36673,G36674,G36675,G36676,G36677,G36678,G36679,G36680,
       G36681,G36682,G36683,G36684,G36685,G36686,G36687,G36688,G36689,G36690,G36691,G36692,G36693,G36694,G36695,G36696,G36697,G36698,G36699,G36700,
       G36701,G36702,G36703,G36704,G36705,G36706,G36707,G36708,G36709,G36710,G36711,G36712,G36713,G36714,G36715,G36716,G36717,G36718,G36719,G36720,
       G36721,G36722,G36723,G36724,G36725,G36726,G36727,G36728,G36729,G36730,G36731,G36732,G36733,G36734,G36735,G36736,G36737,G36738,G36739,G36740,
       G36741,G36742,G36743,G36744,G36745,G36746,G36747,G36748,G36749,G36750,G36751,G36752,G36753,G36754,G36755,G36756,G36757,G36758,G36759,G36760,
       G36761,G36762,G36763,G36764,G36765,G36766,G36767,G36768,G36769,G36770,G36771,G36772,G36773,G36774,G36775,G36776,G36777,G36778,G36779,G36780,
       G36781,G36782,G36783,G36784,G36785,G36786,G36787,G36788,G36789,G36790,G36791,G36792,G36793,G36794,G36795,G36796,G36797,G36798,G36799,G36800,
       G36801,G36802,G36803,G36804,G36805,G36806,G36807,G36808,G36809,G36810,G36811,G36812,G36813,G36814,G36815,G36816,G36817,G36818,G36819,G36820,
       G36821,G36822,G36823,G36824,G36825,G36826,G36827,G36828,G36829,G36830,G36831,G36832,G36833,G36834,G36835,G36836,G36837,G36838,G36839,G36840,
       G36841,G36842,G36843,G36844,G36845,G36846,G36847,G36848,G36849,G36850,G36851,G36852,G36853,G36854,G36855,G36856,G36857,G36858,G36859,G36860,
       G36861,G36862,G36863,G36864,G36865,G36866,G36867,G36868,G36869,G36870,G36871,G36872,G36873,G36874,G36875,G36876,G36877,G36878,G36879,G36880,
       G36881,G36882,G36883,G36884,G36885,G36886,G36887,G36888,G36889,G36890,G36891,G36892,G36893,G36894,G36895,G36896,G36897,G36898,G36899,G36900,
       G36901,G36902,G36903,G36904,G36905,G36906,G36907,G36908,G36909,G36910,G36911,G36912,G36913,G36914,G36915,G36916,G36917,G36918,G36919,G36920,
       G36921,G36922,G36923,G36924,G36925,G36926,G36927,G36928,G36929,G36930,G36931,G36932,G36933,G36934,G36935,G36936,G36937,G36938,G36939,G36940,
       G36941,G36942,G36943,G36944,G36945,G36946,G36947,G36948,G36949,G36950,G36951,G36952,G36953,G36954,G36955,G36956,G36957,G36958,G36959,G36960,
       G36961,G36962,G36963,G36964,G36965,G36966,G36967,G36968,G36969,G36970,G36971,G36972,G36973,G36974,G36975,G36976,G36977,G36978,G36979,G36980,
       G36981,G36982,G36983,G36984,G36985,G36986,G36987,G36988,G36989,G36990,G36991,G36992,G36993,G36994,G36995,G36996,G36997,G36998,G36999,G37000,
       G37001,G37002,G37003,G37004,G37005,G37006,G37007,G37008,G37009,G37010,G37011,G37012,G37013,G37014,G37015,G37016,G37017,G37018,G37019,G37020,
       G37021,G37022,G37023,G37024,G37025,G37026,G37027,G37028,G37029,G37030,G37031,G37032,G37033,G37034,G37035,G37036,G37037,G37038,G37039,G37040,
       G37041,G37042,G37043,G37044,G37045,G37046,G37047,G37048,G37049,G37050,G37051,G37052,G37053,G37054,G37055,G37056,G37057,G37058,G37059,G37060,
       G37061,G37062,G37063,G37064,G37065,G37066,G37067,G37068,G37069,G37070,G37071,G37072,G37073,G37074,G37075,G37076,G37077,G37078,G37079,G37080,
       G37081,G37082,G37083,G37084,G37085,G37086,G37087,G37088,G37089,G37090,G37091,G37092,G37093,G37094,G37095,G37096,G37097,G37098,G37099,G37100,
       G37101,G37102,G37103,G37104,G37105,G37106,G37107,G37108,G37109,G37110,G37111,G37112,G37113,G37114,G37115,G37116,G37117,G37118,G37119,G37120,
       G37121,G37122,G37123,G37124,G37125,G37126,G37127,G37128,G37129,G37130,G37131,G37132,G37133,G37134,G37135,G37136,G37137,G37138,G37139,G37140,
       G37141,G37142,G37143,G37144,G37145,G37146,G37147,G37148,G37149,G37150,G37151,G37152,G37153,G37154,G37155,G37156,G37157,G37158,G37159,G37160,
       G37161,G37162,G37163,G37164,G37165,G37166,G37167,G37168,G37169,G37170,G37171,G37172,G37173,G37174,G37175,G37176,G37177,G37178,G37179,G37180,
       G37181,G37182,G37183,G37184,G37185,G37186,G37187,G37188,G37189,G37190,G37191,G37192,G37193,G37194,G37195,G37196,G37197,G37198,G37199,G37200,
       G37201,G37202,G37203,G37204,G37205,G37206,G37207,G37208,G37209,G37210,G37211,G37212,G37213,G37214,G37215,G37216,G37217,G37218,G37219,G37220,
       G37221,G37222,G37223,G37224,G37225,G37226,G37227,G37228,G37229,G37230,G37231,G37232,G37233,G37234,G37235,G37236,G37237,G37238,G37239,G37240,
       G37241,G37242,G37243,G37244,G37245,G37246,G37247,G37248,G37249,G37250,G37251,G37252,G37253,G37254,G37255,G37256,G37257,G37258,G37259,G37260,
       G37261,G37262,G37263,G37264,G37265,G37266,G37267,G37268,G37269,G37270,G37271,G37272,G37273,G37274,G37275,G37276,G37277,G37278,G37279,G37280,
       G37281,G37282,G37283,G37284,G37285,G37286,G37287,G37288,G37289,G37290,G37291,G37292,G37293,G37294,G37295,G37296,G37297,G37298,G37299,G37300,
       G37301,G37302,G37303,G37304,G37305,G37306,G37307,G37308,G37309,G37310,G37311,G37312,G37313,G37314,G37315,G37316,G37317,G37318,G37319,G37320,
       G37321,G37322,G37323,G37324,G37325,G37326,G37327,G37328,G37329,G37330,G37331,G37332,G37333,G37334,G37335,G37336,G37337,G37338,G37339,G37340,
       G37341,G37342,G37343,G37344,G37345,G37346,G37347,G37348,G37349,G37350,G37351,G37352,G37353,G37354,G37355,G37356,G37357,G37358,G37359,G37360,
       G37361,G37362,G37363,G37364,G37365,G37366,G37367,G37368,G37369,G37370,G37371,G37372,G37373,G37374,G37375,G37376,G37377,G37378,G37379,G37380,
       G37381,G37382,G37383,G37384,G37385,G37386,G37387,G37388,G37389,G37390,G37391,G37392,G37393,G37394,G37395,G37396,G37397,G37398,G37399,G37400,
       G37401,G37402,G37403,G37404,G37405,G37406,G37407,G37408,G37409,G37410,G37411,G37412,G37413,G37414,G37415,G37416,G37417,G37418,G37419,G37420,
       G37421,G37422,G37423,G37424,G37425,G37426,G37427,G37428,G37429,G37430,G37431,G37432,G37433,G37434,G37435,G37436,G37437,G37438,G37439,G37440,
       G37441,G37442,G37443,G37444,G37445,G37446,G37447,G37448,G37449,G37450,G37451,G37452,G37453,G37454,G37455,G37456,G37457,G37458,G37459,G37460,
       G37461,G37462,G37463,G37464,G37465,G37466,G37467,G37468,G37469,G37470,G37471,G37472,G37473,G37474,G37475,G37476,G37477,G37478,G37479,G37480,
       G37481,G37482,G37483,G37484,G37485,G37486,G37487,G37488,G37489,G37490,G37491,G37492,G37493,G37494,G37495,G37496,G37497,G37498,G37499,G37500,
       G37501,G37502,G37503,G37504,G37505,G37506,G37507,G37508,G37509,G37510,G37511,G37512,G37513,G37514,G37515,G37516,G37517,G37518,G37519,G37520,
       G37521,G37522,G37523,G37524,G37525,G37526,G37527,G37528,G37529,G37530,G37531,G37532,G37533,G37534,G37535,G37536,G37537,G37538,G37539,G37540,
       G37541,G37542,G37543,G37544,G37545,G37546,G37547,G37548,G37549,G37550,G37551,G37552,G37553,G37554,G37555,G37556,G37557,G37558,G37559,G37560,
       G37561,G37562,G37563,G37564,G37565,G37566,G37567,G37568,G37569,G37570,G37571,G37572,G37573,G37574,G37575,G37576,G37577,G37578,G37579,G37580,
       G37581,G37582,G37583,G37584,G37585,G37586,G37587,G37588,G37589,G37590,G37591,G37592,G37593,G37594,G37595,G37596,G37597,G37598,G37599,G37600,
       G37601,G37602,G37603,G37604,G37605,G37606,G37607,G37608,G37609,G37610,G37611,G37612,G37613,G37614,G37615,G37616,G37617,G37618,G37619,G37620,
       G37621,G37622,G37623,G37624,G37625,G37626,G37627,G37628,G37629,G37630,G37631,G37632,G37633,G37634,G37635,G37636,G37637,G37638,G37639,G37640,
       G37641,G37642,G37643,G37644,G37645,G37646,G37647,G37648,G37649,G37650,G37651,G37652,G37653,G37654,G37655,G37656,G37657,G37658,G37659,G37660,
       G37661,G37662,G37663,G37664,G37665,G37666,G37667,G37668,G37669,G37670,G37671,G37672,G37673,G37674,G37675,G37676,G37677,G37678,G37679,G37680,
       G37681,G37682,G37683,G37684,G37685,G37686,G37687,G37688,G37689,G37690,G37691,G37692,G37693,G37694,G37695,G37696,G37697,G37698,G37699,G37700,
       G37701,G37702,G37703,G37704,G37705,G37706,G37707,G37708,G37709,G37710,G37711,G37712,G37713,G37714,G37715,G37716,G37717,G37718,G37719,G37720,
       G37721,G37722,G37723,G37724,G37725,G37726,G37727,G37728,G37729,G37730,G37731,G37732,G37733,G37734,G37735,G37736,G37737,G37738,G37739,G37740,
       G37741,G37742,G37743,G37744,G37745,G37746,G37747,G37748,G37749,G37750,G37751,G37752,G37753,G37754,G37755,G37756,G37757,G37758,G37759,G37760,
       G37761,G37762,G37763,G37764,G37765,G37766,G37767,G37768,G37769,G37770,G37771,G37772,G37773,G37774,G37775,G37776,G37777,G37778,G37779,G37780,
       G37781,G37782,G37783,G37784,G37785,G37786,G37787,G37788,G37789,G37790,G37791,G37792,G37793,G37794,G37795,G37796,G37797,G37798,G37799,G37800,
       G37801,G37802,G37803,G37804,G37805,G37806,G37807,G37808,G37809,G37810,G37811,G37812,G37813,G37814,G37815,G37816,G37817,G37818,G37819,G37820,
       G37821,G37822,G37823,G37824,G37825,G37826,G37827,G37828,G37829,G37830,G37831,G37832,G37833,G37834,G37835,G37836,G37837,G37838,G37839,G37840,
       G37841,G37842,G37843,G37844,G37845,G37846,G37847,G37848,G37849,G37850,G37851,G37852,G37853,G37854,G37855,G37856,G37857,G37858,G37859,G37860,
       G37861,G37862,G37863,G37864,G37865,G37866,G37867,G37868,G37869,G37870,G37871,G37872,G37873,G37874,G37875,G37876,G37877,G37878,G37879,G37880,
       G37881,G37882,G37883,G37884,G37885,G37886,G37887,G37888,G37889,G37890,G37891,G37892,G37893,G37894,G37895,G37896,G37897,G37898,G37899,G37900,
       G37901,G37902,G37903,G37904,G37905,G37906,G37907,G37908,G37909,G37910,G37911,G37912,G37913,G37914,G37915,G37916,G37917,G37918,G37919,G37920,
       G37921,G37922,G37923,G37924,G37925,G37926,G37927,G37928,G37929,G37930,G37931,G37932,G37933,G37934,G37935,G37936,G37937,G37938,G37939,G37940,
       G37941,G37942,G37943,G37944,G37945,G37946,G37947,G37948,G37949,G37950,G37951,G37952,G37953,G37954,G37955,G37956,G37957,G37958,G37959,G37960,
       G37961,G37962,G37963,G37964,G37965,G37966,G37967,G37968,G37969,G37970,G37971,G37972,G37973,G37974,G37975,G37976,G37977,G37978,G37979,G37980,
       G37981,G37982,G37983,G37984,G37985,G37986,G37987,G37988,G37989,G37990,G37991,G37992,G37993,G37994,G37995,G37996,G37997,G37998,G37999,G38000,
       G38001,G38002,G38003,G38004,G38005,G38006,G38007,G38008,G38009,G38010,G38011,G38012,G38013,G38014,G38015,G38016,G38017,G38018,G38019,G38020,
       G38021,G38022,G38023,G38024,G38025,G38026,G38027,G38028,G38029,G38030,G38031,G38032,G38033,G38034,G38035,G38036,G38037,G38038,G38039,G38040,
       G38041,G38042,G38043,G38044,G38045,G38046,G38047,G38048,G38049,G38050,G38051,G38052,G38053,G38054,G38055,G38056,G38057,G38058,G38059,G38060,
       G38061,G38062,G38063,G38064,G38065,G38066,G38067,G38068,G38069,G38070,G38071,G38072,G38073,G38074,G38075,G38076,G38077,G38078,G38079,G38080,
       G38081,G38082,G38083,G38084,G38085,G38086,G38087,G38088,G38089,G38090,G38091,G38092,G38093,G38094,G38095,G38096,G38097,G38098,G38099,G38100,
       G38101,G38102,G38103,G38104,G38105,G38106,G38107,G38108,G38109,G38110,G38111,G38112,G38113,G38114,G38115,G38116,G38117,G38118,G38119,G38120,
       G38121,G38122,G38123,G38124,G38125,G38126,G38127,G38128,G38129,G38130,G38131,G38132,G38133,G38134,G38135,G38136,G38137,G38138,G38139,G38140,
       G38141,G38142,G38143,G38144,G38145,G38146,G38147,G38148,G38149,G38150,G38151,G38152,G38153,G38154,G38155,G38156,G38157,G38158,G38159,G38160,
       G38161,G38162,G38163,G38164,G38165,G38166,G38167,G38168,G38169,G38170,G38171,G38172,G38173,G38174,G38175,G38176,G38177,G38178,G38179,G38180,
       G38181,G38182,G38183,G38184,G38185,G38186,G38187,G38188,G38189,G38190,G38191,G38192,G38193,G38194,G38195,G38196,G38197,G38198,G38199,G38200,
       G38201,G38202,G38203,G38204,G38205,G38206,G38207,G38208,G38209,G38210,G38211,G38212,G38213,G38214,G38215,G38216,G38217,G38218,G38219,G38220,
       G38221,G38222,G38223,G38224,G38225,G38226,G38227,G38228,G38229,G38230,G38231,G38232,G38233,G38234,G38235,G38236,G38237,G38238,G38239,G38240,
       G38241,G38242,G38243,G38244,G38245,G38246,G38247,G38248,G38249,G38250,G38251,G38252,G38253,G38254,G38255,G38256,G38257,G38258,G38259,G38260,
       G38261,G38262,G38263,G38264,G38265,G38266,G38267,G38268,G38269,G38270,G38271,G38272,G38273,G38274,G38275,G38276,G38277,G38278,G38279,G38280,
       G38281,G38282,G38283,G38284,G38285,G38286,G38287,G38288,G38289,G38290,G38291,G38292,G38293,G38294,G38295,G38296,G38297,G38298,G38299,G38300,
       G38301,G38302,G38303,G38304,G38305,G38306,G38307,G38308,G38309,G38310,G38311,G38312,G38313,G38314,G38315,G38316,G38317,G38318,G38319,G38320,
       G38321,G38322,G38323,G38324,G38325,G38326,G38327,G38328,G38329,G38330,G38331,G38332,G38333,G38334,G38335,G38336,G38337,G38338,G38339,G38340,
       G38341,G38342,G38343,G38344,G38345,G38346,G38347,G38348,G38349,G38350,G38351,G38352,G38353,G38354,G38355,G38356,G38357,G38358,G38359,G38360,
       G38361,G38362,G38363,G38364,G38365,G38366,G38367,G38368,G38369,G38370,G38371,G38372,G38373,G38374,G38375,G38376,G38377,G38378,G38379,G38380,
       G38381,G38382,G38383,G38384,G38385,G38386,G38387,G38388,G38389,G38390,G38391,G38392,G38393,G38394,G38395,G38396,G38397,G38398,G38399,G38400,
       G38401,G38402,G38403,G38404,G38405,G38406,G38407,G38408,G38409,G38410,G38411,G38412,G38413,G38414,G38415,G38416,G38417,G38418,G38419,G38420,
       G38421,G38422,G38423,G38424,G38425,G38426,G38427,G38428,G38429,G38430,G38431,G38432,G38433,G38434,G38435,G38436,G38437,G38438,G38439,G38440,
       G38441,G38442,G38443,G38444,G38445,G38446,G38447,G38448,G38449,G38450,G38451,G38452,G38453,G38454,G38455,G38456,G38457,G38458,G38459,G38460,
       G38461,G38462,G38463,G38464,G38465,G38466,G38467,G38468,G38469,G38470,G38471,G38472,G38473,G38474,G38475,G38476,G38477,G38478,G38479,G38480,
       G38481,G38482,G38483,G38484,G38485,G38486,G38487,G38488,G38489,G38490,G38491,G38492,G38493,G38494,G38495,G38496,G38497,G38498,G38499,G38500,
       G38501,G38502,G38503,G38504,G38505,G38506,G38507,G38508,G38509,G38510,G38511,G38512,G38513,G38514,G38515,G38516,G38517,G38518,G38519,G38520,
       G38521,G38522,G38523,G38524,G38525,G38526,G38527,G38528,G38529,G38530,G38531,G38532,G38533,G38534,G38535,G38536,G38537,G38538,G38539,G38540,
       G38541,G38542,G38543,G38544,G38545,G38546,G38547,G38548,G38549,G38550,G38551,G38552,G38553,G38554,G38555,G38556,G38557,G38558,G38559,G38560,
       G38561,G38562,G38563,G38564,G38565,G38566,G38567,G38568,G38569,G38570,G38571,G38572,G38573,G38574,G38575,G38576,G38577,G38578,G38579,G38580,
       G38581,G38582,G38583,G38584,G38585,G38586,G38587,G38588,G38589,G38590,G38591,G38592,G38593,G38594,G38595,G38596,G38597,G38598,G38599,G38600,
       G38601,G38602,G38603,G38604,G38605,G38606,G38607,G38608,G38609,G38610,G38611,G38612,G38613,G38614,G38615,G38616,G38617,G38618,G38619,G38620,
       G38621,G38622,G38623,G38624,G38625,G38626,G38627,G38628,G38629,G38630,G38631,G38632,G38633,G38634,G38635,G38636,G38637,G38638,G38639,G38640,
       G38641,G38642,G38643,G38644,G38645,G38646,G38647,G38648,G38649,G38650,G38651,G38652,G38653,G38654,G38655,G38656,G38657,G38658,G38659,G38660,
       G38661,G38662,G38663,G38664,G38665,G38666,G38667,G38668,G38669,G38670,G38671,G38672,G38673,G38674,G38675,G38676,G38677,G38678,G38679,G38680,
       G38681,G38682,G38683,G38684,G38685,G38686,G38687,G38688,G38689,G38690,G38691,G38692,G38693,G38694,G38695,G38696,G38697,G38698,G38699,G38700,
       G38701,G38702,G38703,G38704,G38705,G38706,G38707,G38708,G38709,G38710,G38711,G38712,G38713,G38714,G38715,G38716,G38717,G38718,G38719,G38720,
       G38721,G38722,G38723,G38724,G38725,G38726,G38727,G38728,G38729,G38730,G38731,G38732,G38733,G38734,G38735,G38736,G38737,G38738,G38739,G38740,
       G38741,G38742,G38743,G38744,G38745,G38746,G38747,G38748,G38749,G38750,G38751,G38752,G38753,G38754,G38755,G38756,G38757,G38758,G38759,G38760,
       G38761,G38762,G38763,G38764,G38765,G38766,G38767,G38768,G38769,G38770,G38771,G38772,G38773,G38774,G38775,G38776,G38777,G38778,G38779,G38780,
       G38781,G38782,G38783,G38784,G38785,G38786,G38787,G38788,G38789,G38790,G38791,G38792,G38793,G38794,G38795,G38796,G38797,G38798,G38799,G38800,
       G38801,G38802,G38803,G38804,G38805,G38806,G38807,G38808,G38809,G38810,G38811,G38812,G38813,G38814,G38815,G38816,G38817,G38818,G38819,G38820,
       G38821,G38822,G38823,G38824,G38825,G38826,G38827,G38828,G38829,G38830,G38831,G38832,G38833,G38834,G38835,G38836,G38837,G38838,G38839,G38840,
       G38841,G38842,G38843,G38844,G38845,G38846,G38847,G38848,G38849,G38850,G38851,G38852,G38853,G38854,G38855,G38856,G38857,G38858,G38859,G38860,
       G38861,G38862,G38863,G38864,G38865,G38866,G38867,G38868,G38869,G38870,G38871,G38872,G38873,G38874,G38875,G38876,G38877,G38878,G38879,G38880,
       G38881,G38882,G38883,G38884,G38885,G38886,G38887,G38888,G38889,G38890,G38891,G38892,G38893,G38894,G38895,G38896,G38897,G38898,G38899,G38900,
       G38901,G38902,G38903,G38904,G38905,G38906,G38907,G38908,G38909,G38910,G38911,G38912,G38913,G38914,G38915,G38916,G38917,G38918,G38919,G38920,
       G38921,G38922,G38923,G38924,G38925,G38926,G38927,G38928,G38929,G38930,G38931,G38932,G38933,G38934,G38935,G38936,G38937,G38938,G38939,G38940,
       G38941,G38942,G38943,G38944,G38945,G38946,G38947,G38948,G38949,G38950,G38951,G38952,G38953,G38954,G38955,G38956,G38957,G38958,G38959,G38960,
       G38961,G38962,G38963,G38964,G38965,G38966,G38967,G38968,G38969,G38970,G38971,G38972,G38973,G38974,G38975,G38976,G38977,G38978,G38979,G38980,
       G38981,G38982,G38983,G38984,G38985,G38986,G38987,G38988,G38989,G38990,G38991,G38992,G38993,G38994,G38995,G38996,G38997,G38998,G38999,G39000,
       G39001,G39002,G39003,G39004,G39005,G39006,G39007,G39008,G39009,G39010,G39011,G39012,G39013,G39014,G39015,G39016,G39017,G39018,G39019,G39020,
       G39021,G39022,G39023,G39024,G39025,G39026,G39027,G39028,G39029,G39030,G39031,G39032,G39033,G39034,G39035,G39036,G39037,G39038,G39039,G39040,
       G39041,G39042,G39043,G39044,G39045,G39046,G39047,G39048,G39049,G39050,G39051,G39052,G39053,G39054,G39055,G39056,G39057,G39058,G39059,G39060,
       G39061,G39062,G39063,G39064,G39065,G39066,G39067,G39068,G39069,G39070,G39071,G39072,G39073,G39074,G39075,G39076,G39077,G39078,G39079,G39080,
       G39081,G39082,G39083,G39084,G39085,G39086,G39087,G39088,G39089,G39090,G39091,G39092,G39093,G39094,G39095,G39096,G39097,G39098,G39099,G39100,
       G39101,G39102,G39103,G39104,G39105,G39106,G39107,G39108,G39109,G39110,G39111,G39112,G39113,G39114,G39115,G39116,G39117,G39118,G39119,G39120,
       G39121,G39122,G39123,G39124,G39125,G39126,G39127,G39128,G39129,G39130,G39131,G39132,G39133,G39134,G39135,G39136,G39137,G39138,G39139,G39140,
       G39141,G39142,G39143,G39144,G39145,G39146,G39147,G39148,G39149,G39150,G39151,G39152,G39153,G39154,G39155,G39156,G39157,G39158,G39159,G39160,
       G39161,G39162,G39163,G39164,G39165,G39166,G39167,G39168,G39169,G39170,G39171,G39172,G39173,G39174,G39175,G39176,G39177,G39178,G39179,G39180,
       G39181,G39182,G39183,G39184,G39185,G39186,G39187,G39188,G39189,G39190,G39191,G39192,G39193,G39194,G39195,G39196,G39197,G39198,G39199,G39200,
       G39201,G39202,G39203,G39204,G39205,G39206,G39207,G39208,G39209,G39210,G39211,G39212,G39213,G39214,G39215,G39216,G39217,G39218,G39219,G39220,
       G39221,G39222,G39223,G39224,G39225,G39226,G39227,G39228,G39229,G39230,G39231,G39232,G39233,G39234,G39235,G39236,G39237,G39238,G39239,G39240,
       G39241,G39242,G39243,G39244,G39245,G39246,G39247,G39248,G39249,G39250,G39251,G39252,G39253,G39254,G39255,G39256,G39257,G39258,G39259,G39260,
       G39261,G39262,G39263,G39264,G39265,G39266,G39267,G39268,G39269,G39270,G39271,G39272,G39273,G39274,G39275,G39276,G39277,G39278,G39279,G39280,
       G39281,G39282,G39283,G39284,G39285,G39286,G39287,G39288,G39289,G39290,G39291,G39292,G39293,G39294,G39295,G39296,G39297,G39298,G39299,G39300,
       G39301,G39302,G39303,G39304,G39305,G39306,G39307,G39308,G39309,G39310,G39311,G39312,G39313,G39314,G39315,G39316,G39317,G39318,G39319,G39320,
       G39321,G39322,G39323,G39324,G39325,G39326,G39327,G39328,G39329,G39330,G39331,G39332,G39333,G39334,G39335,G39336,G39337,G39338,G39339,G39340,
       G39341,G39342,G39343,G39344,G39345,G39346,G39347,G39348,G39349,G39350,G39351,G39352,G39353,G39354,G39355,G39356,G39357,G39358,G39359,G39360,
       G39361,G39362,G39363,G39364,G39365,G39366,G39367,G39368,G39369,G39370,G39371,G39372,G39373,G39374,G39375,G39376,G39377,G39378,G39379,G39380,
       G39381,G39382,G39383,G39384,G39385,G39386,G39387,G39388,G39389,G39390,G39391,G39392,G39393,G39394,G39395,G39396,G39397,G39398,G39399,G39400,
       G39401,G39402,G39403,G39404,G39405,G39406,G39407,G39408,G39409,G39410,G39411,G39412,G39413,G39414,G39415,G39416,G39417,G39418,G39419,G39420,
       G39421,G39422,G39423,G39424,G39425,G39426,G39427,G39428,G39429,G39430,G39431,G39432,G39433,G39434,G39435,G39436,G39437,G39438,G39439,G39440,
       G39441,G39442,G39443,G39444,G39445,G39446,G39447,G39448,G39449,G39450,G39451,G39452,G39453,G39454,G39455,G39456,G39457,G39458,G39459,G39460,
       G39461,G39462,G39463,G39464,G39465,G39466,G39467,G39468,G39469,G39470,G39471,G39472,G39473,G39474,G39475,G39476,G39477,G39478,G39479,G39480,
       G39481,G39482,G39483,G39484,G39485,G39486,G39487,G39488,G39489,G39490,G39491,G39492,G39493,G39494,G39495,G39496,G39497,G39498,G39499,G39500,
       G39501,G39502,G39503,G39504,G39505,G39506,G39507,G39508,G39509,G39510,G39511,G39512,G39513,G39514,G39515,G39516,G39517,G39518,G39519,G39520,
       G39521,G39522,G39523,G39524,G39525,G39526,G39527,G39528,G39529,G39530,G39531,G39532,G39533,G39534,G39535,G39536,G39537,G39538,G39539,G39540,
       G39541,G39542,G39543,G39544,G39545,G39546,G39547,G39548,G39549,G39550,G39551,G39552,G39553,G39554,G39555,G39556,G39557,G39558,G39559,G39560,
       G39561,G39562,G39563,G39564,G39565,G39566,G39567,G39568,G39569,G39570,G39571,G39572,G39573,G39574,G39575,G39576,G39577,G39578,G39579,G39580,
       G39581,G39582,G39583,G39584,G39585,G39586,G39587,G39588,G39589,G39590,G39591,G39592,G39593,G39594,G39595,G39596,G39597,G39598,G39599,G39600,
       G39601,G39602,G39603,G39604,G39605,G39606,G39607,G39608,G39609,G39610,G39611,G39612,G39613,G39614,G39615,G39616,G39617,G39618,G39619,G39620,
       G39621,G39622,G39623,G39624,G39625,G39626,G39627,G39628,G39629,G39630,G39631,G39632,G39633,G39634,G39635,G39636,G39637,G39638,G39639,G39640,
       G39641,G39642,G39643,G39644,G39645,G39646,G39647,G39648,G39649,G39650,G39651,G39652,G39653,G39654,G39655,G39656,G39657,G39658,G39659,G39660,
       G39661,G39662,G39663,G39664,G39665,G39666,G39667,G39668,G39669,G39670,G39671,G39672,G39673,G39674,G39675,G39676,G39677,G39678,G39679,G39680,
       G39681,G39682,G39683,G39684,G39685,G39686,G39687,G39688,G39689,G39690,G39691,G39692,G39693,G39694,G39695,G39696,G39697,G39698,G39699,G39700,
       G39701,G39702,G39703,G39704,G39705,G39706,G39707,G39708,G39709,G39710,G39711,G39712,G39713,G39714,G39715,G39716,G39717,G39718,G39719,G39720,
       G39721,G39722,G39723,G39724,G39725,G39726,G39727,G39728,G39729,G39730,G39731,G39732,G39733,G39734,G39735,G39736,G39737,G39738,G39739,G39740,
       G39741,G39742,G39743,G39744,G39745,G39746,G39747,G39748,G39749,G39750,G39751,G39752,G39753,G39754,G39755,G39756,G39757,G39758,G39759,G39760,
       G39761,G39762,G39763,G39764,G39765,G39766,G39767,G39768,G39769,G39770,G39771,G39772,G39773,G39774,G39775,G39776,G39777,G39778,G39779,G39780,
       G39781,G39782,G39783,G39784,G39785,G39786,G39787,G39788,G39789,G39790,G39791,G39792,G39793,G39794,G39795,G39796,G39797,G39798,G39799,G39800,
       G39801,G39802,G39803,G39804,G39805,G39806,G39807,G39808,G39809,G39810,G39811,G39812,G39813,G39814,G39815,G39816,G39817,G39818,G39819,G39820,
       G39821,G39822,G39823,G39824,G39825,G39826,G39827,G39828,G39829,G39830,G39831,G39832,G39833,G39834,G39835,G39836,G39837,G39838,G39839,G39840,
       G39841,G39842,G39843,G39844,G39845,G39846,G39847,G39848,G39849,G39850,G39851,G39852,G39853,G39854,G39855,G39856,G39857,G39858,G39859,G39860,
       G39861,G39862,G39863,G39864,G39865,G39866,G39867,G39868,G39869,G39870,G39871,G39872,G39873,G39874,G39875,G39876,G39877,G39878,G39879,G39880,
       G39881,G39882,G39883,G39884,G39885,G39886,G39887,G39888,G39889,G39890,G39891,G39892,G39893,G39894,G39895,G39896,G39897,G39898,G39899,G39900,
       G39901,G39902,G39903,G39904,G39905,G39906,G39907,G39908,G39909,G39910,G39911,G39912,G39913,G39914,G39915,G39916,G39917,G39918,G39919,G39920,
       G39921,G39922,G39923,G39924,G39925,G39926,G39927,G39928,G39929,G39930,G39931,G39932,G39933,G39934,G39935,G39936,G39937,G39938,G39939,G39940,
       G39941,G39942,G39943,G39944,G39945,G39946,G39947,G39948,G39949,G39950,G39951,G39952,G39953,G39954,G39955,G39956,G39957,G39958,G39959,G39960,
       G39961,G39962,G39963,G39964,G39965,G39966,G39967,G39968,G39969,G39970,G39971,G39972,G39973,G39974,G39975,G39976,G39977,G39978,G39979,G39980,
       G39981,G39982,G39983,G39984,G39985,G39986,G39987,G39988,G39989,G39990,G39991,G39992,G39993,G39994,G39995,G39996,G39997,G39998,G39999,G40000,
       G40001,G40002,G40003,G40004,G40005,G40006,G40007,G40008,G40009,G40010,G40011,G40012,G40013,G40014,G40015,G40016,G40017,G40018,G40019,G40020,
       G40021,G40022,G40023,G40024,G40025,G40026,G40027,G40028,G40029,G40030,G40031,G40032,G40033,G40034,G40035,G40036,G40037,G40038,G40039,G40040,
       G40041,G40042,G40043,G40044,G40045,G40046,G40047,G40048,G40049,G40050,G40051,G40052,G40053,G40054,G40055,G40056,G40057,G40058,G40059,G40060,
       G40061,G40062,G40063,G40064,G40065,G40066,G40067,G40068,G40069,G40070,G40071,G40072,G40073,G40074,G40075,G40076,G40077,G40078,G40079,G40080,
       G40081,G40082,G40083,G40084,G40085,G40086,G40087,G40088,G40089,G40090,G40091,G40092,G40093,G40094,G40095,G40096,G40097,G40098,G40099,G40100,
       G40101,G40102,G40103,G40104,G40105,G40106,G40107,G40108,G40109,G40110,G40111,G40112,G40113,G40114,G40115,G40116,G40117,G40118,G40119,G40120,
       G40121,G40122,G40123,G40124,G40125,G40126,G40127,G40128,G40129,G40130,G40131,G40132,G40133,G40134,G40135,G40136,G40137,G40138,G40139,G40140,
       G40141,G40142,G40143,G40144,G40145,G40146,G40147,G40148,G40149,G40150,G40151,G40152,G40153,G40154,G40155,G40156,G40157,G40158,G40159,G40160,
       G40161,G40162,G40163,G40164,G40165,G40166,G40167,G40168,G40169,G40170,G40171,G40172,G40173,G40174,G40175,G40176,G40177,G40178,G40179,G40180,
       G40181,G40182,G40183,G40184,G40185,G40186,G40187,G40188,G40189,G40190,G40191,G40192,G40193,G40194,G40195,G40196,G40197,G40198,G40199,G40200,
       G40201,G40202,G40203,G40204,G40205,G40206,G40207,G40208,G40209,G40210,G40211,G40212,G40213,G40214,G40215,G40216,G40217,G40218,G40219,G40220,
       G40221,G40222,G40223,G40224,G40225,G40226,G40227,G40228,G40229,G40230,G40231,G40232,G40233,G40234,G40235,G40236,G40237,G40238,G40239,G40240,
       G40241,G40242,G40243,G40244,G40245,G40246,G40247,G40248,G40249,G40250,G40251,G40252,G40253,G40254,G40255,G40256,G40257,G40258,G40259,G40260,
       G40261,G40262,G40263,G40264,G40265,G40266,G40267,G40268,G40269,G40270,G40271,G40272,G40273,G40274,G40275,G40276,G40277,G40278,G40279,G40280,
       G40281,G40282,G40283,G40284,G40285,G40286,G40287,G40288,G40289,G40290,G40291,G40292,G40293,G40294,G40295,G40296,G40297,G40298,G40299,G40300,
       G40301,G40302,G40303,G40304,G40305,G40306,G40307,G40308,G40309,G40310,G40311,G40312,G40313,G40314,G40315,G40316,G40317,G40318,G40319,G40320,
       G40321,G40322,G40323,G40324,G40325,G40326,G40327,G40328,G40329,G40330,G40331,G40332,G40333,G40334,G40335,G40336,G40337,G40338,G40339,G40340,
       G40341,G40342,G40343,G40344,G40345,G40346,G40347,G40348,G40349,G40350,G40351,G40352,G40353,G40354,G40355,G40356,G40357,G40358,G40359,G40360,
       G40361,G40362,G40363,G40364,G40365,G40366,G40367,G40368,G40369,G40370,G40371,G40372,G40373,G40374,G40375,G40376,G40377,G40378,G40379,G40380,
       G40381,G40382,G40383,G40384,G40385,G40386,G40387,G40388,G40389,G40390,G40391,G40392,G40393,G40394,G40395,G40396,G40397,G40398,G40399,G40400,
       G40401,G40402,G40403,G40404,G40405,G40406,G40407,G40408,G40409,G40410,G40411,G40412,G40413,G40414,G40415,G40416,G40417,G40418,G40419,G40420,
       G40421,G40422,G40423,G40424,G40425,G40426,G40427,G40428,G40429,G40430,G40431,G40432,G40433,G40434,G40435,G40436,G40437,G40438,G40439,G40440,
       G40441,G40442,G40443,G40444,G40445,G40446,G40447,G40448,G40449,G40450,G40451,G40452,G40453,G40454,G40455,G40456,G40457,G40458,G40459,G40460,
       G40461,G40462,G40463,G40464,G40465,G40466,G40467,G40468,G40469,G40470,G40471,G40472,G40473,G40474,G40475,G40476,G40477,G40478,G40479,G40480,
       G40481,G40482,G40483,G40484,G40485,G40486,G40487,G40488,G40489,G40490,G40491,G40492,G40493,G40494,G40495,G40496,G40497,G40498,G40499,G40500,
       G40501,G40502,G40503,G40504,G40505,G40506,G40507,G40508,G40509,G40510,G40511,G40512,G40513,G40514,G40515,G40516,G40517,G40518,G40519,G40520,
       G40521,G40522,G40523,G40524,G40525,G40526,G40527,G40528,G40529,G40530,G40531,G40532,G40533,G40534,G40535,G40536,G40537,G40538,G40539,G40540,
       G40541,G40542,G40543,G40544,G40545,G40546,G40547,G40548,G40549,G40550,G40551,G40552,G40553,G40554,G40555,G40556,G40557,G40558,G40559,G40560,
       G40561,G40562,G40563,G40564,G40565,G40566,G40567,G40568,G40569,G40570,G40571,G40572,G40573,G40574,G40575,G40576,G40577,G40578,G40579,G40580,
       G40581,G40582,G40583,G40584,G40585,G40586,G40587,G40588,G40589,G40590,G40591,G40592,G40593,G40594,G40595,G40596,G40597,G40598,G40599,G40600,
       G40601,G40602,G40603,G40604,G40605,G40606,G40607,G40608,G40609,G40610,G40611,G40612,G40613,G40614,G40615,G40616,G40617,G40618,G40619,G40620,
       G40621,G40622,G40623,G40624,G40625,G40626,G40627,G40628,G40629,G40630,G40631,G40632,G40633,G40634,G40635,G40636,G40637,G40638,G40639,G40640,
       G40641,G40642,G40643,G40644,G40645,G40646,G40647,G40648,G40649,G40650,G40651,G40652,G40653,G40654,G40655,G40656,G40657,G40658,G40659,G40660,
       G40661,G40662,G40663,G40664,G40665,G40666,G40667,G40668,G40669,G40670,G40671,G40672,G40673,G40674,G40675,G40676,G40677,G40678,G40679,G40680,
       G40681,G40682,G40683,G40684,G40685,G40686,G40687,G40688,G40689,G40690,G40691,G40692,G40693,G40694,G40695,G40696,G40697,G40698,G40699,G40700,
       G40701,G40702,G40703,G40704,G40705,G40706,G40707,G40708,G40709,G40710,G40711,G40712,G40713,G40714,G40715,G40716,G40717,G40718,G40719,G40720,
       G40721,G40722,G40723,G40724,G40725,G40726,G40727,G40728,G40729,G40730,G40731,G40732,G40733,G40734,G40735,G40736,G40737,G40738,G40739,G40740,
       G40741,G40742,G40743,G40744,G40745,G40746,G40747,G40748,G40749,G40750,G40751,G40752,G40753,G40754,G40755,G40756,G40757,G40758,G40759,G40760,
       G40761,G40762,G40763,G40764,G40765,G40766,G40767,G40768,G40769,G40770,G40771,G40772,G40773,G40774,G40775,G40776,G40777,G40778,G40779,G40780,
       G40781,G40782,G40783,G40784,G40785,G40786,G40787,G40788,G40789,G40790,G40791,G40792,G40793,G40794,G40795,G40796,G40797,G40798,G40799,G40800,
       G40801,G40802,G40803,G40804,G40805,G40806,G40807,G40808,G40809,G40810,G40811,G40812,G40813,G40814,G40815,G40816,G40817,G40818,G40819,G40820,
       G40821,G40822,G40823,G40824,G40825,G40826,G40827,G40828,G40829,G40830,G40831,G40832,G40833,G40834,G40835,G40836,G40837,G40838,G40839,G40840,
       G40841,G40842,G40843,G40844,G40845,G40846,G40847,G40848,G40849,G40850,G40851,G40852,G40853,G40854,G40855,G40856,G40857,G40858,G40859,G40860,
       G40861,G40862,G40863,G40864,G40865,G40866,G40867,G40868,G40869,G40870,G40871,G40872,G40873,G40874,G40875,G40876,G40877,G40878,G40879,G40880,
       G40881,G40882,G40883,G40884,G40885,G40886,G40887,G40888,G40889,G40890,G40891,G40892,G40893,G40894,G40895,G40896,G40897,G40898,G40899,G40900,
       G40901,G40902,G40903,G40904,G40905,G40906,G40907,G40908,G40909,G40910,G40911,G40912,G40913,G40914,G40915,G40916,G40917,G40918,G40919,G40920,
       G40921,G40922,G40923,G40924,G40925,G40926,G40927,G40928,G40929,G40930,G40931,G40932,G40933,G40934,G40935,G40936,G40937,G40938,G40939,G40940,
       G40941,G40942,G40943,G40944,G40945,G40946,G40947,G40948,G40949,G40950,G40951,G40952,G40953,G40954,G40955,G40956,G40957,G40958,G40959,G40960,
       G40961,G40962,G40963,G40964,G40965,G40966,G40967,G40968,G40969,G40970,G40971,G40972,G40973,G40974,G40975,G40976,G40977,G40978,G40979,G40980,
       G40981,G40982,G40983,G40984,G40985,G40986,G40987,G40988,G40989,G40990,G40991,G40992,G40993,G40994,G40995,G40996,G40997,G40998,G40999,G41000,
       G41001,G41002,G41003,G41004,G41005,G41006,G41007,G41008,G41009,G41010,G41011,G41012,G41013,G41014,G41015,G41016,G41017,G41018,G41019,G41020,
       G41021,G41022,G41023,G41024,G41025,G41026,G41027,G41028,G41029,G41030,G41031,G41032,G41033,G41034,G41035,G41036,G41037,G41038,G41039,G41040,
       G41041,G41042,G41043,G41044,G41045,G41046,G41047,G41048,G41049,G41050,G41051,G41052,G41053,G41054,G41055,G41056,G41057,G41058,G41059,G41060,
       G41061,G41062,G41063,G41064,G41065,G41066,G41067,G41068,G41069,G41070,G41071,G41072,G41073,G41074,G41075,G41076,G41077,G41078,G41079,G41080,
       G41081,G41082,G41083,G41084,G41085,G41086,G41087,G41088,G41089,G41090,G41091,G41092,G41093,G41094,G41095,G41096,G41097,G41098,G41099,G41100,
       G41101,G41102,G41103,G41104,G41105,G41106,G41107,G41108,G41109,G41110,G41111,G41112,G41113,G41114,G41115,G41116,G41117,G41118,G41119,G41120,
       G41121,G41122,G41123,G41124,G41125,G41126,G41127,G41128,G41129,G41130,G41131,G41132,G41133,G41134,G41135,G41136,G41137,G41138,G41139,G41140,
       G41141,G41142,G41143,G41144,G41145,G41146,G41147,G41148,G41149,G41150,G41151,G41152,G41153,G41154,G41155,G41156,G41157,G41158,G41159,G41160,
       G41161,G41162,G41163,G41164,G41165,G41166,G41167,G41168,G41169,G41170,G41171,G41172,G41173,G41174,G41175,G41176,G41177,G41178,G41179,G41180,
       G41181,G41182,G41183,G41184,G41185,G41186,G41187,G41188,G41189,G41190,G41191,G41192,G41193,G41194,G41195,G41196,G41197,G41198,G41199,G41200,
       G41201,G41202,G41203,G41204,G41205,G41206,G41207,G41208,G41209,G41210,G41211,G41212,G41213,G41214,G41215,G41216,G41217,G41218,G41219,G41220,
       G41221,G41222,G41223,G41224,G41225,G41226,G41227,G41228,G41229,G41230,G41231,G41232,G41233,G41234,G41235,G41236,G41237,G41238,G41239,G41240,
       G41241,G41242,G41243,G41244,G41245,G41246,G41247,G41248,G41249,G41250,G41251,G41252,G41253,G41254,G41255,G41256,G41257,G41258,G41259,G41260,
       G41261,G41262,G41263,G41264,G41265,G41266,G41267,G41268,G41269,G41270,G41271,G41272,G41273,G41274,G41275,G41276,G41277,G41278,G41279,G41280,
       G41281,G41282,G41283,G41284,G41285,G41286,G41287,G41288,G41289,G41290,G41291,G41292,G41293,G41294,G41295,G41296,G41297,G41298,G41299,G41300,
       G41301,G41302,G41303,G41304,G41305,G41306,G41307,G41308,G41309,G41310,G41311,G41312,G41313,G41314,G41315,G41316,G41317,G41318,G41319,G41320,
       G41321,G41322,G41323,G41324,G41325,G41326,G41327,G41328,G41329,G41330,G41331,G41332,G41333,G41334,G41335,G41336,G41337,G41338,G41339,G41340,
       G41341,G41342,G41343,G41344,G41345,G41346,G41347,G41348,G41349,G41350,G41351,G41352,G41353,G41354,G41355,G41356,G41357,G41358,G41359,G41360,
       G41361,G41362,G41363,G41364,G41365,G41366,G41367,G41368,G41369,G41370,G41371,G41372,G41373,G41374,G41375,G41376,G41377,G41378,G41379,G41380,
       G41381,G41382,G41383,G41384,G41385,G41386,G41387,G41388,G41389,G41390,G41391,G41392,G41393,G41394,G41395,G41396,G41397,G41398,G41399,G41400,
       G41401,G41402,G41403,G41404,G41405,G41406,G41407,G41408,G41409,G41410,G41411,G41412,G41413,G41414,G41415,G41416,G41417,G41418,G41419,G41420,
       G41421,G41422,G41423,G41424,G41425,G41426,G41427,G41428,G41429,G41430,G41431,G41432,G41433,G41434,G41435,G41436,G41437,G41438,G41439,G41440,
       G41441,G41442,G41443,G41444,G41445,G41446,G41447,G41448,G41449,G41450,G41451,G41452,G41453,G41454,G41455,G41456,G41457,G41458,G41459,G41460,
       G41461,G41462,G41463,G41464,G41465,G41466,G41467,G41468,G41469,G41470,G41471,G41472,G41473,G41474,G41475,G41476,G41477,G41478,G41479,G41480,
       G41481,G41482,G41483,G41484,G41485,G41486,G41487,G41488,G41489,G41490,G41491,G41492,G41493,G41494,G41495,G41496,G41497,G41498,G41499,G41500,
       G41501,G41502,G41503,G41504,G41505,G41506,G41507,G41508,G41509,G41510,G41511,G41512,G41513,G41514,G41515,G41516,G41517,G41518,G41519,G41520,
       G41521,G41522,G41523,G41524,G41525,G41526,G41527,G41528,G41529,G41530,G41531,G41532,G41533,G41534,G41535,G41536,G41537,G41538,G41539,G41540,
       G41541,G41542,G41543,G41544,G41545,G41546,G41547,G41548,G41549,G41550,G41551,G41552,G41553,G41554,G41555,G41556,G41557,G41558,G41559,G41560,
       G41561,G41562,G41563,G41564,G41565,G41566,G41567,G41568,G41569,G41570,G41571,G41572,G41573,G41574,G41575,G41576,G41577,G41578,G41579,G41580,
       G41581,G41582,G41583,G41584,G41585,G41586,G41587,G41588,G41589,G41590,G41591,G41592,G41593,G41594,G41595,G41596,G41597,G41598,G41599,G41600,
       G41601,G41602,G41603,G41604,G41605,G41606,G41607,G41608,G41609,G41610,G41611,G41612,G41613,G41614,G41615,G41616,G41617,G41618,G41619,G41620,
       G41621,G41622,G41623,G41624,G41625,G41626,G41627,G41628,G41629,G41630,G41631,G41632,G41633,G41634,G41635,G41636,G41637,G41638,G41639,G41640,
       G41641,G41642,G41643,G41644,G41645,G41646,G41647,G41648,G41649,G41650,G41651,G41652,G41653,G41654,G41655,G41656,G41657,G41658,G41659,G41660,
       G41661,G41662,G41663,G41664,G41665,G41666,G41667,G41668,G41669,G41670,G41671,G41672,G41673,G41674,G41675,G41676,G41677,G41678,G41679,G41680,
       G41681,G41682,G41683,G41684,G41685,G41686,G41687,G41688,G41689,G41690,G41691,G41692,G41693,G41694,G41695,G41696,G41697,G41698,G41699,G41700,
       G41701,G41702,G41703,G41704,G41705,G41706,G41707,G41708,G41709,G41710,G41711,G41712,G41713,G41714,G41715,G41716,G41717,G41718,G41719,G41720,
       G41721,G41722,G41723,G41724,G41725,G41726,G41727,G41728,G41729,G41730,G41731,G41732,G41733,G41734,G41735,G41736,G41737,G41738,G41739,G41740,
       G41741,G41742,G41743,G41744,G41745,G41746,G41747,G41748,G41749,G41750,G41751,G41752,G41753,G41754,G41755,G41756,G41757,G41758,G41759,G41760,
       G41761,G41762,G41763,G41764,G41765,G41766,G41767,G41768,G41769,G41770,G41771,G41772,G41773,G41774,G41775,G41776,G41777,G41778,G41779,G41780,
       G41781,G41782,G41783,G41784,G41785,G41786,G41787,G41788,G41789,G41790,G41791,G41792,G41793,G41794,G41795,G41796,G41797,G41798,G41799,G41800,
       G41801,G41802,G41803,G41804,G41805,G41806,G41807,G41808,G41809,G41810,G41811,G41812,G41813,G41814,G41815,G41816,G41817,G41818,G41819,G41820,
       G41821,G41822,G41823,G41824,G41825,G41826,G41827,G41828,G41829,G41830,G41831,G41832,G41833,G41834,G41835,G41836,G41837,G41838,G41839,G41840,
       G41841,G41842,G41843,G41844,G41845,G41846,G41847,G41848,G41849,G41850,G41851,G41852,G41853,G41854,G41855,G41856,G41857,G41858,G41859,G41860,
       G41861,G41862,G41863,G41864,G41865,G41866,G41867,G41868,G41869,G41870,G41871,G41872,G41873,G41874,G41875,G41876,G41877,G41878,G41879,G41880,
       G41881,G41882,G41883,G41884,G41885,G41886,G41887,G41888,G41889,G41890,G41891,G41892,G41893,G41894,G41895,G41896,G41897,G41898,G41899,G41900,
       G41901,G41902,G41903,G41904,G41905,G41906,G41907,G41908,G41909,G41910,G41911,G41912,G41913,G41914,G41915,G41916,G41917,G41918,G41919,G41920,
       G41921,G41922,G41923,G41924,G41925,G41926,G41927,G41928,G41929,G41930,G41931,G41932,G41933,G41934,G41935,G41936,G41937,G41938,G41939,G41940,
       G41941,G41942,G41943,G41944,G41945,G41946,G41947,G41948,G41949,G41950,G41951,G41952,G41953,G41954,G41955,G41956,G41957,G41958,G41959,G41960,
       G41961,G41962,G41963,G41964,G41965,G41966,G41967,G41968,G41969,G41970,G41971,G41972,G41973,G41974,G41975,G41976,G41977,G41978,G41979,G41980,
       G41981,G41982,G41983,G41984,G41985,G41986,G41987,G41988,G41989,G41990,G41991,G41992,G41993,G41994,G41995,G41996,G41997,G41998,G41999,G42000,
       G42001,G42002,G42003,G42004,G42005,G42006,G42007,G42008,G42009,G42010,G42011,G42012,G42013,G42014,G42015,G42016,G42017,G42018,G42019,G42020,
       G42021,G42022,G42023,G42024,G42025,G42026,G42027,G42028,G42029,G42030,G42031,G42032,G42033,G42034,G42035,G42036,G42037,G42038,G42039,G42040,
       G42041,G42042,G42043,G42044,G42045,G42046,G42047,G42048,G42049,G42050,G42051,G42052,G42053,G42054,G42055,G42056,G42057,G42058,G42059,G42060,
       G42061,G42062,G42063,G42064,G42065,G42066,G42067,G42068,G42069,G42070,G42071,G42072,G42073,G42074,G42075,G42076,G42077,G42078,G42079,G42080,
       G42081,G42082,G42083,G42084,G42085,G42086,G42087,G42088,G42089,G42090,G42091,G42092,G42093,G42094,G42095,G42096,G42097,G42098,G42099,G42100,
       G42101,G42102,G42103,G42104,G42105,G42106,G42107,G42108,G42109,G42110,G42111,G42112,G42113,G42114,G42115,G42116,G42117,G42118,G42119,G42120,
       G42121,G42122,G42123,G42124,G42125,G42126,G42127,G42128,G42129,G42130,G42131,G42132,G42133,G42134,G42135,G42136,G42137,G42138,G42139,G42140,
       G42141,G42142,G42143,G42144,G42145,G42146,G42147,G42148,G42149,G42150,G42151,G42152,G42153,G42154,G42155,G42156,G42157,G42158,G42159,G42160,
       G42161,G42162,G42163,G42164,G42165,G42166,G42167,G42168,G42169,G42170,G42171,G42172,G42173,G42174,G42175,G42176,G42177,G42178,G42179,G42180,
       G42181,G42182,G42183,G42184,G42185,G42186,G42187,G42188,G42189,G42190,G42191,G42192,G42193,G42194,G42195,G42196,G42197,G42198,G42199,G42200,
       G42201,G42202,G42203,G42204,G42205,G42206,G42207,G42208,G42209,G42210,G42211,G42212,G42213,G42214,G42215,G42216,G42217,G42218,G42219,G42220,
       G42221,G42222,G42223,G42224,G42225,G42226,G42227,G42228,G42229,G42230,G42231,G42232,G42233,G42234,G42235,G42236,G42237,G42238,G42239,G42240,
       G42241,G42242,G42243,G42244,G42245,G42246,G42247,G42248,G42249,G42250,G42251,G42252,G42253,G42254,G42255,G42256,G42257,G42258,G42259,G42260,
       G42261,G42262,G42263,G42264,G42265,G42266,G42267,G42268,G42269,G42270,G42271,G42272,G42273,G42274,G42275,G42276,G42277,G42278,G42279,G42280,
       G42281,G42282,G42283,G42284,G42285,G42286,G42287,G42288,G42289,G42290,G42291,G42292,G42293,G42294,G42295,G42296,G42297,G42298,G42299,G42300,
       G42301,G42302,G42303,G42304,G42305,G42306,G42307,G42308,G42309,G42310,G42311,G42312,G42313,G42314,G42315,G42316,G42317,G42318,G42319,G42320,
       G42321,G42322,G42323,G42324,G42325,G42326,G42327,G42328,G42329,G42330,G42331,G42332,G42333,G42334,G42335,G42336,G42337,G42338,G42339,G42340,
       G42341,G42342,G42343,G42344,G42345,G42346,G42347,G42348,G42349,G42350,G42351,G42352,G42353,G42354,G42355,G42356,G42357,G42358,G42359,G42360,
       G42361,G42362,G42363,G42364,G42365,G42366,G42367,G42368,G42369,G42370,G42371,G42372,G42373,G42374,G42375,G42376,G42377,G42378,G42379,G42380,
       G42381,G42382,G42383,G42384,G42385,G42386,G42387,G42388,G42389,G42390,G42391,G42392,G42393,G42394,G42395,G42396,G42397,G42398,G42399,G42400,
       G42401,G42402,G42403,G42404,G42405,G42406,G42407,G42408,G42409,G42410,G42411,G42412,G42413,G42414,G42415,G42416,G42417,G42418,G42419,G42420,
       G42421,G42422,G42423,G42424,G42425,G42426,G42427,G42428,G42429,G42430,G42431,G42432,G42433,G42434,G42435,G42436,G42437,G42438,G42439,G42440,
       G42441,G42442,G42443,G42444,G42445,G42446,G42447,G42448,G42449,G42450,G42451,G42452,G42453,G42454,G42455,G42456,G42457,G42458,G42459,G42460,
       G42461,G42462,G42463,G42464,G42465,G42466,G42467,G42468,G42469,G42470,G42471,G42472,G42473,G42474,G42475,G42476,G42477,G42478,G42479,G42480,
       G42481,G42482,G42483,G42484,G42485,G42486,G42487,G42488,G42489,G42490,G42491,G42492,G42493,G42494,G42495,G42496,G42497,G42498,G42499,G42500,
       G42501,G42502,G42503,G42504,G42505,G42506,G42507,G42508,G42509,G42510,G42511,G42512,G42513,G42514,G42515,G42516,G42517,G42518,G42519,G42520,
       G42521,G42522,G42523,G42524,G42525,G42526,G42527,G42528,G42529,G42530,G42531,G42532,G42533,G42534,G42535,G42536,G42537,G42538,G42539,G42540,
       G42541,G42542,G42543,G42544,G42545,G42546,G42547,G42548,G42549,G42550,G42551,G42552,G42553,G42554,G42555,G42556,G42557,G42558,G42559,G42560,
       G42561,G42562,G42563,G42564,G42565,G42566,G42567,G42568,G42569,G42570,G42571,G42572,G42573,G42574,G42575,G42576,G42577,G42578,G42579,G42580,
       G42581,G42582,G42583,G42584,G42585,G42586,G42587,G42588,G42589,G42590,G42591,G42592,G42593,G42594,G42595,G42596,G42597,G42598,G42599,G42600,
       G42601,G42602,G42603,G42604,G42605,G42606,G42607,G42608,G42609,G42610,G42611,G42612,G42613,G42614,G42615,G42616,G42617,G42618,G42619,G42620,
       G42621,G42622,G42623,G42624,G42625,G42626,G42627,G42628,G42629,G42630,G42631,G42632,G42633,G42634,G42635,G42636,G42637,G42638,G42639,G42640,
       G42641,G42642,G42643,G42644,G42645,G42646,G42647,G42648,G42649,G42650,G42651,G42652,G42653,G42654,G42655,G42656,G42657,G42658,G42659,G42660,
       G42661,G42662,G42663,G42664,G42665,G42666,G42667,G42668,G42669,G42670,G42671,G42672,G42673,G42674,G42675,G42676,G42677,G42678,G42679,G42680,
       G42681,G42682,G42683,G42684,G42685,G42686,G42687,G42688,G42689,G42690,G42691,G42692,G42693,G42694,G42695,G42696,G42697,G42698,G42699,G42700,
       G42701,G42702,G42703,G42704,G42705,G42706,G42707,G42708,G42709,G42710,G42711,G42712,G42713,G42714,G42715,G42716,G42717,G42718,G42719,G42720,
       G42721,G42722,G42723,G42724,G42725,G42726,G42727,G42728,G42729,G42730,G42731,G42732,G42733,G42734,G42735,G42736,G42737,G42738,G42739,G42740,
       G42741,G42742,G42743,G42744,G42745,G42746,G42747,G42748,G42749,G42750,G42751,G42752,G42753,G42754,G42755,G42756,G42757,G42758,G42759,G42760,
       G42761,G42762,G42763,G42764,G42765,G42766,G42767,G42768,G42769,G42770,G42771,G42772,G42773,G42774,G42775,G42776,G42777,G42778,G42779,G42780,
       G42781,G42782,G42783,G42784,G42785,G42786,G42787,G42788,G42789,G42790,G42791,G42792,G42793,G42794,G42795,G42796,G42797,G42798,G42799,G42800,
       G42801,G42802,G42803,G42804,G42805,G42806,G42807,G42808,G42809,G42810,G42811,G42812,G42813,G42814,G42815,G42816,G42817,G42818,G42819,G42820,
       G42821,G42822,G42823,G42824,G42825,G42826,G42827,G42828,G42829,G42830,G42831,G42832,G42833,G42834,G42835,G42836,G42837,G42838,G42839,G42840,
       G42841,G42842,G42843,G42844,G42845,G42846,G42847,G42848,G42849,G42850,G42851,G42852,G42853,G42854,G42855,G42856,G42857,G42858,G42859,G42860,
       G42861,G42862,G42863,G42864,G42865,G42866,G42867,G42868,G42869,G42870,G42871,G42872,G42873,G42874,G42875,G42876,G42877,G42878,G42879,G42880,
       G42881,G42882,G42883,G42884,G42885,G42886,G42887,G42888,G42889,G42890,G42891,G42892,G42893,G42894,G42895,G42896,G42897,G42898,G42899,G42900,
       G42901,G42902,G42903,G42904,G42905,G42906,G42907,G42908,G42909,G42910,G42911,G42912,G42913,G42914,G42915,G42916,G42917,G42918,G42919,G42920,
       G42921,G42922,G42923,G42924,G42925,G42926,G42927,G42928,G42929,G42930,G42931,G42932,G42933,G42934,G42935,G42936,G42937,G42938,G42939,G42940,
       G42941,G42942,G42943,G42944,G42945,G42946,G42947,G42948,G42949,G42950,G42951,G42952,G42953,G42954,G42955,G42956,G42957,G42958,G42959,G42960,
       G42961,G42962,G42963,G42964,G42965,G42966,G42967,G42968,G42969,G42970,G42971,G42972,G42973,G42974,G42975,G42976,G42977,G42978,G42979,G42980,
       G42981,G42982,G42983,G42984,G42985,G42986,G42987,G42988,G42989,G42990,G42991,G42992,G42993,G42994,G42995,G42996,G42997,G42998,G42999,G43000,
       G43001,G43002,G43003,G43004,G43005,G43006,G43007,G43008,G43009,G43010,G43011,G43012,G43013,G43014,G43015,G43016,G43017,G43018,G43019,G43020,
       G43021,G43022,G43023,G43024,G43025,G43026,G43027,G43028,G43029,G43030,G43031,G43032,G43033,G43034,G43035,G43036,G43037,G43038,G43039,G43040,
       G43041,G43042,G43043,G43044,G43045,G43046,G43047,G43048,G43049,G43050,G43051,G43052,G43053,G43054,G43055,G43056,G43057,G43058,G43059,G43060,
       G43061,G43062,G43063,G43064,G43065,G43066,G43067,G43068,G43069,G43070,G43071,G43072,G43073,G43074,G43075,G43076,G43077,G43078,G43079,G43080,
       G43081,G43082,G43083,G43084,G43085,G43086,G43087,G43088,G43089,G43090,G43091,G43092,G43093,G43094,G43095,G43096,G43097,G43098,G43099,G43100,
       G43101,G43102,G43103,G43104,G43105,G43106,G43107,G43108,G43109,G43110,G43111,G43112,G43113,G43114,G43115,G43116,G43117,G43118,G43119,G43120,
       G43121,G43122,G43123,G43124,G43125,G43126,G43127,G43128,G43129,G43130,G43131,G43132,G43133,G43134,G43135,G43136,G43137,G43138,G43139,G43140,
       G43141,G43142,G43143,G43144,G43145,G43146,G43147,G43148,G43149,G43150,G43151,G43152,G43153,G43154,G43155,G43156,G43157,G43158,G43159,G43160,
       G43161,G43162,G43163,G43164,G43165,G43166,G43167,G43168,G43169,G43170,G43171,G43172,G43173,G43174,G43175,G43176,G43177,G43178,G43179,G43180,
       G43181,G43182,G43183,G43184,G43185,G43186,G43187,G43188,G43189,G43190,G43191,G43192,G43193,G43194,G43195,G43196,G43197,G43198,G43199,G43200,
       G43201,G43202,G43203,G43204,G43205,G43206,G43207,G43208,G43209,G43210,G43211,G43212,G43213,G43214,G43215,G43216,G43217,G43218,G43219,G43220,
       G43221,G43222,G43223,G43224,G43225,G43226,G43227,G43228,G43229,G43230,G43231,G43232,G43233,G43234,G43235,G43236,G43237,G43238,G43239,G43240,
       G43241,G43242,G43243,G43244,G43245,G43246,G43247,G43248,G43249,G43250,G43251,G43252,G43253,G43254,G43255,G43256,G43257,G43258,G43259,G43260,
       G43261,G43262,G43263,G43264,G43265,G43266,G43267,G43268,G43269,G43270,G43271,G43272,G43273,G43274,G43275,G43276,G43277,G43278,G43279,G43280,
       G43281,G43282,G43283,G43284,G43285,G43286,G43287,G43288,G43289,G43290,G43291,G43292,G43293,G43294,G43295,G43296,G43297,G43298,G43299,G43300,
       G43301,G43302,G43303,G43304,G43305,G43306,G43307,G43308,G43309,G43310,G43311,G43312,G43313,G43314,G43315,G43316,G43317,G43318,G43319,G43320,
       G43321,G43322,G43323,G43324,G43325,G43326,G43327,G43328,G43329,G43330,G43331,G43332,G43333,G43334,G43335,G43336,G43337,G43338,G43339,G43340,
       G43341,G43342,G43343,G43344,G43345,G43346,G43347,G43348,G43349,G43350,G43351,G43352,G43353,G43354,G43355,G43356,G43357,G43358,G43359,G43360,
       G43361,G43362,G43363,G43364,G43365,G43366,G43367,G43368,G43369,G43370,G43371,G43372,G43373,G43374,G43375,G43376,G43377,G43378,G43379,G43380,
       G43381,G43382,G43383,G43384,G43385,G43386,G43387,G43388,G43389,G43390,G43391,G43392,G43393,G43394,G43395,G43396,G43397,G43398,G43399,G43400,
       G43401,G43402,G43403,G43404,G43405,G43406,G43407,G43408,G43409,G43410,G43411,G43412,G43413,G43414,G43415,G43416,G43417,G43418,G43419,G43420,
       G43421,G43422,G43423,G43424,G43425,G43426,G43427,G43428,G43429,G43430,G43431,G43432,G43433,G43434,G43435,G43436,G43437,G43438,G43439,G43440,
       G43441,G43442,G43443,G43444,G43445,G43446,G43447,G43448,G43449,G43450,G43451,G43452,G43453,G43454,G43455,G43456,G43457,G43458,G43459,G43460,
       G43461,G43462,G43463,G43464,G43465,G43466,G43467,G43468,G43469,G43470,G43471,G43472,G43473,G43474,G43475,G43476,G43477,G43478,G43479,G43480,
       G43481,G43482,G43483,G43484,G43485,G43486,G43487,G43488,G43489,G43490,G43491,G43492,G43493,G43494,G43495,G43496,G43497,G43498,G43499,G43500,
       G43501,G43502,G43503,G43504,G43505,G43506,G43507,G43508,G43509,G43510,G43511,G43512,G43513,G43514,G43515,G43516,G43517,G43518,G43519,G43520,
       G43521,G43522,G43523,G43524,G43525,G43526,G43527,G43528,G43529,G43530,G43531,G43532,G43533,G43534,G43535,G43536,G43537,G43538,G43539,G43540,
       G43541,G43542,G43543,G43544,G43545,G43546,G43547,G43548,G43549,G43550,G43551,G43552,G43553,G43554,G43555,G43556,G43557,G43558,G43559,G43560,
       G43561,G43562,G43563,G43564,G43565,G43566,G43567,G43568,G43569,G43570,G43571,G43572,G43573,G43574,G43575,G43576,G43577,G43578,G43579,G43580,
       G43581,G43582,G43583,G43584,G43585,G43586,G43587,G43588,G43589,G43590,G43591,G43592,G43593,G43594,G43595,G43596,G43597,G43598,G43599,G43600,
       G43601,G43602,G43603,G43604,G43605,G43606,G43607,G43608,G43609,G43610,G43611,G43612,G43613,G43614,G43615,G43616,G43617,G43618,G43619,G43620,
       G43621,G43622,G43623,G43624,G43625,G43626,G43627,G43628,G43629,G43630,G43631,G43632,G43633,G43634,G43635,G43636,G43637,G43638,G43639,G43640,
       G43641,G43642,G43643,G43644,G43645,G43646,G43647,G43648,G43649,G43650,G43651,G43652,G43653,G43654,G43655,G43656,G43657,G43658,G43659,G43660,
       G43661,G43662,G43663,G43664,G43665,G43666,G43667,G43668,G43669,G43670,G43671,G43672,G43673,G43674,G43675,G43676,G43677,G43678,G43679,G43680,
       G43681,G43682,G43683,G43684,G43685,G43686,G43687,G43688,G43689,G43690,G43691,G43692,G43693,G43694,G43695,G43696,G43697,G43698,G43699,G43700,
       G43701,G43702,G43703,G43704,G43705,G43706,G43707,G43708,G43709,G43710,G43711,G43712,G43713,G43714,G43715,G43716,G43717,G43718,G43719,G43720,
       G43721,G43722,G43723,G43724,G43725,G43726,G43727,G43728,G43729,G43730,G43731,G43732,G43733,G43734,G43735,G43736,G43737,G43738,G43739,G43740,
       G43741,G43742,G43743,G43744,G43745,G43746,G43747,G43748,G43749,G43750,G43751,G43752,G43753,G43754,G43755,G43756,G43757,G43758,G43759,G43760,
       G43761,G43762,G43763,G43764,G43765,G43766,G43767,G43768,G43769,G43770,G43771,G43772,G43773,G43774,G43775,G43776,G43777,G43778,G43779,G43780,
       G43781,G43782,G43783,G43784,G43785,G43786,G43787,G43788,G43789,G43790,G43791,G43792,G43793,G43794,G43795,G43796,G43797,G43798,G43799,G43800,
       G43801,G43802,G43803,G43804,G43805,G43806,G43807,G43808,G43809,G43810,G43811,G43812,G43813,G43814,G43815,G43816,G43817,G43818,G43819,G43820,
       G43821,G43822,G43823,G43824,G43825,G43826,G43827,G43828,G43829,G43830,G43831,G43832,G43833,G43834,G43835,G43836,G43837,G43838,G43839,G43840,
       G43841,G43842,G43843,G43844,G43845,G43846,G43847,G43848,G43849,G43850,G43851,G43852,G43853,G43854,G43855,G43856,G43857,G43858,G43859,G43860,
       G43861,G43862,G43863,G43864,G43865,G43866,G43867,G43868,G43869,G43870,G43871,G43872,G43873,G43874,G43875,G43876,G43877,G43878,G43879,G43880,
       G43881,G43882,G43883,G43884,G43885,G43886,G43887,G43888,G43889,G43890,G43891,G43892,G43893,G43894,G43895,G43896,G43897,G43898,G43899,G43900,
       G43901,G43902,G43903,G43904,G43905,G43906,G43907,G43908,G43909,G43910,G43911,G43912,G43913,G43914,G43915,G43916,G43917,G43918,G43919,G43920,
       G43921,G43922,G43923,G43924,G43925,G43926,G43927,G43928,G43929,G43930,G43931,G43932,G43933,G43934,G43935,G43936,G43937,G43938,G43939,G43940,
       G43941,G43942,G43943,G43944,G43945,G43946,G43947,G43948,G43949,G43950,G43951,G43952,G43953,G43954,G43955,G43956,G43957,G43958,G43959,G43960,
       G43961,G43962,G43963,G43964,G43965,G43966,G43967,G43968,G43969,G43970,G43971,G43972,G43973,G43974,G43975,G43976,G43977,G43978,G43979,G43980,
       G43981,G43982,G43983,G43984,G43985,G43986,G43987,G43988,G43989,G43990,G43991,G43992,G43993,G43994,G43995,G43996,G43997,G43998,G43999,G44000,
       G44001,G44002,G44003,G44004,G44005,G44006,G44007,G44008,G44009,G44010,G44011,G44012,G44013,G44014,G44015,G44016,G44017,G44018,G44019,G44020,
       G44021,G44022,G44023,G44024,G44025,G44026,G44027,G44028,G44029,G44030,G44031,G44032,G44033,G44034,G44035,G44036,G44037,G44038,G44039,G44040,
       G44041,G44042,G44043,G44044,G44045,G44046,G44047,G44048,G44049,G44050,G44051,G44052,G44053,G44054,G44055,G44056,G44057,G44058,G44059,G44060,
       G44061,G44062,G44063,G44064,G44065,G44066,G44067,G44068,G44069,G44070,G44071,G44072,G44073,G44074,G44075,G44076,G44077,G44078,G44079,G44080,
       G44081,G44082,G44083,G44084,G44085,G44086,G44087,G44088,G44089,G44090,G44091,G44092,G44093,G44094,G44095,G44096,G44097,G44098,G44099,G44100,
       G44101,G44102,G44103,G44104,G44105,G44106,G44107,G44108,G44109,G44110,G44111,G44112,G44113,G44114,G44115,G44116,G44117,G44118,G44119,G44120,
       G44121,G44122,G44123,G44124,G44125,G44126,G44127,G44128,G44129,G44130,G44131,G44132,G44133,G44134,G44135,G44136,G44137,G44138,G44139,G44140,
       G44141,G44142,G44143,G44144,G44145,G44146,G44147,G44148,G44149,G44150,G44151,G44152,G44153,G44154,G44155,G44156,G44157,G44158,G44159,G44160,
       G44161,G44162,G44163,G44164,G44165,G44166,G44167,G44168,G44169,G44170,G44171,G44172,G44173,G44174,G44175,G44176,G44177,G44178,G44179,G44180,
       G44181,G44182,G44183,G44184,G44185,G44186,G44187,G44188,G44189,G44190,G44191,G44192,G44193,G44194,G44195,G44196,G44197,G44198,G44199,G44200,
       G44201,G44202,G44203,G44204,G44205,G44206,G44207,G44208,G44209,G44210,G44211,G44212,G44213,G44214,G44215,G44216,G44217,G44218,G44219,G44220,
       G44221,G44222,G44223,G44224,G44225,G44226,G44227,G44228,G44229,G44230,G44231,G44232,G44233,G44234,G44235,G44236,G44237,G44238,G44239,G44240,
       G44241,G44242,G44243,G44244,G44245,G44246,G44247,G44248,G44249,G44250,G44251,G44252,G44253,G44254,G44255,G44256,G44257,G44258,G44259,G44260,
       G44261,G44262,G44263,G44264,G44265,G44266,G44267,G44268,G44269,G44270,G44271,G44272,G44273,G44274,G44275,G44276,G44277,G44278,G44279,G44280,
       G44281,G44282,G44283,G44284,G44285,G44286,G44287,G44288,G44289,G44290,G44291,G44292,G44293,G44294,G44295,G44296,G44297,G44298,G44299,G44300,
       G44301,G44302,G44303,G44304,G44305,G44306,G44307,G44308,G44309,G44310,G44311,G44312,G44313,G44314,G44315,G44316,G44317,G44318,G44319,G44320,
       G44321,G44322,G44323,G44324,G44325,G44326,G44327,G44328,G44329,G44330,G44331,G44332,G44333,G44334,G44335,G44336,G44337,G44338,G44339,G44340,
       G44341,G44342,G44343,G44344,G44345,G44346,G44347,G44348,G44349,G44350,G44351,G44352,G44353,G44354,G44355,G44356,G44357,G44358,G44359,G44360,
       G44361,G44362,G44363,G44364,G44365,G44366,G44367,G44368,G44369,G44370,G44371,G44372,G44373,G44374,G44375,G44376,G44377,G44378,G44379,G44380,
       G44381,G44382,G44383,G44384,G44385,G44386,G44387,G44388,G44389,G44390,G44391,G44392,G44393,G44394,G44395,G44396,G44397,G44398,G44399,G44400,
       G44401,G44402,G44403,G44404,G44405,G44406,G44407,G44408,G44409,G44410,G44411,G44412,G44413,G44414,G44415,G44416,G44417,G44418,G44419,G44420,
       G44421,G44422,G44423,G44424,G44425,G44426,G44427,G44428,G44429,G44430,G44431,G44432,G44433,G44434,G44435,G44436,G44437,G44438,G44439,G44440,
       G44441,G44442,G44443,G44444,G44445,G44446,G44447,G44448,G44449,G44450,G44451,G44452,G44453,G44454,G44455,G44456,G44457,G44458,G44459,G44460,
       G44461,G44462,G44463,G44464,G44465,G44466,G44467,G44468,G44469,G44470,G44471,G44472,G44473,G44474,G44475,G44476,G44477,G44478,G44479,G44480,
       G44481,G44482,G44483,G44484,G44485,G44486,G44487,G44488,G44489,G44490,G44491,G44492,G44493,G44494,G44495,G44496,G44497,G44498,G44499,G44500,
       G44501,G44502,G44503,G44504,G44505,G44506,G44507,G44508,G44509,G44510,G44511,G44512,G44513,G44514,G44515,G44516,G44517,G44518,G44519,G44520,
       G44521,G44522,G44523,G44524,G44525,G44526,G44527,G44528,G44529,G44530,G44531,G44532,G44533,G44534,G44535,G44536,G44537,G44538,G44539,G44540,
       G44541,G44542,G44543,G44544,G44545,G44546,G44547,G44548,G44549,G44550,G44551,G44552,G44553,G44554,G44555,G44556,G44557,G44558,G44559,G44560,
       G44561,G44562,G44563,G44564,G44565,G44566,G44567,G44568,G44569,G44570,G44571,G44572,G44573,G44574,G44575,G44576,G44577,G44578,G44579,G44580,
       G44581,G44582,G44583,G44584,G44585,G44586,G44587,G44588,G44589,G44590,G44591,G44592,G44593,G44594,G44595,G44596,G44597,G44598,G44599,G44600,
       G44601,G44602,G44603,G44604,G44605,G44606,G44607,G44608,G44609,G44610,G44611,G44612,G44613,G44614,G44615,G44616,G44617,G44618,G44619,G44620,
       G44621,G44622,G44623,G44624,G44625,G44626,G44627,G44628,G44629,G44630,G44631,G44632,G44633,G44634,G44635,G44636,G44637,G44638,G44639,G44640,
       G44641,G44642,G44643,G44644,G44645,G44646,G44647,G44648,G44649,G44650,G44651,G44652,G44653,G44654,G44655,G44656,G44657,G44658,G44659,G44660,
       G44661,G44662,G44663,G44664,G44665,G44666,G44667,G44668,G44669,G44670,G44671,G44672,G44673,G44674,G44675,G44676,G44677,G44678,G44679,G44680,
       G44681,G44682,G44683,G44684,G44685,G44686,G44687,G44688,G44689,G44690,G44691,G44692,G44693,G44694,G44695,G44696,G44697,G44698,G44699,G44700,
       G44701,G44702,G44703,G44704,G44705,G44706,G44707,G44708,G44709,G44710,G44711,G44712,G44713,G44714,G44715,G44716,G44717,G44718,G44719,G44720,
       G44721,G44722,G44723,G44724,G44725,G44726,G44727,G44728,G44729,G44730,G44731,G44732,G44733,G44734,G44735,G44736,G44737,G44738,G44739,G44740,
       G44741,G44742,G44743,G44744,G44745,G44746,G44747,G44748,G44749,G44750,G44751,G44752,G44753,G44754,G44755,G44756,G44757,G44758,G44759,G44760,
       G44761,G44762,G44763,G44764,G44765,G44766,G44767,G44768,G44769,G44770,G44771,G44772,G44773,G44774,G44775,G44776,G44777,G44778,G44779,G44780,
       G44781,G44782,G44783,G44784,G44785,G44786,G44787,G44788,G44789,G44790,G44791,G44792,G44793,G44794,G44795,G44796,G44797,G44798,G44799,G44800,
       G44801,G44802,G44803,G44804,G44805,G44806,G44807,G44808,G44809,G44810,G44811,G44812,G44813,G44814,G44815,G44816,G44817,G44818,G44819,G44820,
       G44821,G44822,G44823,G44824,G44825,G44826,G44827,G44828,G44829,G44830,G44831,G44832,G44833,G44834,G44835,G44836,G44837,G44838,G44839,G44840,
       G44841,G44842,G44843,G44844,G44845,G44846,G44847,G44848,G44849,G44850,G44851,G44852,G44853,G44854,G44855,G44856,G44857,G44858,G44859,G44860,
       G44861,G44862,G44863,G44864,G44865,G44866,G44867,G44868,G44869,G44870,G44871,G44872,G44873,G44874,G44875,G44876,G44877,G44878,G44879,G44880,
       G44881,G44882,G44883,G44884,G44885,G44886,G44887,G44888,G44889,G44890,G44891,G44892,G44893,G44894,G44895,G44896,G44897,G44898,G44899,G44900,
       G44901,G44902,G44903,G44904,G44905,G44906,G44907,G44908,G44909,G44910,G44911,G44912,G44913,G44914,G44915,G44916,G44917,G44918,G44919,G44920,
       G44921,G44922,G44923,G44924,G44925,G44926,G44927,G44928,G44929,G44930,G44931,G44932,G44933,G44934,G44935,G44936,G44937,G44938,G44939,G44940,
       G44941,G44942,G44943,G44944,G44945,G44946,G44947,G44948,G44949,G44950,G44951,G44952,G44953,G44954,G44955,G44956,G44957,G44958,G44959,G44960,
       G44961,G44962,G44963,G44964,G44965,G44966,G44967,G44968,G44969,G44970,G44971,G44972,G44973,G44974,G44975,G44976,G44977,G44978,G44979,G44980,
       G44981,G44982,G44983,G44984,G44985,G44986,G44987,G44988,G44989,G44990,G44991,G44992,G44993,G44994,G44995,G44996,G44997,G44998,G44999,G45000,
       G45001,G45002,G45003,G45004,G45005,G45006,G45007,G45008,G45009,G45010,G45011,G45012,G45013,G45014,G45015,G45016,G45017,G45018,G45019,G45020,
       G45021,G45022,G45023,G45024,G45025,G45026,G45027,G45028,G45029,G45030,G45031,G45032,G45033,G45034,G45035,G45036,G45037,G45038,G45039,G45040,
       G45041,G45042,G45043,G45044,G45045,G45046,G45047,G45048,G45049,G45050,G45051,G45052,G45053,G45054,G45055,G45056,G45057,G45058,G45059,G45060,
       G45061,G45062,G45063,G45064,G45065,G45066,G45067,G45068,G45069,G45070,G45071,G45072,G45073,G45074,G45075,G45076,G45077,G45078,G45079,G45080,
       G45081,G45082,G45083,G45084,G45085,G45086,G45087,G45088,G45089,G45090,G45091,G45092,G45093,G45094,G45095,G45096,G45097,G45098,G45099,G45100,
       G45101,G45102,G45103,G45104,G45105,G45106,G45107,G45108,G45109,G45110,G45111,G45112,G45113,G45114,G45115,G45116,G45117,G45118,G45119,G45120,
       G45121,G45122,G45123,G45124,G45125,G45126,G45127,G45128,G45129,G45130,G45131,G45132,G45133,G45134,G45135,G45136,G45137,G45138,G45139,G45140,
       G45141,G45142,G45143,G45144,G45145,G45146,G45147,G45148,G45149,G45150,G45151,G45152,G45153,G45154,G45155,G45156,G45157,G45158,G45159,G45160,
       G45161,G45162,G45163,G45164,G45165,G45166,G45167,G45168,G45169,G45170,G45171,G45172,G45173,G45174,G45175,G45176,G45177,G45178,G45179,G45180,
       G45181,G45182,G45183,G45184,G45185,G45186,G45187,G45188,G45189,G45190,G45191,G45192,G45193,G45194,G45195,G45196,G45197,G45198,G45199,G45200,
       G45201,G45202,G45203,G45204,G45205,G45206,G45207,G45208,G45209,G45210,G45211,G45212,G45213,G45214,G45215,G45216,G45217,G45218,G45219,G45220,
       G45221,G45222,G45223,G45224,G45225,G45226,G45227,G45228,G45229,G45230,G45231,G45232,G45233,G45234,G45235,G45236,G45237,G45238,G45239,G45240,
       G45241,G45242,G45243,G45244,G45245,G45246,G45247,G45248,G45249,G45250,G45251,G45252,G45253,G45254,G45255,G45256,G45257,G45258,G45259,G45260,
       G45261,G45262,G45263,G45264,G45265,G45266,G45267,G45268,G45269,G45270,G45271,G45272,G45273,G45274,G45275,G45276,G45277,G45278,G45279,G45280,
       G45281,G45282,G45283,G45284,G45285,G45286,G45287,G45288,G45289,G45290,G45291,G45292,G45293,G45294,G45295,G45296,G45297,G45298,G45299,G45300,
       G45301,G45302,G45303,G45304,G45305,G45306,G45307,G45308,G45309,G45310,G45311,G45312,G45313,G45314,G45315,G45316,G45317,G45318,G45319,G45320,
       G45321,G45322,G45323,G45324,G45325,G45326,G45327,G45328,G45329,G45330,G45331,G45332,G45333,G45334,G45335,G45336,G45337,G45338,G45339,G45340,
       G45341,G45342,G45343,G45344,G45345,G45346,G45347,G45348,G45349,G45350,G45351,G45352,G45353,G45354,G45355,G45356,G45357,G45358,G45359,G45360,
       G45361,G45362,G45363,G45364,G45365,G45366,G45367,G45368,G45369,G45370,G45371,G45372,G45373,G45374,G45375,G45376,G45377,G45378,G45379,G45380,
       G45381,G45382,G45383,G45384,G45385,G45386,G45387,G45388,G45389,G45390,G45391,G45392,G45393,G45394,G45395,G45396,G45397,G45398,G45399,G45400,
       G45401,G45402,G45403,G45404,G45405,G45406,G45407,G45408,G45409,G45410,G45411,G45412,G45413,G45414,G45415,G45416,G45417,G45418,G45419,G45420,
       G45421,G45422,G45423,G45424,G45425,G45426,G45427,G45428,G45429,G45430,G45431,G45432,G45433,G45434,G45435,G45436,G45437,G45438,G45439,G45440,
       G45441,G45442,G45443,G45444,G45445,G45446,G45447,G45448,G45449,G45450,G45451,G45452,G45453,G45454,G45455,G45456,G45457,G45458,G45459,G45460,
       G45461,G45462,G45463,G45464,G45465,G45466,G45467,G45468,G45469,G45470,G45471,G45472,G45473,G45474,G45475,G45476,G45477,G45478,G45479,G45480,
       G45481,G45482,G45483,G45484,G45485,G45486,G45487,G45488,G45489,G45490,G45491,G45492,G45493,G45494,G45495,G45496,G45497,G45498,G45499,G45500,
       G45501,G45502,G45503,G45504,G45505,G45506,G45507,G45508,G45509,G45510,G45511,G45512,G45513,G45514,G45515,G45516,G45517,G45518,G45519,G45520,
       G45521,G45522,G45523,G45524,G45525,G45526,G45527,G45528,G45529,G45530,G45531,G45532,G45533,G45534,G45535,G45536,G45537,G45538,G45539,G45540,
       G45541,G45542,G45543,G45544,G45545,G45546,G45547,G45548,G45549,G45550,G45551,G45552,G45553,G45554,G45555,G45556,G45557,G45558,G45559,G45560,
       G45561,G45562,G45563,G45564,G45565,G45566,G45567,G45568,G45569,G45570,G45571,G45572,G45573,G45574,G45575,G45576,G45577,G45578,G45579,G45580,
       G45581,G45582,G45583,G45584,G45585,G45586,G45587,G45588,G45589,G45590,G45591,G45592,G45593,G45594,G45595,G45596,G45597,G45598,G45599,G45600,
       G45601,G45602,G45603,G45604,G45605,G45606,G45607,G45608,G45609,G45610,G45611,G45612,G45613,G45614,G45615,G45616,G45617,G45618,G45619,G45620,
       G45621,G45622,G45623,G45624,G45625,G45626,G45627,G45628,G45629,G45630,G45631,G45632,G45633,G45634,G45635,G45636,G45637,G45638,G45639,G45640,
       G45641,G45642,G45643,G45644,G45645,G45646,G45647,G45648,G45649,G45650,G45651,G45652,G45653,G45654,G45655,G45656,G45657,G45658,G45659,G45660,
       G45661,G45662,G45663,G45664,G45665,G45666,G45667,G45668,G45669,G45670,G45671,G45672,G45673,G45674,G45675,G45676,G45677,G45678,G45679,G45680,
       G45681,G45682,G45683,G45684,G45685,G45686,G45687,G45688,G45689,G45690,G45691,G45692,G45693,G45694,G45695,G45696,G45697,G45698,G45699,G45700,
       G45701,G45702,G45703,G45704,G45705,G45706,G45707,G45708,G45709,G45710,G45711,G45712,G45713,G45714,G45715,G45716,G45717,G45718,G45719,G45720,
       G45721,G45722,G45723,G45724,G45725,G45726,G45727,G45728,G45729,G45730,G45731,G45732,G45733,G45734,G45735,G45736,G45737,G45738,G45739,G45740,
       G45741,G45742,G45743,G45744,G45745,G45746,G45747,G45748,G45749,G45750,G45751,G45752,G45753,G45754,G45755,G45756,G45757,G45758,G45759,G45760,
       G45761,G45762,G45763,G45764,G45765,G45766,G45767,G45768,G45769,G45770,G45771,G45772,G45773,G45774,G45775,G45776,G45777,G45778,G45779,G45780,
       G45781,G45782,G45783,G45784,G45785,G45786,G45787,G45788,G45789,G45790,G45791,G45792,G45793,G45794,G45795,G45796,G45797,G45798,G45799,G45800,
       G45801,G45802,G45803,G45804,G45805,G45806,G45807,G45808,G45809,G45810,G45811,G45812,G45813,G45814,G45815,G45816,G45817,G45818,G45819,G45820,
       G45821,G45822,G45823,G45824,G45825,G45826,G45827,G45828,G45829,G45830,G45831,G45832,G45833,G45834,G45835,G45836,G45837,G45838,G45839,G45840,
       G45841,G45842,G45843,G45844,G45845,G45846,G45847,G45848,G45849,G45850,G45851,G45852,G45853,G45854,G45855,G45856,G45857,G45858,G45859,G45860,
       G45861,G45862,G45863,G45864,G45865,G45866,G45867,G45868,G45869,G45870,G45871,G45872,G45873,G45874,G45875,G45876,G45877,G45878,G45879,G45880,
       G45881,G45882,G45883,G45884,G45885,G45886,G45887,G45888,G45889,G45890,G45891,G45892,G45893,G45894,G45895,G45896,G45897,G45898,G45899,G45900,
       G45901,G45902,G45903,G45904,G45905,G45906,G45907,G45908,G45909,G45910,G45911,G45912,G45913,G45914,G45915,G45916,G45917,G45918,G45919,G45920,
       G45921,G45922,G45923,G45924,G45925,G45926,G45927,G45928,G45929,G45930,G45931,G45932,G45933,G45934,G45935,G45936,G45937,G45938,G45939,G45940,
       G45941,G45942,G45943,G45944,G45945,G45946,G45947,G45948,G45949,G45950,G45951,G45952,G45953,G45954,G45955,G45956,G45957,G45958,G45959,G45960,
       G45961,G45962,G45963,G45964,G45965,G45966,G45967,G45968,G45969,G45970,G45971,G45972,G45973,G45974,G45975,G45976,G45977,G45978,G45979,G45980,
       G45981,G45982,G45983,G45984,G45985,G45986,G45987,G45988,G45989,G45990,G45991,G45992,G45993,G45994,G45995,G45996,G45997,G45998,G45999,G46000,
       G46001,G46002,G46003,G46004,G46005,G46006,G46007,G46008,G46009,G46010,G46011,G46012,G46013,G46014,G46015,G46016,G46017,G46018,G46019,G46020,
       G46021,G46022,G46023,G46024,G46025,G46026,G46027,G46028,G46029,G46030,G46031,G46032,G46033,G46034,G46035,G46036,G46037,G46038,G46039,G46040,
       G46041,G46042,G46043,G46044,G46045,G46046,G46047,G46048,G46049,G46050,G46051,G46052,G46053,G46054,G46055,G46056,G46057,G46058,G46059,G46060,
       G46061,G46062,G46063,G46064,G46065,G46066,G46067,G46068,G46069,G46070,G46071,G46072,G46073,G46074,G46075,G46076,G46077,G46078,G46079,G46080,
       G46081,G46082,G46083,G46084,G46085,G46086,G46087,G46088,G46089,G46090,G46091,G46092,G46093,G46094,G46095,G46096,G46097,G46098,G46099,G46100,
       G46101,G46102,G46103,G46104,G46105,G46106,G46107,G46108,G46109,G46110,G46111,G46112,G46113,G46114,G46115,G46116,G46117,G46118,G46119,G46120,
       G46121,G46122,G46123,G46124,G46125,G46126,G46127,G46128,G46129,G46130,G46131,G46132,G46133,G46134,G46135,G46136,G46137,G46138,G46139,G46140,
       G46141,G46142,G46143,G46144,G46145,G46146,G46147,G46148,G46149,G46150,G46151,G46152,G46153,G46154,G46155,G46156,G46157,G46158,G46159,G46160,
       G46161,G46162,G46163,G46164,G46165,G46166,G46167,G46168,G46169,G46170,G46171,G46172,G46173,G46174,G46175,G46176,G46177,G46178,G46179,G46180,
       G46181,G46182,G46183,G46184,G46185,G46186,G46187,G46188,G46189,G46190,G46191,G46192,G46193,G46194,G46195,G46196,G46197,G46198,G46199,G46200,
       G46201,G46202,G46203,G46204,G46205,G46206,G46207,G46208,G46209,G46210,G46211,G46212,G46213,G46214,G46215,G46216,G46217,G46218,G46219,G46220,
       G46221,G46222,G46223,G46224,G46225,G46226,G46227,G46228,G46229,G46230,G46231,G46232,G46233,G46234,G46235,G46236,G46237,G46238,G46239,G46240,
       G46241,G46242,G46243,G46244,G46245,G46246,G46247,G46248,G46249,G46250,G46251,G46252,G46253,G46254,G46255,G46256,G46257,G46258,G46259,G46260,
       G46261,G46262,G46263,G46264,G46265,G46266,G46267,G46268,G46269,G46270,G46271,G46272,G46273,G46274,G46275,G46276,G46277,G46278,G46279,G46280,
       G46281,G46282,G46283,G46284,G46285,G46286,G46287,G46288,G46289,G46290,G46291,G46292,G46293,G46294,G46295,G46296,G46297,G46298,G46299,G46300,
       G46301,G46302,G46303,G46304,G46305,G46306,G46307,G46308,G46309,G46310,G46311,G46312,G46313,G46314,G46315,G46316,G46317,G46318,G46319,G46320,
       G46321,G46322,G46323,G46324,G46325,G46326,G46327,G46328,G46329,G46330,G46331,G46332,G46333,G46334,G46335,G46336,G46337,G46338,G46339,G46340,
       G46341,G46342,G46343,G46344,G46345,G46346,G46347,G46348,G46349,G46350,G46351,G46352,G46353,G46354,G46355,G46356,G46357,G46358,G46359,G46360,
       G46361,G46362,G46363,G46364,G46365,G46366,G46367,G46368,G46369,G46370,G46371,G46372,G46373,G46374,G46375,G46376,G46377,G46378,G46379,G46380,
       G46381,G46382,G46383,G46384,G46385,G46386,G46387,G46388,G46389,G46390,G46391,G46392,G46393,G46394,G46395,G46396,G46397,G46398,G46399,G46400,
       G46401,G46402,G46403,G46404,G46405,G46406,G46407,G46408,G46409,G46410,G46411,G46412,G46413,G46414,G46415,G46416,G46417,G46418,G46419,G46420,
       G46421,G46422,G46423,G46424,G46425,G46426,G46427,G46428,G46429,G46430,G46431,G46432,G46433,G46434,G46435,G46436,G46437,G46438,G46439,G46440,
       G46441,G46442,G46443,G46444,G46445,G46446,G46447,G46448,G46449,G46450,G46451,G46452,G46453,G46454,G46455,G46456,G46457,G46458,G46459,G46460,
       G46461,G46462,G46463,G46464,G46465,G46466,G46467,G46468,G46469,G46470,G46471,G46472,G46473,G46474,G46475,G46476,G46477,G46478,G46479,G46480,
       G46481,G46482,G46483,G46484,G46485,G46486,G46487,G46488,G46489,G46490,G46491,G46492,G46493,G46494,G46495,G46496,G46497,G46498,G46499,G46500,
       G46501,G46502,G46503,G46504,G46505,G46506,G46507,G46508,G46509,G46510,G46511,G46512,G46513,G46514,G46515,G46516,G46517,G46518,G46519,G46520,
       G46521,G46522,G46523,G46524,G46525,G46526,G46527,G46528,G46529,G46530,G46531,G46532,G46533,G46534,G46535,G46536,G46537,G46538,G46539,G46540,
       G46541,G46542,G46543,G46544,G46545,G46546,G46547,G46548,G46549,G46550,G46551,G46552,G46553,G46554,G46555,G46556,G46557,G46558,G46559,G46560,
       G46561,G46562,G46563,G46564,G46565,G46566,G46567,G46568,G46569,G46570,G46571,G46572,G46573,G46574,G46575,G46576,G46577,G46578,G46579,G46580,
       G46581,G46582,G46583,G46584,G46585,G46586,G46587,G46588,G46589,G46590,G46591,G46592,G46593,G46594,G46595,G46596,G46597,G46598,G46599,G46600,
       G46601,G46602,G46603,G46604,G46605,G46606,G46607,G46608,G46609,G46610,G46611,G46612,G46613,G46614,G46615,G46616,G46617,G46618,G46619,G46620,
       G46621,G46622,G46623,G46624,G46625,G46626,G46627,G46628,G46629,G46630,G46631,G46632,G46633,G46634,G46635,G46636,G46637,G46638,G46639,G46640,
       G46641,G46642,G46643,G46644,G46645,G46646,G46647,G46648,G46649,G46650,G46651,G46652,G46653,G46654,G46655,G46656,G46657,G46658,G46659,G46660,
       G46661,G46662,G46663,G46664,G46665,G46666,G46667,G46668,G46669,G46670,G46671,G46672,G46673,G46674,G46675,G46676,G46677,G46678,G46679,G46680,
       G46681,G46682,G46683,G46684,G46685,G46686,G46687,G46688,G46689,G46690,G46691,G46692,G46693,G46694,G46695,G46696,G46697,G46698,G46699,G46700,
       G46701,G46702,G46703,G46704,G46705,G46706,G46707,G46708,G46709,G46710,G46711,G46712,G46713,G46714,G46715,G46716,G46717,G46718,G46719,G46720,
       G46721,G46722,G46723,G46724,G46725,G46726,G46727,G46728,G46729,G46730,G46731,G46732,G46733,G46734,G46735,G46736,G46737,G46738,G46739,G46740,
       G46741,G46742,G46743,G46744,G46745,G46746,G46747,G46748,G46749,G46750,G46751,G46752,G46753,G46754,G46755,G46756,G46757,G46758,G46759,G46760,
       G46761,G46762,G46763,G46764,G46765,G46766,G46767,G46768,G46769,G46770,G46771,G46772,G46773,G46774,G46775,G46776,G46777,G46778,G46779,G46780,
       G46781,G46782,G46783,G46784,G46785,G46786,G46787,G46788,G46789,G46790,G46791,G46792,G46793,G46794,G46795,G46796,G46797,G46798,G46799,G46800,
       G46801,G46802,G46803,G46804,G46805,G46806,G46807,G46808,G46809,G46810,G46811,G46812,G46813,G46814,G46815,G46816,G46817,G46818,G46819,G46820,
       G46821,G46822,G46823,G46824,G46825,G46826,G46827,G46828,G46829,G46830,G46831,G46832,G46833,G46834,G46835,G46836,G46837,G46838,G46839,G46840,
       G46841,G46842,G46843,G46844,G46845,G46846,G46847,G46848,G46849,G46850,G46851,G46852,G46853,G46854,G46855,G46856,G46857,G46858,G46859,G46860,
       G46861,G46862,G46863,G46864,G46865,G46866,G46867,G46868,G46869,G46870,G46871,G46872,G46873,G46874,G46875,G46876,G46877,G46878,G46879,G46880,
       G46881,G46882,G46883,G46884,G46885,G46886,G46887,G46888,G46889,G46890,G46891,G46892,G46893,G46894,G46895,G46896,G46897,G46898,G46899,G46900,
       G46901,G46902,G46903,G46904,G46905,G46906,G46907,G46908,G46909,G46910,G46911,G46912,G46913,G46914,G46915,G46916,G46917,G46918,G46919,G46920,
       G46921,G46922,G46923,G46924,G46925,G46926,G46927,G46928,G46929,G46930,G46931,G46932,G46933,G46934,G46935,G46936,G46937,G46938,G46939,G46940,
       G46941,G46942,G46943,G46944,G46945,G46946,G46947,G46948,G46949,G46950,G46951,G46952,G46953,G46954,G46955,G46956,G46957,G46958,G46959,G46960,
       G46961,G46962,G46963,G46964,G46965,G46966,G46967,G46968,G46969,G46970,G46971,G46972,G46973,G46974,G46975,G46976,G46977,G46978,G46979,G46980,
       G46981,G46982,G46983,G46984,G46985,G46986,G46987,G46988,G46989,G46990,G46991,G46992,G46993,G46994,G46995,G46996,G46997,G46998,G46999,G47000,
       G47001,G47002,G47003,G47004,G47005,G47006,G47007,G47008,G47009,G47010,G47011,G47012,G47013,G47014,G47015,G47016,G47017,G47018,G47019,G47020,
       G47021,G47022,G47023,G47024,G47025,G47026,G47027,G47028,G47029,G47030,G47031,G47032,G47033,G47034,G47035,G47036,G47037,G47038,G47039,G47040,
       G47041,G47042,G47043,G47044,G47045,G47046,G47047,G47048,G47049,G47050,G47051,G47052,G47053,G47054,G47055,G47056,G47057,G47058,G47059,G47060,
       G47061,G47062,G47063,G47064,G47065,G47066,G47067,G47068,G47069,G47070,G47071,G47072,G47073,G47074,G47075,G47076,G47077,G47078,G47079,G47080,
       G47081,G47082,G47083,G47084,G47085,G47086,G47087,G47088,G47089,G47090,G47091,G47092,G47093,G47094,G47095,G47096,G47097,G47098,G47099,G47100,
       G47101,G47102,G47103,G47104,G47105,G47106,G47107,G47108,G47109,G47110,G47111,G47112,G47113,G47114,G47115,G47116,G47117,G47118,G47119,G47120,
       G47121,G47122,G47123,G47124,G47125,G47126,G47127,G47128,G47129,G47130,G47131,G47132,G47133,G47134,G47135,G47136,G47137,G47138,G47139,G47140,
       G47141,G47142,G47143,G47144,G47145,G47146,G47147,G47148,G47149,G47150,G47151,G47152,G47153,G47154,G47155,G47156,G47157,G47158,G47159,G47160,
       G47161,G47162,G47163,G47164,G47165,G47166,G47167,G47168,G47169,G47170,G47171,G47172,G47173,G47174,G47175,G47176,G47177,G47178,G47179,G47180,
       G47181,G47182,G47183,G47184,G47185,G47186,G47187,G47188,G47189,G47190,G47191,G47192,G47193,G47194,G47195,G47196,G47197,G47198,G47199,G47200,
       G47201,G47202,G47203,G47204,G47205,G47206,G47207,G47208,G47209,G47210,G47211,G47212,G47213,G47214,G47215,G47216,G47217,G47218,G47219,G47220,
       G47221,G47222,G47223,G47224,G47225,G47226,G47227,G47228,G47229,G47230,G47231,G47232,G47233,G47234,G47235,G47236,G47237,G47238,G47239,G47240,
       G47241,G47242,G47243,G47244,G47245,G47246,G47247,G47248,G47249,G47250,G47251,G47252,G47253,G47254,G47255,G47256,G47257,G47258,G47259,G47260,
       G47261,G47262,G47263,G47264,G47265,G47266,G47267,G47268,G47269,G47270,G47271,G47272,G47273,G47274,G47275,G47276,G47277,G47278,G47279,G47280,
       G47281,G47282,G47283,G47284,G47285,G47286,G47287,G47288,G47289,G47290,G47291,G47292,G47293,G47294,G47295,G47296,G47297,G47298,G47299,G47300,
       G47301,G47302,G47303,G47304,G47305,G47306,G47307,G47308,G47309,G47310,G47311,G47312,G47313,G47314,G47315,G47316,G47317,G47318,G47319,G47320,
       G47321,G47322,G47323,G47324,G47325,G47326,G47327,G47328,G47329,G47330,G47331,G47332,G47333,G47334,G47335,G47336,G47337,G47338,G47339,G47340,
       G47341,G47342,G47343,G47344,G47345,G47346,G47347,G47348,G47349,G47350,G47351,G47352,G47353,G47354,G47355,G47356,G47357,G47358,G47359,G47360,
       G47361,G47362,G47363,G47364,G47365,G47366,G47367,G47368,G47369,G47370,G47371,G47372,G47373,G47374,G47375,G47376,G47377,G47378,G47379,G47380,
       G47381,G47382,G47383,G47384,G47385,G47386,G47387,G47388,G47389,G47390,G47391,G47392,G47393,G47394,G47395,G47396,G47397,G47398,G47399,G47400,
       G47401,G47402,G47403,G47404,G47405,G47406,G47407,G47408,G47409,G47410,G47411,G47412,G47413,G47414,G47415,G47416,G47417,G47418,G47419,G47420,
       G47421,G47422,G47423,G47424,G47425,G47426,G47427,G47428,G47429,G47430,G47431,G47432,G47433,G47434,G47435,G47436,G47437,G47438,G47439,G47440,
       G47441,G47442,G47443,G47444,G47445,G47446,G47447,G47448,G47449,G47450,G47451,G47452,G47453,G47454,G47455,G47456,G47457,G47458,G47459,G47460,
       G47461,G47462,G47463,G47464,G47465,G47466,G47467,G47468,G47469,G47470,G47471,G47472,G47473,G47474,G47475,G47476,G47477,G47478,G47479,G47480,
       G47481,G47482,G47483,G47484,G47485,G47486,G47487,G47488,G47489,G47490,G47491,G47492,G47493,G47494,G47495,G47496,G47497,G47498,G47499,G47500,
       G47501,G47502,G47503,G47504,G47505,G47506,G47507,G47508,G47509,G47510,G47511,G47512,G47513,G47514,G47515,G47516,G47517,G47518,G47519,G47520,
       G47521,G47522,G47523,G47524,G47525,G47526,G47527,G47528,G47529,G47530,G47531,G47532,G47533,G47534,G47535,G47536,G47537,G47538,G47539,G47540,
       G47541,G47542,G47543,G47544,G47545,G47546,G47547,G47548,G47549,G47550,G47551,G47552,G47553,G47554,G47555,G47556,G47557,G47558,G47559,G47560,
       G47561,G47562,G47563,G47564,G47565,G47566,G47567,G47568,G47569,G47570,G47571,G47572,G47573,G47574,G47575,G47576,G47577,G47578,G47579,G47580,
       G47581,G47582,G47583,G47584,G47585,G47586,G47587,G47588,G47589,G47590,G47591,G47592,G47593,G47594,G47595,G47596,G47597,G47598,G47599,G47600,
       G47601,G47602,G47603,G47604,G47605,G47606,G47607,G47608,G47609,G47610,G47611,G47612,G47613,G47614,G47615,G47616,G47617,G47618,G47619,G47620,
       G47621,G47622,G47623,G47624,G47625,G47626,G47627,G47628,G47629,G47630,G47631,G47632,G47633,G47634,G47635,G47636,G47637,G47638,G47639,G47640,
       G47641,G47642,G47643,G47644,G47645,G47646,G47647,G47648,G47649,G47650,G47651,G47652,G47653,G47654,G47655,G47656,G47657,G47658,G47659,G47660,
       G47661,G47662,G47663,G47664,G47665,G47666,G47667,G47668,G47669,G47670,G47671,G47672,G47673,G47674,G47675,G47676,G47677,G47678,G47679,G47680,
       G47681,G47682,G47683,G47684,G47685,G47686,G47687,G47688,G47689,G47690,G47691,G47692,G47693,G47694,G47695,G47696,G47697,G47698,G47699,G47700,
       G47701,G47702,G47703,G47704,G47705,G47706,G47707,G47708,G47709,G47710,G47711,G47712,G47713,G47714,G47715,G47716,G47717,G47718,G47719,G47720,
       G47721,G47722,G47723,G47724,G47725,G47726,G47727,G47728,G47729,G47730,G47731,G47732,G47733,G47734,G47735,G47736,G47737,G47738,G47739,G47740,
       G47741,G47742,G47743,G47744,G47745,G47746,G47747,G47748,G47749,G47750,G47751,G47752,G47753,G47754,G47755,G47756,G47757,G47758,G47759,G47760,
       G47761,G47762,G47763,G47764,G47765,G47766,G47767,G47768,G47769,G47770,G47771,G47772,G47773,G47774,G47775,G47776,G47777,G47778,G47779,G47780,
       G47781,G47782,G47783,G47784,G47785,G47786,G47787,G47788,G47789,G47790,G47791,G47792,G47793,G47794,G47795,G47796,G47797,G47798,G47799,G47800,
       G47801,G47802,G47803,G47804,G47805,G47806,G47807,G47808,G47809,G47810,G47811,G47812,G47813,G47814,G47815,G47816,G47817,G47818,G47819,G47820,
       G47821,G47822,G47823,G47824,G47825,G47826,G47827,G47828,G47829,G47830,G47831,G47832,G47833,G47834,G47835,G47836,G47837,G47838,G47839,G47840,
       G47841,G47842,G47843,G47844,G47845,G47846,G47847,G47848,G47849,G47850,G47851,G47852,G47853,G47854,G47855,G47856,G47857,G47858,G47859,G47860,
       G47861,G47862,G47863,G47864,G47865,G47866,G47867,G47868,G47869,G47870,G47871,G47872,G47873,G47874,G47875,G47876,G47877,G47878,G47879,G47880,
       G47881,G47882,G47883,G47884,G47885,G47886,G47887,G47888,G47889,G47890,G47891,G47892,G47893,G47894,G47895,G47896,G47897,G47898,G47899,G47900,
       G47901,G47902,G47903,G47904,G47905,G47906,G47907,G47908,G47909,G47910,G47911,G47912,G47913,G47914,G47915,G47916,G47917,G47918,G47919,G47920,
       G47921,G47922,G47923,G47924,G47925,G47926,G47927,G47928,G47929,G47930,G47931,G47932,G47933,G47934,G47935,G47936,G47937,G47938,G47939,G47940,
       G47941,G47942,G47943,G47944,G47945,G47946,G47947,G47948,G47949,G47950,G47951,G47952,G47953,G47954,G47955,G47956,G47957,G47958,G47959,G47960,
       G47961,G47962,G47963,G47964,G47965,G47966,G47967,G47968,G47969,G47970,G47971,G47972,G47973,G47974,G47975,G47976,G47977,G47978,G47979,G47980,
       G47981,G47982,G47983,G47984,G47985,G47986,G47987,G47988,G47989,G47990,G47991,G47992,G47993,G47994,G47995,G47996,G47997,G47998,G47999,G48000,
       G48001,G48002,G48003,G48004,G48005,G48006,G48007,G48008,G48009,G48010,G48011,G48012,G48013,G48014,G48015,G48016,G48017,G48018,G48019,G48020,
       G48021,G48022,G48023,G48024,G48025,G48026,G48027,G48028,G48029,G48030,G48031,G48032,G48033,G48034,G48035,G48036,G48037,G48038,G48039,G48040,
       G48041,G48042,G48043,G48044,G48045,G48046,G48047,G48048,G48049,G48050,G48051,G48052,G48053,G48054,G48055,G48056,G48057,G48058,G48059,G48060,
       G48061,G48062,G48063,G48064,G48065,G48066,G48067,G48068,G48069,G48070,G48071,G48072,G48073,G48074,G48075,G48076,G48077,G48078,G48079,G48080,
       G48081,G48082,G48083,G48084,G48085,G48086,G48087,G48088,G48089,G48090,G48091,G48092,G48093,G48094,G48095,G48096,G48097,G48098,G48099,G48100,
       G48101,G48102,G48103,G48104,G48105,G48106,G48107,G48108,G48109,G48110,G48111,G48112,G48113,G48114,G48115,G48116,G48117,G48118,G48119,G48120,
       G48121,G48122,G48123,G48124,G48125,G48126,G48127,G48128,G48129,G48130,G48131,G48132,G48133,G48134,G48135,G48136,G48137,G48138,G48139,G48140,
       G48141,G48142,G48143,G48144,G48145,G48146,G48147,G48148,G48149,G48150,G48151,G48152,G48153,G48154,G48155,G48156,G48157,G48158,G48159,G48160,
       G48161,G48162,G48163,G48164,G48165,G48166,G48167,G48168,G48169,G48170,G48171,G48172,G48173,G48174,G48175,G48176,G48177,G48178,G48179,G48180,
       G48181,G48182,G48183,G48184,G48185,G48186,G48187,G48188,G48189,G48190,G48191,G48192,G48193,G48194,G48195,G48196,G48197,G48198,G48199,G48200,
       G48201,G48202,G48203,G48204,G48205,G48206,G48207,G48208,G48209,G48210,G48211,G48212,G48213,G48214,G48215,G48216,G48217,G48218,G48219,G48220,
       G48221,G48222,G48223,G48224,G48225,G48226,G48227,G48228,G48229,G48230,G48231,G48232,G48233,G48234,G48235,G48236,G48237,G48238,G48239,G48240,
       G48241,G48242,G48243,G48244,G48245,G48246,G48247,G48248,G48249,G48250,G48251,G48252,G48253,G48254,G48255,G48256,G48257,G48258,G48259,G48260,
       G48261,G48262,G48263,G48264,G48265,G48266,G48267,G48268,G48269,G48270,G48271,G48272,G48273,G48274,G48275,G48276,G48277,G48278,G48279,G48280,
       G48281,G48282,G48283,G48284,G48285,G48286,G48287,G48288,G48289,G48290,G48291,G48292,G48293,G48294,G48295,G48296,G48297,G48298,G48299,G48300,
       G48301,G48302,G48303,G48304,G48305,G48306,G48307,G48308,G48309,G48310,G48311,G48312,G48313,G48314,G48315,G48316,G48317,G48318,G48319,G48320,
       G48321,G48322,G48323,G48324,G48325,G48326,G48327,G48328,G48329,G48330,G48331,G48332,G48333,G48334,G48335,G48336,G48337,G48338,G48339,G48340,
       G48341,G48342,G48343,G48344,G48345,G48346,G48347,G48348,G48349,G48350,G48351,G48352,G48353,G48354,G48355,G48356,G48357,G48358,G48359,G48360,
       G48361,G48362,G48363,G48364,G48365,G48366,G48367,G48368,G48369,G48370,G48371,G48372,G48373,G48374,G48375,G48376,G48377,G48378,G48379,G48380,
       G48381,G48382,G48383,G48384,G48385,G48386,G48387,G48388,G48389,G48390,G48391,G48392,G48393,G48394,G48395,G48396,G48397,G48398,G48399,G48400,
       G48401,G48402,G48403,G48404,G48405,G48406,G48407,G48408,G48409,G48410,G48411,G48412,G48413,G48414,G48415,G48416,G48417,G48418,G48419,G48420,
       G48421,G48422,G48423,G48424,G48425,G48426,G48427,G48428,G48429,G48430,G48431,G48432,G48433,G48434,G48435,G48436,G48437,G48438,G48439,G48440,
       G48441,G48442,G48443,G48444,G48445,G48446,G48447,G48448,G48449,G48450,G48451,G48452,G48453,G48454,G48455,G48456,G48457,G48458,G48459,G48460,
       G48461,G48462,G48463,G48464,G48465,G48466,G48467,G48468,G48469,G48470,G48471,G48472,G48473,G48474,G48475,G48476,G48477,G48478,G48479,G48480,
       G48481,G48482,G48483,G48484,G48485,G48486,G48487,G48488,G48489,G48490,G48491,G48492,G48493,G48494,G48495,G48496,G48497,G48498,G48499,G48500,
       G48501,G48502,G48503,G48504,G48505,G48506,G48507,G48508,G48509,G48510,G48511,G48512,G48513,G48514,G48515,G48516,G48517,G48518,G48519,G48520,
       G48521,G48522,G48523,G48524,G48525,G48526,G48527,G48528,G48529,G48530,G48531,G48532,G48533,G48534,G48535,G48536,G48537,G48538,G48539,G48540,
       G48541,G48542,G48543,G48544,G48545,G48546,G48547,G48548,G48549,G48550,G48551,G48552,G48553,G48554,G48555,G48556,G48557,G48558,G48559,G48560,
       G48561,G48562,G48563,G48564,G48565,G48566,G48567,G48568,G48569,G48570,G48571,G48572,G48573,G48574,G48575,G48576,G48577,G48578,G48579,G48580,
       G48581,G48582,G48583,G48584,G48585,G48586,G48587,G48588,G48589,G48590,G48591,G48592,G48593,G48594,G48595,G48596,G48597,G48598,G48599,G48600,
       G48601,G48602,G48603,G48604,G48605,G48606,G48607,G48608,G48609,G48610,G48611,G48612,G48613,G48614,G48615,G48616,G48617,G48618,G48619,G48620,
       G48621,G48622,G48623,G48624,G48625,G48626,G48627,G48628,G48629,G48630,G48631,G48632,G48633,G48634,G48635,G48636,G48637,G48638,G48639,G48640,
       G48641,G48642,G48643,G48644,G48645,G48646,G48647,G48648,G48649,G48650,G48651,G48652,G48653,G48654,G48655,G48656,G48657,G48658,G48659,G48660,
       G48661,G48662,G48663,G48664,G48665,G48666,G48667,G48668,G48669,G48670,G48671,G48672,G48673,G48674,G48675,G48676,G48677,G48678,G48679,G48680,
       G48681,G48682,G48683,G48684,G48685,G48686,G48687,G48688,G48689,G48690,G48691,G48692,G48693,G48694,G48695,G48696,G48697,G48698,G48699,G48700,
       G48701,G48702,G48703,G48704,G48705,G48706,G48707,G48708,G48709,G48710,G48711,G48712,G48713,G48714,G48715,G48716,G48717,G48718,G48719,G48720,
       G48721,G48722,G48723,G48724,G48725,G48726,G48727,G48728,G48729,G48730,G48731,G48732,G48733,G48734,G48735,G48736,G48737,G48738,G48739,G48740,
       G48741,G48742,G48743,G48744,G48745,G48746,G48747,G48748,G48749,G48750,G48751,G48752,G48753,G48754,G48755,G48756,G48757,G48758,G48759,G48760,
       G48761,G48762,G48763,G48764,G48765,G48766,G48767,G48768,G48769,G48770,G48771,G48772,G48773,G48774,G48775,G48776,G48777,G48778,G48779,G48780,
       G48781,G48782,G48783,G48784,G48785,G48786,G48787,G48788,G48789,G48790,G48791,G48792,G48793,G48794,G48795,G48796,G48797,G48798,G48799,G48800,
       G48801,G48802,G48803,G48804,G48805,G48806,G48807,G48808,G48809,G48810,G48811,G48812,G48813,G48814,G48815,G48816,G48817,G48818,G48819,G48820,
       G48821,G48822,G48823,G48824,G48825,G48826,G48827,G48828,G48829,G48830,G48831,G48832,G48833,G48834,G48835,G48836,G48837,G48838,G48839,G48840,
       G48841,G48842,G48843,G48844,G48845,G48846,G48847,G48848,G48849,G48850,G48851,G48852,G48853,G48854,G48855,G48856,G48857,G48858,G48859,G48860,
       G48861,G48862,G48863,G48864,G48865,G48866,G48867,G48868,G48869,G48870,G48871,G48872,G48873,G48874,G48875,G48876,G48877,G48878,G48879,G48880,
       G48881,G48882,G48883,G48884,G48885,G48886,G48887,G48888,G48889,G48890,G48891,G48892,G48893,G48894,G48895,G48896,G48897,G48898,G48899,G48900,
       G48901,G48902,G48903,G48904,G48905,G48906,G48907,G48908,G48909,G48910,G48911,G48912,G48913,G48914,G48915,G48916,G48917,G48918,G48919,G48920,
       G48921,G48922,G48923,G48924,G48925,G48926,G48927,G48928,G48929,G48930,G48931,G48932,G48933,G48934,G48935,G48936,G48937,G48938,G48939,G48940,
       G48941,G48942,G48943,G48944,G48945,G48946,G48947,G48948,G48949,G48950,G48951,G48952,G48953,G48954,G48955,G48956,G48957,G48958,G48959,G48960,
       G48961,G48962,G48963,G48964,G48965,G48966,G48967,G48968,G48969,G48970,G48971,G48972,G48973,G48974,G48975,G48976,G48977,G48978,G48979,G48980,
       G48981,G48982,G48983,G48984,G48985,G48986,G48987,G48988,G48989,G48990,G48991,G48992,G48993,G48994,G48995,G48996,G48997,G48998,G48999,G49000,
       G49001,G49002,G49003,G49004,G49005,G49006,G49007,G49008,G49009,G49010,G49011,G49012,G49013,G49014,G49015,G49016,G49017,G49018,G49019,G49020,
       G49021,G49022,G49023,G49024,G49025,G49026,G49027,G49028,G49029,G49030,G49031,G49032,G49033,G49034,G49035,G49036,G49037,G49038,G49039,G49040,
       G49041,G49042,G49043,G49044,G49045,G49046,G49047,G49048,G49049,G49050,G49051,G49052,G49053,G49054,G49055,G49056,G49057,G49058,G49059,G49060,
       G49061,G49062,G49063,G49064,G49065,G49066,G49067,G49068,G49069,G49070,G49071,G49072,G49073,G49074,G49075,G49076,G49077,G49078,G49079,G49080,
       G49081,G49082,G49083,G49084,G49085,G49086,G49087,G49088,G49089,G49090,G49091,G49092,G49093,G49094,G49095,G49096,G49097,G49098,G49099,G49100,
       G49101,G49102,G49103,G49104,G49105,G49106,G49107,G49108,G49109,G49110,G49111,G49112,G49113,G49114,G49115,G49116,G49117,G49118,G49119,G49120,
       G49121,G49122,G49123,G49124,G49125,G49126,G49127,G49128,G49129,G49130,G49131,G49132,G49133,G49134,G49135,G49136,G49137,G49138,G49139,G49140,
       G49141,G49142,G49143,G49144,G49145,G49146,G49147,G49148,G49149,G49150,G49151,G49152,G49153,G49154,G49155,G49156,G49157,G49158,G49159,G49160,
       G49161,G49162,G49163,G49164,G49165,G49166,G49167,G49168,G49169,G49170,G49171,G49172,G49173,G49174,G49175,G49176,G49177,G49178,G49179,G49180,
       G49181,G49182,G49183,G49184,G49185,G49186,G49187,G49188,G49189,G49190,G49191,G49192,G49193,G49194,G49195,G49196,G49197,G49198,G49199,G49200,
       G49201,G49202,G49203,G49204,G49205,G49206,G49207,G49208,G49209,G49210,G49211,G49212,G49213,G49214,G49215,G49216,G49217,G49218,G49219,G49220,
       G49221,G49222,G49223,G49224,G49225,G49226,G49227,G49228,G49229,G49230,G49231,G49232,G49233,G49234,G49235,G49236,G49237,G49238,G49239,G49240,
       G49241,G49242,G49243,G49244,G49245,G49246,G49247,G49248,G49249,G49250,G49251,G49252,G49253,G49254,G49255,G49256,G49257,G49258,G49259,G49260,
       G49261,G49262,G49263,G49264,G49265,G49266,G49267,G49268,G49269,G49270,G49271,G49272,G49273,G49274,G49275,G49276,G49277,G49278,G49279,G49280,
       G49281,G49282,G49283,G49284,G49285,G49286,G49287,G49288,G49289,G49290,G49291,G49292,G49293,G49294,G49295,G49296,G49297,G49298,G49299,G49300,
       G49301,G49302,G49303,G49304,G49305,G49306,G49307,G49308,G49309,G49310,G49311,G49312,G49313,G49314,G49315,G49316,G49317,G49318,G49319,G49320,
       G49321,G49322,G49323,G49324,G49325,G49326,G49327,G49328,G49329,G49330,G49331,G49332,G49333,G49334,G49335,G49336,G49337,G49338,G49339,G49340,
       G49341,G49342,G49343,G49344,G49345,G49346,G49347,G49348,G49349,G49350,G49351,G49352,G49353,G49354,G49355,G49356,G49357,G49358,G49359,G49360,
       G49361,G49362,G49363,G49364,G49365,G49366,G49367,G49368,G49369,G49370,G49371,G49372,G49373,G49374,G49375,G49376,G49377,G49378,G49379,G49380,
       G49381,G49382,G49383,G49384,G49385,G49386,G49387,G49388,G49389,G49390,G49391,G49392,G49393,G49394,G49395,G49396,G49397,G49398,G49399,G49400,
       G49401,G49402,G49403,G49404,G49405,G49406,G49407,G49408,G49409,G49410,G49411,G49412,G49413,G49414,G49415,G49416,G49417,G49418,G49419,G49420,
       G49421,G49422,G49423,G49424,G49425,G49426,G49427,G49428,G49429,G49430,G49431,G49432,G49433,G49434,G49435,G49436,G49437,G49438,G49439,G49440,
       G49441,G49442,G49443,G49444,G49445,G49446,G49447,G49448,G49449,G49450,G49451,G49452,G49453,G49454,G49455,G49456,G49457,G49458,G49459,G49460,
       G49461,G49462,G49463,G49464,G49465,G49466,G49467,G49468,G49469,G49470,G49471,G49472,G49473,G49474,G49475,G49476,G49477,G49478,G49479,G49480,
       G49481,G49482,G49483,G49484,G49485,G49486,G49487,G49488,G49489,G49490,G49491,G49492,G49493,G49494,G49495,G49496,G49497,G49498,G49499,G49500,
       G49501,G49502,G49503,G49504,G49505,G49506,G49507,G49508,G49509,G49510,G49511,G49512,G49513,G49514,G49515,G49516,G49517,G49518,G49519,G49520,
       G49521,G49522,G49523,G49524,G49525,G49526,G49527,G49528,G49529,G49530,G49531,G49532,G49533,G49534,G49535,G49536,G49537,G49538,G49539,G49540,
       G49541,G49542,G49543,G49544,G49545,G49546,G49547,G49548,G49549,G49550,G49551,G49552,G49553,G49554,G49555,G49556,G49557,G49558,G49559,G49560,
       G49561,G49562,G49563,G49564,G49565,G49566,G49567,G49568,G49569,G49570,G49571,G49572,G49573,G49574,G49575,G49576,G49577,G49578,G49579,G49580,
       G49581,G49582,G49583,G49584,G49585,G49586,G49587,G49588,G49589,G49590,G49591,G49592,G49593,G49594,G49595,G49596,G49597,G49598,G49599,G49600,
       G49601,G49602,G49603,G49604,G49605,G49606,G49607,G49608,G49609,G49610,G49611,G49612,G49613,G49614,G49615,G49616,G49617,G49618,G49619,G49620,
       G49621,G49622,G49623,G49624,G49625,G49626,G49627,G49628,G49629,G49630,G49631,G49632,G49633,G49634,G49635,G49636,G49637,G49638,G49639,G49640,
       G49641,G49642,G49643,G49644,G49645,G49646,G49647,G49648,G49649,G49650,G49651,G49652,G49653,G49654,G49655,G49656,G49657,G49658,G49659,G49660,
       G49661,G49662,G49663,G49664,G49665,G49666,G49667,G49668,G49669,G49670,G49671,G49672,G49673,G49674,G49675,G49676,G49677,G49678,G49679,G49680,
       G49681,G49682,G49683,G49684,G49685,G49686,G49687,G49688,G49689,G49690,G49691,G49692,G49693,G49694,G49695,G49696,G49697,G49698,G49699,G49700,
       G49701,G49702,G49703,G49704,G49705,G49706,G49707,G49708,G49709,G49710,G49711,G49712,G49713,G49714,G49715,G49716,G49717,G49718,G49719,G49720,
       G49721,G49722,G49723,G49724,G49725,G49726,G49727,G49728,G49729,G49730,G49731,G49732,G49733,G49734,G49735,G49736,G49737,G49738,G49739,G49740,
       G49741,G49742,G49743,G49744,G49745,G49746,G49747,G49748,G49749,G49750,G49751,G49752,G49753,G49754,G49755,G49756,G49757,G49758,G49759,G49760,
       G49761,G49762,G49763,G49764,G49765,G49766,G49767,G49768,G49769,G49770,G49771,G49772,G49773,G49774,G49775,G49776,G49777,G49778,G49779,G49780,
       G49781,G49782,G49783,G49784,G49785,G49786,G49787,G49788,G49789,G49790,G49791,G49792,G49793,G49794,G49795,G49796,G49797,G49798,G49799,G49800,
       G49801,G49802,G49803,G49804,G49805,G49806,G49807,G49808,G49809,G49810,G49811,G49812,G49813,G49814,G49815,G49816,G49817,G49818,G49819,G49820,
       G49821,G49822,G49823,G49824,G49825,G49826,G49827,G49828,G49829,G49830,G49831,G49832,G49833,G49834,G49835,G49836,G49837,G49838,G49839,G49840,
       G49841,G49842,G49843,G49844,G49845,G49846,G49847,G49848,G49849,G49850,G49851,G49852,G49853,G49854,G49855,G49856,G49857,G49858,G49859,G49860,
       G49861,G49862,G49863,G49864,G49865,G49866,G49867,G49868,G49869,G49870,G49871,G49872,G49873,G49874,G49875,G49876,G49877,G49878,G49879,G49880,
       G49881,G49882,G49883,G49884,G49885,G49886,G49887,G49888,G49889,G49890,G49891,G49892,G49893,G49894,G49895,G49896,G49897,G49898,G49899,G49900,
       G49901,G49902,G49903,G49904,G49905,G49906,G49907,G49908,G49909,G49910,G49911,G49912,G49913,G49914,G49915,G49916,G49917,G49918,G49919,G49920,
       G49921,G49922,G49923,G49924,G49925,G49926,G49927,G49928,G49929,G49930,G49931,G49932,G49933,G49934,G49935,G49936,G49937,G49938,G49939,G49940,
       G49941,G49942,G49943,G49944,G49945,G49946,G49947,G49948,G49949,G49950,G49951,G49952,G49953,G49954,G49955,G49956,G49957,G49958,G49959,G49960,
       G49961,G49962,G49963,G49964,G49965,G49966,G49967,G49968,G49969,G49970,G49971,G49972,G49973,G49974,G49975,G49976,G49977,G49978,G49979,G49980,
       G49981,G49982,G49983,G49984,G49985,G49986,G49987,G49988,G49989,G49990,G49991,G49992,G49993,G49994,G49995,G49996,G49997,G49998,G49999,G50000,
       G50001,G50002,G50003,G50004,G50005,G50006,G50007,G50008,G50009,G50010,G50011,G50012,G50013,G50014,G50015,G50016,G50017,G50018,G50019,G50020,
       G50021,G50022,G50023,G50024,G50025,G50026,G50027,G50028,G50029,G50030,G50031,G50032,G50033,G50034,G50035,G50036,G50037,G50038,G50039,G50040,
       G50041,G50042,G50043,G50044,G50045,G50046,G50047,G50048,G50049,G50050,G50051,G50052,G50053,G50054,G50055,G50056,G50057,G50058,G50059,G50060,
       G50061,G50062,G50063,G50064,G50065,G50066,G50067,G50068,G50069,G50070,G50071,G50072,G50073,G50074,G50075,G50076,G50077,G50078,G50079,G50080,
       G50081,G50082,G50083,G50084,G50085,G50086,G50087,G50088,G50089,G50090,G50091,G50092,G50093,G50094,G50095,G50096,G50097,G50098,G50099,G50100,
       G50101,G50102,G50103,G50104,G50105,G50106,G50107,G50108,G50109,G50110,G50111,G50112,G50113,G50114,G50115,G50116,G50117,G50118,G50119,G50120,
       G50121,G50122,G50123,G50124,G50125,G50126,G50127,G50128,G50129,G50130,G50131,G50132,G50133,G50134,G50135,G50136,G50137,G50138,G50139,G50140,
       G50141,G50142,G50143,G50144,G50145,G50146,G50147,G50148,G50149,G50150,G50151,G50152,G50153,G50154,G50155,G50156,G50157,G50158,G50159,G50160,
       G50161,G50162,G50163,G50164,G50165,G50166,G50167,G50168,G50169,G50170,G50171,G50172,G50173,G50174,G50175,G50176,G50177,G50178,G50179,G50180,
       G50181,G50182,G50183,G50184,G50185,G50186,G50187,G50188,G50189,G50190,G50191,G50192,G50193,G50194,G50195,G50196,G50197,G50198,G50199,G50200,
       G50201,G50202,G50203,G50204,G50205,G50206,G50207,G50208,G50209,G50210,G50211,G50212,G50213,G50214,G50215,G50216,G50217,G50218,G50219,G50220,
       G50221,G50222,G50223,G50224,G50225,G50226,G50227,G50228,G50229,G50230,G50231,G50232,G50233,G50234,G50235,G50236,G50237,G50238,G50239,G50240,
       G50241,G50242,G50243,G50244,G50245,G50246,G50247,G50248,G50249,G50250,G50251,G50252,G50253,G50254,G50255,G50256,G50257,G50258,G50259,G50260,
       G50261,G50262,G50263,G50264,G50265,G50266,G50267,G50268,G50269,G50270,G50271,G50272,G50273,G50274,G50275,G50276,G50277,G50278,G50279,G50280,
       G50281,G50282,G50283,G50284,G50285,G50286,G50287,G50288,G50289,G50290,G50291,G50292,G50293,G50294,G50295,G50296,G50297,G50298,G50299,G50300,
       G50301,G50302,G50303,G50304,G50305,G50306,G50307,G50308,G50309,G50310,G50311,G50312,G50313,G50314,G50315,G50316,G50317,G50318,G50319,G50320,
       G50321,G50322,G50323,G50324,G50325,G50326,G50327,G50328,G50329,G50330,G50331,G50332,G50333,G50334,G50335,G50336,G50337,G50338,G50339,G50340,
       G50341,G50342,G50343,G50344,G50345,G50346,G50347,G50348,G50349,G50350,G50351,G50352,G50353,G50354,G50355,G50356,G50357,G50358,G50359,G50360,
       G50361,G50362,G50363,G50364,G50365,G50366,G50367,G50368,G50369,G50370,G50371,G50372,G50373,G50374,G50375,G50376,G50377,G50378,G50379,G50380,
       G50381,G50382,G50383,G50384,G50385,G50386,G50387,G50388,G50389,G50390,G50391,G50392,G50393,G50394,G50395,G50396,G50397,G50398,G50399,G50400,
       G50401,G50402,G50403,G50404,G50405,G50406,G50407,G50408,G50409,G50410,G50411,G50412,G50413,G50414,G50415,G50416,G50417,G50418,G50419,G50420,
       G50421,G50422,G50423,G50424,G50425,G50426,G50427,G50428,G50429,G50430,G50431,G50432,G50433,G50434,G50435,G50436,G50437,G50438,G50439,G50440,
       G50441,G50442,G50443,G50444,G50445,G50446,G50447,G50448,G50449,G50450,G50451,G50452,G50453,G50454,G50455,G50456,G50457,G50458,G50459,G50460,
       G50461,G50462,G50463,G50464,G50465,G50466,G50467,G50468,G50469,G50470,G50471,G50472,G50473,G50474,G50475,G50476,G50477,G50478,G50479,G50480,
       G50481,G50482,G50483,G50484,G50485,G50486,G50487,G50488,G50489,G50490,G50491,G50492,G50493,G50494,G50495,G50496,G50497,G50498,G50499,G50500,
       G50501,G50502,G50503,G50504,G50505,G50506,G50507,G50508,G50509,G50510,G50511,G50512,G50513,G50514,G50515,G50516,G50517,G50518,G50519,G50520,
       G50521,G50522,G50523,G50524,G50525,G50526,G50527,G50528,G50529,G50530,G50531,G50532,G50533,G50534,G50535,G50536,G50537,G50538,G50539,G50540,
       G50541,G50542,G50543,G50544,G50545,G50546,G50547,G50548,G50549,G50550,G50551,G50552,G50553,G50554,G50555,G50556,G50557,G50558,G50559,G50560,
       G50561,G50562,G50563,G50564,G50565,G50566,G50567,G50568,G50569,G50570,G50571,G50572,G50573,G50574,G50575,G50576,G50577,G50578,G50579,G50580,
       G50581,G50582,G50583,G50584,G50585,G50586,G50587,G50588,G50589,G50590,G50591,G50592,G50593,G50594,G50595,G50596,G50597,G50598,G50599,G50600,
       G50601,G50602,G50603,G50604,G50605,G50606,G50607,G50608,G50609,G50610,G50611,G50612,G50613,G50614,G50615,G50616,G50617,G50618,G50619,G50620,
       G50621,G50622,G50623,G50624,G50625,G50626,G50627,G50628,G50629,G50630,G50631,G50632,G50633,G50634,G50635,G50636,G50637,G50638,G50639,G50640,
       G50641,G50642,G50643,G50644,G50645,G50646,G50647,G50648,G50649,G50650,G50651,G50652,G50653,G50654,G50655,G50656,G50657,G50658,G50659,G50660,
       G50661,G50662,G50663,G50664,G50665,G50666,G50667,G50668,G50669,G50670,G50671,G50672,G50673,G50674,G50675,G50676,G50677,G50678,G50679,G50680,
       G50681,G50682,G50683,G50684,G50685,G50686,G50687,G50688,G50689,G50690,G50691,G50692,G50693,G50694,G50695,G50696,G50697,G50698,G50699,G50700,
       G50701,G50702,G50703,G50704,G50705,G50706,G50707,G50708,G50709,G50710,G50711,G50712,G50713,G50714,G50715,G50716,G50717,G50718,G50719,G50720,
       G50721,G50722,G50723,G50724,G50725,G50726,G50727,G50728,G50729,G50730,G50731,G50732,G50733,G50734,G50735,G50736,G50737,G50738,G50739,G50740,
       G50741,G50742,G50743,G50744,G50745,G50746,G50747,G50748,G50749,G50750,G50751,G50752,G50753,G50754,G50755,G50756,G50757,G50758,G50759,G50760,
       G50761,G50762,G50763,G50764,G50765,G50766,G50767,G50768,G50769,G50770,G50771,G50772,G50773,G50774,G50775,G50776,G50777,G50778,G50779,G50780,
       G50781,G50782,G50783,G50784,G50785,G50786,G50787,G50788,G50789,G50790,G50791,G50792,G50793,G50794,G50795,G50796,G50797,G50798,G50799,G50800,
       G50801,G50802,G50803,G50804,G50805,G50806,G50807,G50808,G50809,G50810,G50811,G50812,G50813,G50814,G50815,G50816,G50817,G50818,G50819,G50820,
       G50821,G50822,G50823,G50824,G50825,G50826,G50827,G50828,G50829,G50830,G50831,G50832,G50833,G50834,G50835,G50836,G50837,G50838,G50839,G50840,
       G50841,G50842,G50843,G50844,G50845,G50846,G50847,G50848,G50849,G50850,G50851,G50852,G50853,G50854,G50855,G50856,G50857,G50858,G50859,G50860,
       G50861,G50862,G50863,G50864,G50865,G50866,G50867,G50868,G50869,G50870,G50871,G50872,G50873,G50874,G50875,G50876,G50877,G50878,G50879,G50880,
       G50881,G50882,G50883,G50884,G50885,G50886,G50887,G50888,G50889,G50890,G50891,G50892,G50893,G50894,G50895,G50896,G50897,G50898,G50899,G50900,
       G50901,G50902,G50903,G50904,G50905,G50906,G50907,G50908,G50909,G50910,G50911,G50912,G50913,G50914,G50915,G50916,G50917,G50918,G50919,G50920,
       G50921,G50922,G50923,G50924,G50925,G50926,G50927,G50928,G50929,G50930,G50931,G50932,G50933,G50934,G50935,G50936,G50937,G50938,G50939,G50940,
       G50941,G50942,G50943,G50944,G50945,G50946,G50947,G50948,G50949,G50950,G50951,G50952,G50953,G50954,G50955,G50956,G50957,G50958,G50959,G50960,
       G50961,G50962,G50963,G50964,G50965,G50966,G50967,G50968,G50969,G50970,G50971,G50972,G50973,G50974,G50975,G50976,G50977,G50978,G50979,G50980,
       G50981,G50982,G50983,G50984,G50985,G50986,G50987,G50988,G50989,G50990,G50991,G50992,G50993,G50994,G50995,G50996,G50997,G50998,G50999,G51000,
       G51001,G51002,G51003,G51004,G51005,G51006,G51007,G51008,G51009,G51010,G51011,G51012,G51013,G51014,G51015,G51016,G51017,G51018,G51019,G51020,
       G51021,G51022,G51023,G51024,G51025,G51026,G51027,G51028,G51029,G51030,G51031,G51032,G51033,G51034,G51035,G51036,G51037,G51038,G51039,G51040,
       G51041,G51042,G51043,G51044,G51045,G51046,G51047,G51048,G51049,G51050,G51051,G51052,G51053,G51054,G51055,G51056,G51057,G51058,G51059,G51060,
       G51061,G51062,G51063,G51064,G51065,G51066,G51067,G51068,G51069,G51070,G51071,G51072,G51073,G51074,G51075,G51076,G51077,G51078,G51079,G51080,
       G51081,G51082,G51083,G51084,G51085,G51086,G51087,G51088,G51089,G51090,G51091,G51092,G51093,G51094,G51095,G51096,G51097,G51098,G51099,G51100,
       G51101,G51102,G51103,G51104,G51105,G51106,G51107,G51108,G51109,G51110,G51111,G51112,G51113,G51114,G51115,G51116,G51117,G51118,G51119,G51120,
       G51121,G51122,G51123,G51124,G51125,G51126,G51127,G51128,G51129,G51130,G51131,G51132,G51133,G51134,G51135,G51136,G51137,G51138,G51139,G51140,
       G51141,G51142,G51143,G51144,G51145,G51146,G51147,G51148,G51149,G51150,G51151,G51152,G51153,G51154,G51155,G51156,G51157,G51158,G51159,G51160,
       G51161,G51162,G51163,G51164,G51165,G51166,G51167,G51168,G51169,G51170,G51171,G51172,G51173,G51174,G51175,G51176,G51177,G51178,G51179,G51180,
       G51181,G51182,G51183,G51184,G51185,G51186,G51187,G51188,G51189,G51190,G51191,G51192,G51193,G51194,G51195,G51196,G51197,G51198,G51199,G51200,
       G51201,G51202,G51203,G51204,G51205,G51206,G51207,G51208,G51209,G51210,G51211,G51212,G51213,G51214,G51215,G51216,G51217,G51218,G51219,G51220,
       G51221,G51222,G51223,G51224,G51225,G51226,G51227,G51228,G51229,G51230,G51231,G51232,G51233,G51234,G51235,G51236,G51237,G51238,G51239,G51240,
       G51241,G51242,G51243,G51244,G51245,G51246,G51247,G51248,G51249,G51250,G51251,G51252,G51253,G51254,G51255,G51256,G51257,G51258,G51259,G51260,
       G51261,G51262,G51263,G51264,G51265,G51266,G51267,G51268,G51269,G51270,G51271,G51272,G51273,G51274,G51275,G51276,G51277,G51278,G51279,G51280,
       G51281,G51282,G51283,G51284,G51285,G51286,G51287,G51288,G51289,G51290,G51291,G51292,G51293,G51294,G51295,G51296,G51297,G51298,G51299,G51300,
       G51301,G51302,G51303,G51304,G51305,G51306,G51307,G51308,G51309,G51310,G51311,G51312,G51313,G51314,G51315,G51316,G51317,G51318,G51319,G51320,
       G51321,G51322,G51323,G51324,G51325,G51326,G51327,G51328,G51329,G51330,G51331,G51332,G51333,G51334,G51335,G51336,G51337,G51338,G51339,G51340,
       G51341,G51342,G51343,G51344,G51345,G51346,G51347,G51348,G51349,G51350,G51351,G51352,G51353,G51354,G51355,G51356,G51357,G51358,G51359,G51360,
       G51361,G51362,G51363,G51364,G51365,G51366,G51367,G51368,G51369,G51370,G51371,G51372,G51373,G51374,G51375,G51376,G51377,G51378,G51379,G51380,
       G51381,G51382,G51383,G51384,G51385,G51386,G51387,G51388,G51389,G51390,G51391,G51392,G51393,G51394,G51395,G51396,G51397,G51398,G51399,G51400,
       G51401,G51402,G51403,G51404,G51405,G51406,G51407,G51408,G51409,G51410,G51411,G51412,G51413,G51414,G51415,G51416,G51417,G51418,G51419,G51420,
       G51421,G51422,G51423,G51424,G51425,G51426,G51427,G51428,G51429,G51430,G51431,G51432,G51433,G51434,G51435,G51436,G51437,G51438,G51439,G51440,
       G51441,G51442,G51443,G51444,G51445,G51446,G51447,G51448,G51449,G51450,G51451,G51452,G51453,G51454,G51455,G51456,G51457,G51458,G51459,G51460,
       G51461,G51462,G51463,G51464,G51465,G51466,G51467,G51468,G51469,G51470,G51471,G51472,G51473,G51474,G51475,G51476,G51477,G51478,G51479,G51480,
       G51481,G51482,G51483,G51484,G51485,G51486,G51487,G51488,G51489,G51490,G51491,G51492,G51493,G51494,G51495,G51496,G51497,G51498,G51499,G51500,
       G51501,G51502,G51503,G51504,G51505,G51506,G51507,G51508,G51509,G51510,G51511,G51512,G51513,G51514,G51515,G51516,G51517,G51518,G51519,G51520,
       G51521,G51522,G51523,G51524,G51525,G51526,G51527,G51528,G51529,G51530,G51531,G51532,G51533,G51534,G51535,G51536,G51537,G51538,G51539,G51540,
       G51541,G51542,G51543,G51544,G51545,G51546,G51547,G51548,G51549,G51550,G51551,G51552,G51553,G51554,G51555,G51556,G51557,G51558,G51559,G51560,
       G51561,G51562,G51563,G51564,G51565,G51566,G51567,G51568,G51569,G51570,G51571,G51572,G51573,G51574,G51575,G51576,G51577,G51578,G51579,G51580,
       G51581,G51582,G51583,G51584,G51585,G51586,G51587,G51588,G51589,G51590,G51591,G51592,G51593,G51594,G51595,G51596,G51597,G51598,G51599,G51600,
       G51601,G51602,G51603,G51604,G51605,G51606,G51607,G51608,G51609,G51610,G51611,G51612,G51613,G51614,G51615,G51616,G51617,G51618,G51619,G51620,
       G51621,G51622,G51623,G51624,G51625,G51626,G51627,G51628,G51629,G51630,G51631,G51632,G51633,G51634,G51635,G51636,G51637,G51638,G51639,G51640,
       G51641,G51642,G51643,G51644,G51645,G51646,G51647,G51648,G51649,G51650,G51651,G51652,G51653,G51654,G51655,G51656,G51657,G51658,G51659,G51660,
       G51661,G51662,G51663,G51664,G51665,G51666,G51667,G51668,G51669,G51670,G51671,G51672,G51673,G51674,G51675,G51676,G51677,G51678,G51679,G51680,
       G51681,G51682,G51683,G51684,G51685,G51686,G51687,G51688,G51689,G51690,G51691,G51692,G51693,G51694,G51695,G51696,G51697,G51698,G51699,G51700,
       G51701,G51702,G51703,G51704,G51705,G51706,G51707,G51708,G51709,G51710,G51711,G51712,G51713,G51714,G51715,G51716,G51717,G51718,G51719,G51720,
       G51721,G51722,G51723,G51724,G51725,G51726,G51727,G51728,G51729,G51730,G51731,G51732,G51733,G51734,G51735,G51736,G51737,G51738,G51739,G51740,
       G51741,G51742,G51743,G51744,G51745,G51746,G51747,G51748,G51749,G51750,G51751,G51752,G51753,G51754,G51755,G51756,G51757,G51758,G51759,G51760,
       G51761,G51762,G51763,G51764,G51765,G51766,G51767,G51768,G51769,G51770,G51771,G51772,G51773,G51774,G51775,G51776,G51777,G51778,G51779,G51780,
       G51781,G51782,G51783,G51784,G51785,G51786,G51787,G51788,G51789,G51790,G51791,G51792,G51793,G51794,G51795,G51796,G51797,G51798,G51799,G51800,
       G51801,G51802,G51803,G51804,G51805,G51806,G51807,G51808,G51809,G51810,G51811,G51812,G51813,G51814,G51815,G51816,G51817,G51818,G51819,G51820,
       G51821,G51822,G51823,G51824,G51825,G51826,G51827,G51828,G51829,G51830,G51831,G51832,G51833,G51834,G51835,G51836,G51837,G51838,G51839,G51840,
       G51841,G51842,G51843,G51844,G51845,G51846,G51847,G51848,G51849,G51850,G51851,G51852,G51853,G51854,G51855,G51856,G51857,G51858,G51859,G51860,
       G51861,G51862,G51863,G51864,G51865,G51866,G51867,G51868,G51869,G51870,G51871,G51872,G51873,G51874,G51875,G51876,G51877,G51878,G51879,G51880,
       G51881,G51882,G51883,G51884,G51885,G51886,G51887,G51888,G51889,G51890,G51891,G51892,G51893,G51894,G51895,G51896,G51897,G51898,G51899,G51900,
       G51901,G51902,G51903,G51904,G51905,G51906,G51907,G51908,G51909,G51910,G51911,G51912,G51913,G51914,G51915,G51916,G51917,G51918,G51919,G51920,
       G51921,G51922,G51923,G51924,G51925,G51926,G51927,G51928,G51929,G51930,G51931,G51932,G51933,G51934,G51935,G51936,G51937,G51938,G51939,G51940,
       G51941,G51942,G51943,G51944,G51945,G51946,G51947,G51948,G51949,G51950,G51951,G51952,G51953,G51954,G51955,G51956,G51957,G51958,G51959,G51960,
       G51961,G51962,G51963,G51964,G51965,G51966,G51967,G51968,G51969,G51970,G51971,G51972,G51973,G51974,G51975,G51976,G51977,G51978,G51979,G51980,
       G51981,G51982,G51983,G51984,G51985,G51986,G51987,G51988,G51989,G51990,G51991,G51992,G51993,G51994,G51995,G51996,G51997,G51998,G51999,G52000,
       G52001,G52002,G52003,G52004,G52005,G52006,G52007,G52008,G52009,G52010,G52011,G52012,G52013,G52014,G52015,G52016,G52017,G52018,G52019,G52020,
       G52021,G52022,G52023,G52024,G52025,G52026,G52027,G52028,G52029,G52030,G52031,G52032,G52033,G52034,G52035,G52036,G52037,G52038,G52039,G52040,
       G52041,G52042,G52043,G52044,G52045,G52046,G52047,G52048,G52049,G52050,G52051,G52052,G52053,G52054,G52055,G52056,G52057,G52058,G52059,G52060,
       G52061,G52062,G52063,G52064,G52065,G52066,G52067,G52068,G52069,G52070,G52071,G52072,G52073,G52074,G52075,G52076,G52077,G52078,G52079,G52080,
       G52081,G52082,G52083,G52084,G52085,G52086,G52087,G52088,G52089,G52090,G52091,G52092,G52093,G52094,G52095,G52096,G52097,G52098,G52099,G52100,
       G52101,G52102,G52103,G52104,G52105,G52106,G52107,G52108,G52109,G52110,G52111,G52112,G52113,G52114,G52115,G52116,G52117,G52118,G52119,G52120,
       G52121,G52122,G52123,G52124,G52125,G52126,G52127,G52128,G52129,G52130,G52131,G52132,G52133,G52134,G52135,G52136,G52137,G52138,G52139,G52140,
       G52141,G52142,G52143,G52144,G52145,G52146,G52147,G52148,G52149,G52150,G52151,G52152,G52153,G52154,G52155,G52156,G52157,G52158,G52159,G52160,
       G52161,G52162,G52163,G52164,G52165,G52166,G52167,G52168,G52169,G52170,G52171,G52172,G52173,G52174,G52175,G52176,G52177,G52178,G52179,G52180,
       G52181,G52182,G52183,G52184,G52185,G52186,G52187,G52188,G52189,G52190,G52191,G52192,G52193,G52194,G52195,G52196,G52197,G52198,G52199,G52200,
       G52201,G52202,G52203,G52204,G52205,G52206,G52207,G52208,G52209,G52210,G52211,G52212,G52213,G52214,G52215,G52216,G52217,G52218,G52219,G52220,
       G52221,G52222,G52223,G52224,G52225,G52226,G52227,G52228,G52229,G52230,G52231,G52232,G52233,G52234,G52235,G52236,G52237,G52238,G52239,G52240,
       G52241,G52242,G52243,G52244,G52245,G52246,G52247,G52248,G52249,G52250,G52251,G52252,G52253,G52254,G52255,G52256,G52257,G52258,G52259,G52260,
       G52261,G52262,G52263,G52264,G52265,G52266,G52267,G52268,G52269,G52270,G52271,G52272,G52273,G52274,G52275,G52276,G52277,G52278,G52279,G52280,
       G52281,G52282,G52283,G52284,G52285,G52286,G52287,G52288,G52289,G52290,G52291,G52292,G52293,G52294,G52295,G52296,G52297,G52298,G52299,G52300,
       G52301,G52302,G52303,G52304,G52305,G52306,G52307,G52308,G52309,G52310,G52311,G52312,G52313,G52314,G52315,G52316,G52317,G52318,G52319,G52320,
       G52321,G52322,G52323,G52324,G52325,G52326,G52327,G52328,G52329,G52330,G52331,G52332,G52333,G52334,G52335,G52336,G52337,G52338,G52339,G52340,
       G52341,G52342,G52343,G52344,G52345,G52346,G52347,G52348,G52349,G52350,G52351,G52352,G52353,G52354,G52355,G52356,G52357,G52358,G52359,G52360,
       G52361,G52362,G52363,G52364,G52365,G52366,G52367,G52368,G52369,G52370,G52371,G52372,G52373,G52374,G52375,G52376,G52377,G52378,G52379,G52380,
       G52381,G52382,G52383,G52384,G52385,G52386,G52387,G52388,G52389,G52390,G52391,G52392,G52393,G52394,G52395,G52396,G52397,G52398,G52399,G52400,
       G52401,G52402,G52403,G52404,G52405,G52406,G52407,G52408,G52409,G52410,G52411,G52412,G52413,G52414,G52415,G52416,G52417,G52418,G52419,G52420,
       G52421,G52422,G52423,G52424,G52425,G52426,G52427,G52428,G52429,G52430,G52431,G52432,G52433,G52434,G52435,G52436,G52437,G52438,G52439,G52440,
       G52441,G52442,G52443,G52444,G52445,G52446,G52447,G52448,G52449,G52450,G52451,G52452,G52453,G52454,G52455,G52456,G52457,G52458,G52459,G52460,
       G52461,G52462,G52463,G52464,G52465,G52466,G52467,G52468,G52469,G52470,G52471,G52472,G52473,G52474,G52475,G52476,G52477,G52478,G52479,G52480,
       G52481,G52482,G52483,G52484,G52485,G52486,G52487,G52488,G52489,G52490,G52491,G52492,G52493,G52494,G52495,G52496,G52497,G52498,G52499,G52500,
       G52501,G52502,G52503,G52504,G52505,G52506,G52507,G52508,G52509,G52510,G52511,G52512,G52513,G52514,G52515,G52516,G52517,G52518,G52519,G52520,
       G52521,G52522,G52523,G52524,G52525,G52526,G52527,G52528,G52529,G52530,G52531,G52532,G52533,G52534,G52535,G52536,G52537,G52538,G52539,G52540,
       G52541,G52542,G52543,G52544,G52545,G52546,G52547,G52548,G52549,G52550,G52551,G52552,G52553,G52554,G52555,G52556,G52557,G52558,G52559,G52560,
       G52561,G52562,G52563,G52564,G52565,G52566,G52567,G52568,G52569,G52570,G52571,G52572,G52573,G52574,G52575,G52576,G52577,G52578,G52579,G52580,
       G52581,G52582,G52583,G52584,G52585,G52586,G52587,G52588,G52589,G52590,G52591,G52592,G52593,G52594,G52595,G52596,G52597,G52598,G52599,G52600,
       G52601,G52602,G52603,G52604,G52605,G52606,G52607,G52608,G52609,G52610,G52611,G52612,G52613,G52614,G52615,G52616,G52617,G52618,G52619,G52620,
       G52621,G52622,G52623,G52624,G52625,G52626,G52627,G52628,G52629,G52630,G52631,G52632,G52633,G52634,G52635,G52636,G52637,G52638,G52639,G52640,
       G52641,G52642,G52643,G52644,G52645,G52646,G52647,G52648,G52649,G52650,G52651,G52652,G52653,G52654,G52655,G52656,G52657,G52658,G52659,G52660,
       G52661,G52662,G52663,G52664,G52665,G52666,G52667,G52668,G52669,G52670,G52671,G52672,G52673,G52674,G52675,G52676,G52677,G52678,G52679,G52680,
       G52681,G52682,G52683,G52684,G52685,G52686,G52687,G52688,G52689,G52690,G52691,G52692,G52693,G52694,G52695,G52696,G52697,G52698,G52699,G52700,
       G52701,G52702,G52703,G52704,G52705,G52706,G52707,G52708,G52709,G52710,G52711,G52712,G52713,G52714,G52715,G52716,G52717,G52718,G52719,G52720,
       G52721,G52722,G52723,G52724,G52725,G52726,G52727,G52728,G52729,G52730,G52731,G52732,G52733,G52734,G52735,G52736,G52737,G52738,G52739,G52740,
       G52741,G52742,G52743,G52744,G52745,G52746,G52747,G52748,G52749,G52750,G52751,G52752,G52753,G52754,G52755,G52756,G52757,G52758,G52759,G52760,
       G52761,G52762,G52763,G52764,G52765,G52766,G52767,G52768,G52769,G52770,G52771,G52772,G52773,G52774,G52775,G52776,G52777,G52778,G52779,G52780,
       G52781,G52782,G52783,G52784,G52785,G52786,G52787,G52788,G52789,G52790,G52791,G52792,G52793,G52794,G52795,G52796,G52797,G52798,G52799,G52800,
       G52801,G52802,G52803,G52804,G52805,G52806,G52807,G52808,G52809,G52810,G52811,G52812,G52813,G52814,G52815,G52816,G52817,G52818,G52819,G52820,
       G52821,G52822,G52823,G52824,G52825,G52826,G52827,G52828,G52829,G52830,G52831,G52832,G52833,G52834,G52835,G52836,G52837,G52838,G52839,G52840,
       G52841,G52842,G52843,G52844,G52845,G52846,G52847,G52848,G52849,G52850,G52851,G52852,G52853,G52854,G52855,G52856,G52857,G52858,G52859,G52860,
       G52861,G52862,G52863,G52864,G52865,G52866,G52867,G52868,G52869,G52870,G52871,G52872,G52873,G52874,G52875,G52876,G52877,G52878,G52879,G52880,
       G52881,G52882,G52883,G52884,G52885,G52886,G52887,G52888,G52889,G52890,G52891,G52892,G52893,G52894,G52895,G52896,G52897,G52898,G52899,G52900,
       G52901,G52902,G52903,G52904,G52905,G52906,G52907,G52908,G52909,G52910,G52911,G52912,G52913,G52914,G52915,G52916,G52917,G52918,G52919,G52920,
       G52921,G52922,G52923,G52924,G52925,G52926,G52927,G52928,G52929,G52930,G52931,G52932,G52933,G52934,G52935,G52936,G52937,G52938,G52939,G52940,
       G52941,G52942,G52943,G52944,G52945,G52946,G52947,G52948,G52949,G52950,G52951,G52952,G52953,G52954,G52955,G52956,G52957,G52958,G52959,G52960,
       G52961,G52962,G52963,G52964,G52965,G52966,G52967,G52968,G52969,G52970,G52971,G52972,G52973,G52974,G52975,G52976,G52977,G52978,G52979,G52980,
       G52981,G52982,G52983,G52984,G52985,G52986,G52987,G52988,G52989,G52990,G52991,G52992,G52993,G52994,G52995,G52996,G52997,G52998,G52999,G53000,
       G53001,G53002,G53003,G53004,G53005,G53006,G53007,G53008,G53009,G53010,G53011,G53012,G53013,G53014,G53015,G53016,G53017,G53018,G53019,G53020,
       G53021,G53022,G53023,G53024,G53025,G53026,G53027,G53028,G53029,G53030,G53031,G53032,G53033,G53034,G53035,G53036,G53037,G53038,G53039,G53040,
       G53041,G53042,G53043,G53044,G53045,G53046,G53047,G53048,G53049,G53050,G53051,G53052,G53053,G53054,G53055,G53056,G53057,G53058,G53059,G53060,
       G53061,G53062,G53063,G53064,G53065,G53066,G53067,G53068,G53069,G53070,G53071,G53072,G53073,G53074,G53075,G53076,G53077,G53078,G53079,G53080,
       G53081,G53082,G53083,G53084,G53085,G53086,G53087,G53088,G53089,G53090,G53091,G53092,G53093,G53094,G53095,G53096,G53097,G53098,G53099,G53100,
       G53101,G53102,G53103,G53104,G53105,G53106,G53107,G53108,G53109,G53110,G53111,G53112,G53113,G53114,G53115,G53116,G53117,G53118,G53119,G53120,
       G53121,G53122,G53123,G53124,G53125,G53126,G53127,G53128,G53129,G53130,G53131,G53132,G53133,G53134,G53135,G53136,G53137,G53138,G53139,G53140,
       G53141,G53142,G53143,G53144,G53145,G53146,G53147,G53148,G53149,G53150,G53151,G53152,G53153,G53154,G53155,G53156,G53157,G53158,G53159,G53160,
       G53161,G53162,G53163,G53164,G53165,G53166,G53167,G53168,G53169,G53170,G53171,G53172,G53173,G53174,G53175,G53176,G53177,G53178,G53179,G53180,
       G53181,G53182,G53183,G53184,G53185,G53186,G53187,G53188,G53189,G53190,G53191,G53192,G53193,G53194,G53195,G53196,G53197,G53198,G53199,G53200,
       G53201,G53202,G53203,G53204,G53205,G53206,G53207,G53208,G53209,G53210,G53211,G53212,G53213,G53214,G53215,G53216,G53217,G53218,G53219,G53220,
       G53221,G53222,G53223,G53224,G53225,G53226,G53227,G53228,G53229,G53230,G53231,G53232,G53233,G53234,G53235,G53236,G53237,G53238,G53239,G53240,
       G53241,G53242,G53243,G53244,G53245,G53246,G53247,G53248,G53249,G53250,G53251,G53252,G53253,G53254,G53255,G53256,G53257,G53258,G53259,G53260,
       G53261,G53262,G53263,G53264,G53265,G53266,G53267,G53268,G53269,G53270,G53271,G53272,G53273,G53274,G53275,G53276,G53277,G53278,G53279,G53280,
       G53281,G53282,G53283,G53284,G53285,G53286,G53287,G53288,G53289,G53290,G53291,G53292,G53293,G53294,G53295,G53296,G53297,G53298,G53299,G53300,
       G53301,G53302,G53303,G53304,G53305,G53306,G53307,G53308,G53309,G53310,G53311,G53312,G53313,G53314,G53315,G53316,G53317,G53318,G53319,G53320,
       G53321,G53322,G53323,G53324,G53325,G53326,G53327,G53328,G53329,G53330,G53331,G53332,G53333,G53334,G53335,G53336,G53337,G53338,G53339,G53340,
       G53341,G53342,G53343,G53344,G53345,G53346,G53347,G53348,G53349,G53350,G53351,G53352,G53353,G53354,G53355,G53356,G53357,G53358,G53359,G53360,
       G53361,G53362,G53363,G53364,G53365,G53366,G53367,G53368,G53369,G53370,G53371,G53372,G53373,G53374,G53375,G53376,G53377,G53378,G53379,G53380,
       G53381,G53382,G53383,G53384,G53385,G53386,G53387,G53388,G53389,G53390,G53391,G53392,G53393,G53394,G53395,G53396,G53397,G53398,G53399,G53400,
       G53401,G53402,G53403,G53404,G53405,G53406,G53407,G53408,G53409,G53410,G53411,G53412,G53413,G53414,G53415,G53416,G53417,G53418,G53419,G53420,
       G53421,G53422,G53423,G53424,G53425,G53426,G53427,G53428,G53429,G53430,G53431,G53432,G53433,G53434,G53435,G53436,G53437,G53438,G53439,G53440,
       G53441,G53442,G53443,G53444,G53445,G53446,G53447,G53448,G53449,G53450,G53451,G53452,G53453,G53454,G53455,G53456,G53457,G53458,G53459,G53460,
       G53461,G53462,G53463,G53464,G53465,G53466,G53467,G53468,G53469,G53470,G53471,G53472,G53473,G53474,G53475,G53476,G53477,G53478,G53479,G53480,
       G53481,G53482,G53483,G53484,G53485,G53486,G53487,G53488,G53489,G53490,G53491,G53492,G53493,G53494,G53495,G53496,G53497,G53498,G53499,G53500,
       G53501,G53502,G53503,G53504,G53505,G53506,G53507,G53508,G53509,G53510,G53511,G53512,G53513,G53514,G53515,G53516,G53517,G53518,G53519,G53520,
       G53521,G53522,G53523,G53524,G53525,G53526,G53527,G53528,G53529,G53530,G53531,G53532,G53533,G53534,G53535,G53536,G53537,G53538,G53539,G53540,
       G53541,G53542,G53543,G53544,G53545,G53546,G53547,G53548,G53549,G53550,G53551,G53552,G53553,G53554,G53555,G53556,G53557,G53558,G53559,G53560,
       G53561,G53562,G53563,G53564,G53565,G53566,G53567,G53568,G53569,G53570,G53571,G53572,G53573,G53574,G53575,G53576,G53577,G53578,G53579,G53580,
       G53581,G53582,G53583,G53584,G53585,G53586,G53587,G53588,G53589,G53590,G53591,G53592,G53593,G53594,G53595,G53596,G53597,G53598,G53599,G53600,
       G53601,G53602,G53603,G53604,G53605,G53606,G53607,G53608,G53609,G53610,G53611,G53612,G53613,G53614,G53615,G53616,G53617,G53618,G53619,G53620,
       G53621,G53622,G53623,G53624,G53625,G53626,G53627,G53628,G53629,G53630,G53631,G53632,G53633,G53634,G53635,G53636,G53637,G53638,G53639,G53640,
       G53641,G53642,G53643,G53644,G53645,G53646,G53647,G53648,G53649,G53650,G53651,G53652,G53653,G53654,G53655,G53656,G53657,G53658,G53659,G53660,
       G53661,G53662,G53663,G53664,G53665,G53666,G53667,G53668,G53669,G53670,G53671,G53672,G53673,G53674,G53675,G53676,G53677,G53678,G53679,G53680,
       G53681,G53682,G53683,G53684,G53685,G53686,G53687,G53688,G53689,G53690,G53691,G53692,G53693,G53694,G53695,G53696,G53697,G53698,G53699,G53700,
       G53701,G53702,G53703,G53704,G53705,G53706,G53707,G53708,G53709,G53710,G53711,G53712,G53713,G53714,G53715,G53716,G53717,G53718,G53719,G53720,
       G53721,G53722,G53723,G53724,G53725,G53726,G53727,G53728,G53729,G53730,G53731,G53732,G53733,G53734,G53735,G53736,G53737,G53738,G53739,G53740,
       G53741,G53742,G53743,G53744,G53745,G53746,G53747,G53748,G53749,G53750,G53751,G53752,G53753,G53754,G53755,G53756,G53757,G53758,G53759,G53760,
       G53761,G53762,G53763,G53764,G53765,G53766,G53767,G53768,G53769,G53770,G53771,G53772,G53773,G53774,G53775,G53776,G53777,G53778,G53779,G53780,
       G53781,G53782,G53783,G53784,G53785,G53786,G53787,G53788,G53789,G53790,G53791,G53792,G53793,G53794,G53795,G53796,G53797,G53798,G53799,G53800,
       G53801,G53802,G53803,G53804,G53805,G53806,G53807,G53808,G53809,G53810,G53811,G53812,G53813,G53814,G53815,G53816,G53817,G53818,G53819,G53820,
       G53821,G53822,G53823,G53824,G53825,G53826,G53827,G53828,G53829,G53830,G53831,G53832,G53833,G53834,G53835,G53836,G53837,G53838,G53839,G53840,
       G53841,G53842,G53843,G53844,G53845,G53846,G53847,G53848,G53849,G53850,G53851,G53852,G53853,G53854,G53855,G53856,G53857,G53858,G53859,G53860,
       G53861,G53862,G53863,G53864,G53865,G53866,G53867,G53868,G53869,G53870,G53871,G53872,G53873,G53874,G53875,G53876,G53877,G53878,G53879,G53880,
       G53881,G53882,G53883,G53884,G53885,G53886,G53887,G53888,G53889,G53890,G53891,G53892,G53893,G53894,G53895,G53896,G53897,G53898,G53899,G53900,
       G53901,G53902,G53903,G53904,G53905,G53906,G53907,G53908,G53909,G53910,G53911,G53912,G53913,G53914,G53915,G53916,G53917,G53918,G53919,G53920,
       G53921,G53922,G53923,G53924,G53925,G53926,G53927,G53928,G53929,G53930,G53931,G53932,G53933,G53934,G53935,G53936,G53937,G53938,G53939,G53940,
       G53941,G53942,G53943,G53944,G53945,G53946,G53947,G53948,G53949,G53950,G53951,G53952,G53953,G53954,G53955,G53956,G53957,G53958,G53959,G53960,
       G53961,G53962,G53963,G53964,G53965,G53966,G53967,G53968,G53969,G53970,G53971,G53972,G53973,G53974,G53975,G53976,G53977,G53978,G53979,G53980,
       G53981,G53982,G53983,G53984,G53985,G53986,G53987,G53988,G53989,G53990,G53991,G53992,G53993,G53994,G53995,G53996,G53997,G53998,G53999,G54000,
       G54001,G54002,G54003,G54004,G54005,G54006,G54007,G54008,G54009,G54010,G54011,G54012,G54013,G54014,G54015,G54016,G54017,G54018,G54019,G54020,
       G54021,G54022,G54023,G54024,G54025,G54026,G54027,G54028,G54029,G54030,G54031,G54032,G54033,G54034,G54035,G54036,G54037,G54038,G54039,G54040,
       G54041,G54042,G54043,G54044,G54045,G54046,G54047,G54048,G54049,G54050,G54051,G54052,G54053,G54054,G54055,G54056,G54057,G54058,G54059,G54060,
       G54061,G54062,G54063,G54064,G54065,G54066,G54067,G54068,G54069,G54070,G54071,G54072,G54073,G54074,G54075,G54076,G54077,G54078,G54079,G54080,
       G54081,G54082,G54083,G54084,G54085,G54086,G54087,G54088,G54089,G54090,G54091,G54092,G54093,G54094,G54095,G54096,G54097,G54098,G54099,G54100,
       G54101,G54102,G54103,G54104,G54105,G54106,G54107,G54108,G54109,G54110,G54111,G54112,G54113,G54114,G54115,G54116,G54117,G54118,G54119,G54120,
       G54121,G54122,G54123,G54124,G54125,G54126,G54127,G54128,G54129,G54130,G54131,G54132,G54133,G54134,G54135,G54136,G54137,G54138,G54139,G54140,
       G54141,G54142,G54143,G54144,G54145,G54146,G54147,G54148,G54149,G54150,G54151,G54152,G54153,G54154,G54155,G54156,G54157,G54158,G54159,G54160,
       G54161,G54162,G54163,G54164,G54165,G54166,G54167,G54168,G54169,G54170,G54171,G54172,G54173,G54174,G54175,G54176,G54177,G54178,G54179,G54180,
       G54181,G54182,G54183,G54184,G54185,G54186,G54187,G54188,G54189,G54190,G54191,G54192,G54193,G54194,G54195,G54196,G54197,G54198,G54199,G54200,
       G54201,G54202,G54203,G54204,G54205,G54206,G54207,G54208,G54209,G54210,G54211,G54212,G54213,G54214,G54215,G54216,G54217,G54218,G54219,G54220,
       G54221,G54222,G54223,G54224,G54225,G54226,G54227,G54228,G54229,G54230,G54231,G54232,G54233,G54234,G54235,G54236,G54237,G54238,G54239,G54240,
       G54241,G54242,G54243,G54244,G54245,G54246,G54247,G54248,G54249,G54250,G54251,G54252,G54253,G54254,G54255,G54256,G54257,G54258,G54259,G54260,
       G54261,G54262,G54263,G54264,G54265,G54266,G54267,G54268,G54269,G54270,G54271,G54272,G54273,G54274,G54275,G54276,G54277,G54278,G54279,G54280,
       G54281,G54282,G54283,G54284,G54285,G54286,G54287,G54288,G54289,G54290,G54291,G54292,G54293,G54294,G54295,G54296,G54297,G54298,G54299,G54300,
       G54301,G54302,G54303,G54304,G54305,G54306,G54307,G54308,G54309,G54310,G54311,G54312,G54313,G54314,G54315,G54316,G54317,G54318,G54319,G54320,
       G54321,G54322,G54323,G54324,G54325,G54326,G54327,G54328,G54329,G54330,G54331,G54332,G54333,G54334,G54335,G54336,G54337,G54338,G54339,G54340,
       G54341,G54342,G54343,G54344,G54345,G54346,G54347,G54348,G54349,G54350,G54351,G54352,G54353,G54354,G54355,G54356,G54357,G54358,G54359,G54360,
       G54361,G54362,G54363,G54364,G54365,G54366,G54367,G54368,G54369,G54370,G54371,G54372,G54373,G54374,G54375,G54376,G54377,G54378,G54379,G54380,
       G54381,G54382,G54383,G54384,G54385,G54386,G54387,G54388,G54389,G54390,G54391,G54392,G54393,G54394,G54395,G54396,G54397,G54398,G54399,G54400,
       G54401,G54402,G54403,G54404,G54405,G54406,G54407,G54408,G54409,G54410,G54411,G54412,G54413,G54414,G54415,G54416,G54417,G54418,G54419,G54420,
       G54421,G54422,G54423,G54424,G54425,G54426,G54427,G54428,G54429,G54430,G54431,G54432,G54433,G54434,G54435,G54436,G54437,G54438,G54439,G54440,
       G54441,G54442,G54443,G54444,G54445,G54446,G54447,G54448,G54449,G54450,G54451,G54452,G54453,G54454,G54455,G54456,G54457,G54458,G54459,G54460,
       G54461,G54462,G54463,G54464,G54465,G54466,G54467,G54468,G54469,G54470,G54471,G54472,G54473,G54474,G54475,G54476,G54477,G54478,G54479,G54480,
       G54481,G54482,G54483,G54484,G54485,G54486,G54487,G54488,G54489,G54490,G54491,G54492,G54493,G54494,G54495,G54496,G54497,G54498,G54499,G54500,
       G54501,G54502,G54503,G54504,G54505,G54506,G54507,G54508,G54509,G54510,G54511,G54512,G54513,G54514,G54515,G54516,G54517,G54518,G54519,G54520,
       G54521,G54522,G54523,G54524,G54525,G54526,G54527,G54528,G54529,G54530,G54531,G54532,G54533,G54534,G54535,G54536,G54537,G54538,G54539,G54540,
       G54541,G54542,G54543,G54544,G54545,G54546,G54547,G54548,G54549,G54550,G54551,G54552,G54553,G54554,G54555,G54556,G54557,G54558,G54559,G54560,
       G54561,G54562,G54563,G54564,G54565,G54566,G54567,G54568,G54569,G54570,G54571,G54572,G54573,G54574,G54575,G54576,G54577,G54578,G54579,G54580,
       G54581,G54582,G54583,G54584,G54585,G54586,G54587,G54588,G54589,G54590,G54591,G54592,G54593,G54594,G54595,G54596,G54597,G54598,G54599,G54600,
       G54601,G54602,G54603,G54604,G54605,G54606,G54607,G54608,G54609,G54610,G54611,G54612,G54613,G54614,G54615,G54616,G54617,G54618,G54619,G54620,
       G54621,G54622,G54623,G54624,G54625,G54626,G54627,G54628,G54629,G54630,G54631,G54632,G54633,G54634,G54635,G54636,G54637,G54638,G54639,G54640,
       G54641,G54642,G54643,G54644,G54645,G54646,G54647,G54648,G54649,G54650,G54651,G54652,G54653,G54654,G54655,G54656,G54657,G54658,G54659,G54660,
       G54661,G54662,G54663,G54664,G54665,G54666,G54667,G54668,G54669,G54670,G54671,G54672,G54673,G54674,G54675,G54676,G54677,G54678,G54679,G54680,
       G54681,G54682,G54683,G54684,G54685,G54686,G54687,G54688,G54689,G54690,G54691,G54692,G54693,G54694,G54695,G54696,G54697,G54698,G54699,G54700,
       G54701,G54702,G54703,G54704,G54705,G54706,G54707,G54708,G54709,G54710,G54711,G54712,G54713,G54714,G54715,G54716,G54717,G54718,G54719,G54720,
       G54721,G54722,G54723,G54724,G54725,G54726,G54727,G54728,G54729,G54730,G54731,G54732,G54733,G54734,G54735,G54736,G54737,G54738,G54739,G54740,
       G54741,G54742,G54743,G54744,G54745,G54746,G54747,G54748,G54749,G54750,G54751,G54752,G54753,G54754,G54755,G54756,G54757,G54758,G54759,G54760,
       G54761,G54762,G54763,G54764,G54765,G54766,G54767,G54768,G54769,G54770,G54771,G54772,G54773,G54774,G54775,G54776,G54777,G54778,G54779,G54780,
       G54781,G54782,G54783,G54784,G54785,G54786,G54787,G54788,G54789,G54790,G54791,G54792,G54793,G54794,G54795,G54796,G54797,G54798,G54799,G54800,
       G54801,G54802,G54803,G54804,G54805,G54806,G54807,G54808,G54809,G54810,G54811,G54812,G54813,G54814,G54815,G54816,G54817,G54818,G54819,G54820,
       G54821,G54822,G54823,G54824,G54825,G54826,G54827,G54828,G54829,G54830,G54831,G54832,G54833,G54834,G54835,G54836,G54837,G54838,G54839,G54840,
       G54841,G54842,G54843,G54844,G54845,G54846,G54847,G54848,G54849,G54850,G54851,G54852,G54853,G54854,G54855,G54856,G54857,G54858,G54859,G54860,
       G54861,G54862,G54863,G54864,G54865,G54866,G54867,G54868,G54869,G54870,G54871,G54872,G54873,G54874,G54875,G54876,G54877,G54878,G54879,G54880,
       G54881,G54882,G54883,G54884,G54885,G54886,G54887,G54888,G54889,G54890,G54891,G54892,G54893,G54894,G54895,G54896,G54897,G54898,G54899,G54900,
       G54901,G54902,G54903,G54904,G54905,G54906,G54907,G54908,G54909,G54910,G54911,G54912,G54913,G54914,G54915,G54916,G54917,G54918,G54919,G54920,
       G54921,G54922,G54923,G54924,G54925,G54926,G54927,G54928,G54929,G54930,G54931,G54932,G54933,G54934,G54935,G54936,G54937,G54938,G54939,G54940,
       G54941,G54942,G54943,G54944,G54945,G54946,G54947,G54948,G54949,G54950,G54951,G54952,G54953,G54954,G54955,G54956,G54957,G54958,G54959,G54960,
       G54961,G54962,G54963,G54964,G54965,G54966,G54967,G54968,G54969,G54970,G54971,G54972,G54973,G54974,G54975,G54976,G54977,G54978,G54979,G54980,
       G54981,G54982,G54983,G54984,G54985,G54986,G54987,G54988,G54989,G54990,G54991,G54992,G54993,G54994,G54995,G54996,G54997,G54998,G54999,G55000,
       G55001,G55002,G55003,G55004,G55005,G55006,G55007,G55008,G55009,G55010,G55011,G55012,G55013,G55014,G55015,G55016,G55017,G55018,G55019,G55020,
       G55021,G55022,G55023,G55024,G55025,G55026,G55027,G55028,G55029,G55030,G55031,G55032,G55033,G55034,G55035,G55036,G55037,G55038,G55039,G55040,
       G55041,G55042,G55043,G55044,G55045,G55046,G55047,G55048,G55049,G55050,G55051,G55052,G55053,G55054,G55055,G55056,G55057,G55058,G55059,G55060,
       G55061,G55062,G55063,G55064,G55065,G55066,G55067,G55068,G55069,G55070,G55071,G55072,G55073,G55074,G55075,G55076,G55077,G55078,G55079,G55080,
       G55081,G55082,G55083,G55084,G55085,G55086,G55087,G55088,G55089,G55090,G55091,G55092,G55093,G55094,G55095,G55096,G55097,G55098,G55099,G55100,
       G55101,G55102,G55103,G55104,G55105,G55106,G55107,G55108,G55109,G55110,G55111,G55112,G55113,G55114,G55115,G55116,G55117,G55118,G55119,G55120,
       G55121,G55122,G55123,G55124,G55125,G55126,G55127,G55128,G55129,G55130,G55131,G55132,G55133,G55134,G55135,G55136,G55137,G55138,G55139,G55140,
       G55141,G55142,G55143,G55144,G55145,G55146,G55147,G55148,G55149,G55150,G55151,G55152,G55153,G55154,G55155,G55156,G55157,G55158,G55159,G55160,
       G55161,G55162,G55163,G55164,G55165,G55166,G55167,G55168,G55169,G55170,G55171,G55172,G55173,G55174,G55175,G55176,G55177,G55178,G55179,G55180,
       G55181,G55182,G55183,G55184,G55185,G55186,G55187,G55188,G55189,G55190,G55191,G55192,G55193,G55194,G55195,G55196,G55197,G55198,G55199,G55200,
       G55201,G55202,G55203,G55204,G55205,G55206,G55207,G55208,G55209,G55210,G55211,G55212,G55213,G55214,G55215,G55216,G55217,G55218,G55219,G55220,
       G55221,G55222,G55223,G55224,G55225,G55226,G55227,G55228,G55229,G55230,G55231,G55232,G55233,G55234,G55235,G55236,G55237,G55238,G55239,G55240,
       G55241,G55242,G55243,G55244,G55245,G55246,G55247,G55248,G55249,G55250,G55251,G55252,G55253,G55254,G55255,G55256,G55257,G55258,G55259,G55260,
       G55261,G55262,G55263,G55264,G55265,G55266,G55267,G55268,G55269,G55270,G55271,G55272,G55273,G55274,G55275,G55276,G55277,G55278,G55279,G55280,
       G55281,G55282,G55283,G55284,G55285,G55286,G55287,G55288,G55289,G55290,G55291,G55292,G55293,G55294,G55295,G55296,G55297,G55298,G55299,G55300,
       G55301,G55302,G55303,G55304,G55305,G55306,G55307,G55308,G55309,G55310,G55311,G55312,G55313,G55314,G55315,G55316,G55317,G55318,G55319,G55320,
       G55321,G55322,G55323,G55324,G55325,G55326,G55327,G55328,G55329,G55330,G55331,G55332,G55333,G55334,G55335,G55336,G55337,G55338,G55339,G55340,
       G55341,G55342,G55343,G55344,G55345,G55346,G55347,G55348,G55349,G55350,G55351,G55352,G55353,G55354,G55355,G55356,G55357,G55358,G55359,G55360,
       G55361,G55362,G55363,G55364,G55365,G55366,G55367,G55368,G55369,G55370,G55371,G55372,G55373,G55374,G55375,G55376,G55377,G55378,G55379,G55380,
       G55381,G55382,G55383,G55384,G55385,G55386,G55387,G55388,G55389,G55390,G55391,G55392,G55393,G55394,G55395,G55396,G55397,G55398,G55399,G55400,
       G55401,G55402,G55403,G55404,G55405,G55406,G55407,G55408,G55409,G55410,G55411,G55412,G55413,G55414,G55415,G55416,G55417,G55418,G55419,G55420,
       G55421,G55422,G55423,G55424,G55425,G55426,G55427,G55428,G55429,G55430,G55431,G55432,G55433,G55434,G55435,G55436,G55437,G55438,G55439,G55440,
       G55441,G55442,G55443,G55444,G55445,G55446,G55447,G55448,G55449,G55450,G55451,G55452,G55453,G55454,G55455,G55456,G55457,G55458,G55459,G55460,
       G55461,G55462,G55463,G55464,G55465,G55466,G55467,G55468,G55469,G55470,G55471,G55472,G55473,G55474,G55475,G55476,G55477,G55478,G55479,G55480,
       G55481,G55482,G55483,G55484,G55485,G55486,G55487,G55488,G55489,G55490,G55491,G55492,G55493,G55494,G55495,G55496,G55497,G55498,G55499,G55500,
       G55501,G55502,G55503,G55504,G55505,G55506,G55507,G55508,G55509,G55510,G55511,G55512,G55513,G55514,G55515,G55516,G55517,G55518,G55519,G55520,
       G55521,G55522,G55523,G55524,G55525,G55526,G55527,G55528,G55529,G55530,G55531,G55532,G55533,G55534,G55535,G55536,G55537,G55538,G55539,G55540,
       G55541,G55542,G55543,G55544,G55545,G55546,G55547,G55548,G55549,G55550,G55551,G55552,G55553,G55554,G55555,G55556,G55557,G55558,G55559,G55560,
       G55561,G55562,G55563,G55564,G55565,G55566,G55567,G55568,G55569,G55570,G55571,G55572,G55573,G55574,G55575,G55576,G55577,G55578,G55579,G55580,
       G55581,G55582,G55583,G55584,G55585,G55586,G55587,G55588,G55589,G55590,G55591,G55592,G55593,G55594,G55595,G55596,G55597,G55598,G55599,G55600,
       G55601,G55602,G55603,G55604,G55605,G55606,G55607,G55608,G55609,G55610,G55611,G55612,G55613,G55614,G55615,G55616,G55617,G55618,G55619,G55620,
       G55621,G55622,G55623,G55624,G55625,G55626,G55627,G55628,G55629,G55630,G55631,G55632,G55633,G55634,G55635,G55636,G55637,G55638,G55639,G55640,
       G55641,G55642,G55643,G55644,G55645,G55646,G55647,G55648,G55649,G55650,G55651,G55652,G55653,G55654,G55655,G55656,G55657,G55658,G55659,G55660,
       G55661,G55662,G55663,G55664,G55665,G55666,G55667,G55668,G55669,G55670,G55671,G55672,G55673,G55674,G55675,G55676,G55677,G55678,G55679,G55680,
       G55681,G55682,G55683,G55684,G55685,G55686,G55687,G55688,G55689,G55690,G55691,G55692,G55693,G55694,G55695,G55696,G55697,G55698,G55699,G55700,
       G55701,G55702,G55703,G55704,G55705,G55706,G55707,G55708,G55709,G55710,G55711,G55712,G55713,G55714,G55715,G55716,G55717,G55718,G55719,G55720,
       G55721,G55722,G55723,G55724,G55725,G55726,G55727,G55728,G55729,G55730,G55731,G55732,G55733,G55734,G55735,G55736,G55737,G55738,G55739,G55740,
       G55741,G55742,G55743,G55744,G55745,G55746,G55747,G55748,G55749,G55750,G55751,G55752,G55753,G55754,G55755,G55756,G55757,G55758,G55759,G55760,
       G55761,G55762,G55763,G55764,G55765,G55766,G55767,G55768,G55769,G55770,G55771,G55772,G55773,G55774,G55775,G55776,G55777,G55778,G55779,G55780,
       G55781,G55782,G55783,G55784,G55785,G55786,G55787,G55788,G55789,G55790,G55791,G55792,G55793,G55794,G55795,G55796,G55797,G55798,G55799,G55800,
       G55801,G55802,G55803,G55804,G55805,G55806,G55807,G55808,G55809,G55810,G55811,G55812,G55813,G55814,G55815,G55816,G55817,G55818,G55819,G55820,
       G55821,G55822,G55823,G55824,G55825,G55826,G55827,G55828,G55829,G55830,G55831,G55832,G55833,G55834,G55835,G55836,G55837,G55838,G55839,G55840,
       G55841,G55842,G55843,G55844,G55845,G55846,G55847,G55848,G55849,G55850,G55851,G55852,G55853,G55854,G55855,G55856,G55857,G55858,G55859,G55860,
       G55861,G55862,G55863,G55864,G55865,G55866,G55867,G55868,G55869,G55870,G55871,G55872,G55873,G55874,G55875,G55876,G55877,G55878,G55879,G55880,
       G55881,G55882,G55883,G55884,G55885,G55886,G55887,G55888,G55889,G55890,G55891,G55892,G55893,G55894,G55895,G55896,G55897,G55898,G55899,G55900,
       G55901,G55902,G55903,G55904,G55905,G55906,G55907,G55908,G55909,G55910,G55911,G55912,G55913,G55914,G55915,G55916,G55917,G55918,G55919,G55920,
       G55921,G55922,G55923,G55924,G55925,G55926,G55927,G55928,G55929,G55930,G55931,G55932,G55933,G55934,G55935,G55936,G55937,G55938,G55939,G55940,
       G55941,G55942,G55943,G55944,G55945,G55946,G55947,G55948,G55949,G55950,G55951,G55952,G55953,G55954,G55955,G55956,G55957,G55958,G55959,G55960,
       G55961,G55962,G55963,G55964,G55965,G55966,G55967,G55968,G55969,G55970,G55971,G55972,G55973,G55974,G55975,G55976,G55977,G55978,G55979,G55980,
       G55981,G55982,G55983,G55984,G55985,G55986,G55987,G55988,G55989,G55990,G55991,G55992,G55993,G55994,G55995,G55996,G55997,G55998,G55999,G56000,
       G56001,G56002,G56003,G56004,G56005,G56006,G56007,G56008,G56009,G56010,G56011,G56012,G56013,G56014,G56015,G56016,G56017,G56018,G56019,G56020,
       G56021,G56022,G56023,G56024,G56025,G56026,G56027,G56028,G56029,G56030,G56031,G56032,G56033,G56034,G56035,G56036,G56037,G56038,G56039,G56040,
       G56041,G56042,G56043,G56044,G56045,G56046,G56047,G56048,G56049,G56050,G56051,G56052,G56053,G56054,G56055,G56056,G56057,G56058,G56059,G56060,
       G56061,G56062,G56063,G56064,G56065,G56066,G56067,G56068,G56069,G56070,G56071,G56072,G56073,G56074,G56075,G56076,G56077,G56078,G56079,G56080,
       G56081,G56082,G56083,G56084,G56085,G56086,G56087,G56088,G56089,G56090,G56091,G56092,G56093,G56094,G56095,G56096,G56097,G56098,G56099,G56100,
       G56101,G56102,G56103,G56104,G56105,G56106,G56107,G56108,G56109,G56110,G56111,G56112,G56113,G56114,G56115,G56116,G56117,G56118,G56119,G56120,
       G56121,G56122,G56123,G56124,G56125,G56126,G56127,G56128,G56129,G56130,G56131,G56132,G56133,G56134,G56135,G56136,G56137,G56138,G56139,G56140,
       G56141,G56142,G56143,G56144,G56145,G56146,G56147,G56148,G56149,G56150,G56151,G56152,G56153,G56154,G56155,G56156,G56157,G56158,G56159,G56160,
       G56161,G56162,G56163,G56164,G56165,G56166,G56167,G56168,G56169,G56170,G56171,G56172,G56173,G56174,G56175,G56176,G56177,G56178,G56179,G56180,
       G56181,G56182,G56183,G56184,G56185,G56186,G56187,G56188,G56189,G56190,G56191,G56192,G56193,G56194,G56195,G56196,G56197,G56198,G56199,G56200,
       G56201,G56202,G56203,G56204,G56205,G56206,G56207,G56208,G56209,G56210,G56211,G56212,G56213,G56214,G56215,G56216,G56217,G56218,G56219,G56220,
       G56221,G56222,G56223,G56224,G56225,G56226,G56227,G56228,G56229,G56230,G56231,G56232,G56233,G56234,G56235,G56236,G56237,G56238,G56239,G56240,
       G56241,G56242,G56243,G56244,G56245,G56246,G56247,G56248,G56249,G56250,G56251,G56252,G56253,G56254,G56255,G56256,G56257,G56258,G56259,G56260,
       G56261,G56262,G56263,G56264,G56265,G56266,G56267,G56268,G56269,G56270,G56271,G56272,G56273,G56274,G56275,G56276,G56277,G56278,G56279,G56280,
       G56281,G56282,G56283,G56284,G56285,G56286,G56287,G56288,G56289,G56290,G56291,G56292,G56293,G56294,G56295,G56296,G56297,G56298,G56299,G56300,
       G56301,G56302,G56303,G56304,G56305,G56306,G56307,G56308,G56309,G56310,G56311,G56312,G56313,G56314,G56315,G56316,G56317,G56318,G56319,G56320,
       G56321,G56322,G56323,G56324,G56325,G56326,G56327,G56328,G56329,G56330,G56331,G56332,G56333,G56334,G56335,G56336,G56337,G56338,G56339,G56340,
       G56341,G56342,G56343,G56344,G56345,G56346,G56347,G56348,G56349,G56350,G56351,G56352,G56353,G56354,G56355,G56356,G56357,G56358,G56359,G56360,
       G56361,G56362,G56363,G56364,G56365,G56366,G56367,G56368,G56369,G56370,G56371,G56372,G56373,G56374,G56375,G56376,G56377,G56378,G56379,G56380,
       G56381,G56382,G56383,G56384,G56385,G56386,G56387,G56388,G56389,G56390,G56391,G56392,G56393,G56394,G56395,G56396,G56397,G56398,G56399,G56400,
       G56401,G56402,G56403,G56404,G56405,G56406,G56407,G56408,G56409,G56410,G56411,G56412,G56413,G56414,G56415,G56416,G56417,G56418,G56419,G56420,
       G56421,G56422,G56423,G56424,G56425,G56426,G56427,G56428,G56429,G56430,G56431,G56432,G56433,G56434,G56435,G56436,G56437,G56438,G56439,G56440,
       G56441,G56442,G56443,G56444,G56445,G56446,G56447,G56448,G56449,G56450,G56451,G56452,G56453,G56454,G56455,G56456,G56457,G56458,G56459,G56460,
       G56461,G56462,G56463,G56464,G56465,G56466,G56467,G56468,G56469,G56470,G56471,G56472,G56473,G56474,G56475,G56476,G56477,G56478,G56479,G56480,
       G56481,G56482,G56483,G56484,G56485,G56486,G56487,G56488,G56489,G56490,G56491,G56492,G56493,G56494,G56495,G56496,G56497,G56498,G56499,G56500,
       G56501,G56502,G56503,G56504,G56505,G56506,G56507,G56508,G56509,G56510,G56511,G56512,G56513,G56514,G56515,G56516,G56517,G56518,G56519,G56520,
       G56521,G56522,G56523,G56524,G56525,G56526,G56527,G56528,G56529,G56530,G56531,G56532,G56533,G56534,G56535,G56536,G56537,G56538,G56539,G56540,
       G56541,G56542,G56543,G56544,G56545,G56546,G56547,G56548,G56549,G56550,G56551,G56552,G56553,G56554,G56555,G56556,G56557,G56558,G56559,G56560,
       G56561,G56562,G56563,G56564,G56565,G56566,G56567,G56568,G56569,G56570,G56571,G56572,G56573,G56574,G56575,G56576,G56577,G56578,G56579,G56580,
       G56581,G56582,G56583,G56584,G56585,G56586,G56587,G56588,G56589,G56590,G56591,G56592,G56593,G56594,G56595,G56596,G56597,G56598,G56599,G56600,
       G56601,G56602,G56603,G56604,G56605,G56606,G56607,G56608,G56609,G56610,G56611,G56612,G56613,G56614,G56615,G56616,G56617,G56618,G56619,G56620,
       G56621,G56622,G56623,G56624,G56625,G56626,G56627,G56628,G56629,G56630,G56631,G56632,G56633,G56634,G56635,G56636,G56637,G56638,G56639,G56640,
       G56641,G56642,G56643,G56644,G56645,G56646,G56647,G56648,G56649,G56650,G56651,G56652,G56653,G56654,G56655,G56656,G56657,G56658,G56659,G56660,
       G56661,G56662,G56663,G56664,G56665,G56666,G56667,G56668,G56669,G56670,G56671,G56672,G56673,G56674,G56675,G56676,G56677,G56678,G56679,G56680,
       G56681,G56682,G56683,G56684,G56685,G56686,G56687,G56688,G56689,G56690,G56691,G56692,G56693,G56694,G56695,G56696,G56697,G56698,G56699,G56700,
       G56701,G56702,G56703,G56704,G56705,G56706,G56707,G56708,G56709,G56710,G56711,G56712,G56713,G56714,G56715,G56716,G56717,G56718,G56719,G56720,
       G56721,G56722,G56723,G56724,G56725,G56726,G56727,G56728,G56729,G56730,G56731,G56732,G56733,G56734,G56735,G56736,G56737,G56738,G56739,G56740,
       G56741,G56742,G56743,G56744,G56745,G56746,G56747,G56748,G56749,G56750,G56751,G56752,G56753,G56754,G56755,G56756,G56757,G56758,G56759,G56760,
       G56761,G56762,G56763,G56764,G56765,G56766,G56767,G56768,G56769,G56770,G56771,G56772,G56773,G56774,G56775,G56776,G56777,G56778,G56779,G56780,
       G56781,G56782,G56783,G56784,G56785,G56786,G56787,G56788,G56789,G56790,G56791,G56792,G56793,G56794,G56795,G56796,G56797,G56798,G56799,G56800,
       G56801,G56802,G56803,G56804,G56805,G56806,G56807,G56808,G56809,G56810,G56811,G56812,G56813,G56814,G56815,G56816,G56817,G56818,G56819,G56820,
       G56821,G56822,G56823,G56824,G56825,G56826,G56827,G56828,G56829,G56830,G56831,G56832,G56833,G56834,G56835,G56836,G56837,G56838,G56839,G56840,
       G56841,G56842,G56843,G56844,G56845,G56846,G56847,G56848,G56849,G56850,G56851,G56852,G56853,G56854,G56855,G56856,G56857,G56858,G56859,G56860,
       G56861,G56862,G56863,G56864,G56865,G56866,G56867,G56868,G56869,G56870,G56871,G56872,G56873,G56874,G56875,G56876,G56877,G56878,G56879,G56880,
       G56881,G56882,G56883,G56884,G56885,G56886,G56887,G56888,G56889,G56890,G56891,G56892,G56893,G56894,G56895,G56896,G56897,G56898,G56899,G56900,
       G56901,G56902,G56903,G56904,G56905,G56906,G56907,G56908,G56909,G56910,G56911,G56912,G56913,G56914,G56915,G56916,G56917,G56918,G56919,G56920,
       G56921,G56922,G56923,G56924,G56925,G56926,G56927,G56928,G56929,G56930,G56931,G56932,G56933,G56934,G56935,G56936,G56937,G56938,G56939,G56940,
       G56941,G56942,G56943,G56944,G56945,G56946,G56947,G56948,G56949,G56950,G56951,G56952,G56953,G56954,G56955,G56956,G56957,G56958,G56959,G56960,
       G56961,G56962,G56963,G56964,G56965,G56966,G56967,G56968,G56969,G56970,G56971,G56972,G56973,G56974,G56975,G56976,G56977,G56978,G56979,G56980,
       G56981,G56982,G56983,G56984,G56985,G56986,G56987,G56988,G56989,G56990,G56991,G56992,G56993,G56994,G56995,G56996,G56997,G56998,G56999,G57000,
       G57001,G57002,G57003,G57004,G57005,G57006,G57007,G57008,G57009,G57010,G57011,G57012,G57013,G57014,G57015,G57016,G57017,G57018,G57019,G57020,
       G57021,G57022,G57023,G57024,G57025,G57026,G57027,G57028,G57029,G57030,G57031,G57032,G57033,G57034,G57035,G57036,G57037,G57038,G57039,G57040,
       G57041,G57042,G57043,G57044,G57045,G57046,G57047,G57048,G57049,G57050,G57051,G57052,G57053,G57054,G57055,G57056,G57057,G57058,G57059,G57060,
       G57061,G57062,G57063,G57064,G57065,G57066,G57067,G57068,G57069,G57070,G57071,G57072,G57073,G57074,G57075,G57076,G57077,G57078,G57079,G57080,
       G57081,G57082,G57083,G57084,G57085,G57086,G57087,G57088,G57089,G57090,G57091,G57092,G57093,G57094,G57095,G57096,G57097,G57098,G57099,G57100,
       G57101,G57102,G57103,G57104,G57105,G57106,G57107,G57108,G57109,G57110,G57111,G57112,G57113,G57114,G57115,G57116,G57117,G57118,G57119,G57120,
       G57121,G57122,G57123,G57124,G57125,G57126,G57127,G57128,G57129,G57130,G57131,G57132,G57133,G57134,G57135,G57136,G57137,G57138,G57139,G57140,
       G57141,G57142,G57143,G57144,G57145,G57146,G57147,G57148,G57149,G57150,G57151,G57152,G57153,G57154,G57155,G57156,G57157,G57158,G57159,G57160,
       G57161,G57162,G57163,G57164,G57165,G57166,G57167,G57168,G57169,G57170,G57171,G57172,G57173,G57174,G57175,G57176,G57177,G57178,G57179,G57180,
       G57181,G57182,G57183,G57184,G57185,G57186,G57187,G57188,G57189,G57190,G57191,G57192,G57193,G57194,G57195,G57196,G57197,G57198,G57199,G57200,
       G57201,G57202,G57203,G57204,G57205,G57206,G57207,G57208,G57209,G57210,G57211,G57212,G57213,G57214,G57215,G57216,G57217,G57218,G57219,G57220,
       G57221,G57222,G57223,G57224,G57225,G57226,G57227,G57228,G57229,G57230,G57231,G57232,G57233,G57234,G57235,G57236,G57237,G57238,G57239,G57240,
       G57241,G57242,G57243,G57244,G57245,G57246,G57247,G57248,G57249,G57250,G57251,G57252,G57253,G57254,G57255,G57256,G57257,G57258,G57259,G57260,
       G57261,G57262,G57263,G57264,G57265,G57266,G57267,G57268,G57269,G57270,G57271,G57272,G57273,G57274,G57275,G57276,G57277,G57278,G57279,G57280,
       G57281,G57282,G57283,G57284,G57285,G57286,G57287,G57288,G57289,G57290,G57291,G57292,G57293,G57294,G57295,G57296,G57297,G57298,G57299,G57300,
       G57301,G57302,G57303,G57304,G57305,G57306,G57307,G57308,G57309,G57310,G57311,G57312,G57313,G57314,G57315,G57316,G57317,G57318,G57319,G57320,
       G57321,G57322,G57323,G57324,G57325,G57326,G57327,G57328,G57329,G57330,G57331,G57332,G57333,G57334,G57335,G57336,G57337,G57338,G57339,G57340,
       G57341,G57342,G57343,G57344,G57345,G57346,G57347,G57348,G57349,G57350,G57351,G57352,G57353,G57354,G57355,G57356,G57357,G57358,G57359,G57360,
       G57361,G57362,G57363,G57364,G57365,G57366,G57367,G57368,G57369,G57370,G57371,G57372,G57373,G57374,G57375,G57376,G57377,G57378,G57379,G57380,
       G57381,G57382,G57383,G57384,G57385,G57386,G57387,G57388,G57389,G57390,G57391,G57392,G57393,G57394,G57395,G57396,G57397,G57398,G57399,G57400,
       G57401,G57402,G57403,G57404,G57405,G57406,G57407,G57408,G57409,G57410,G57411,G57412,G57413,G57414,G57415,G57416,G57417,G57418,G57419,G57420,
       G57421,G57422,G57423,G57424,G57425,G57426,G57427,G57428,G57429,G57430,G57431,G57432,G57433,G57434,G57435,G57436,G57437,G57438,G57439,G57440,
       G57441,G57442,G57443,G57444,G57445,G57446,G57447,G57448,G57449,G57450,G57451,G57452,G57453,G57454,G57455,G57456,G57457,G57458,G57459,G57460,
       G57461,G57462,G57463,G57464,G57465,G57466,G57467,G57468,G57469,G57470,G57471,G57472,G57473,G57474,G57475,G57476,G57477,G57478,G57479,G57480,
       G57481,G57482,G57483,G57484,G57485,G57486,G57487,G57488,G57489,G57490,G57491,G57492,G57493,G57494,G57495,G57496,G57497,G57498,G57499,G57500,
       G57501,G57502,G57503,G57504,G57505,G57506,G57507,G57508,G57509,G57510,G57511,G57512,G57513,G57514,G57515,G57516,G57517,G57518,G57519,G57520,
       G57521,G57522,G57523,G57524,G57525,G57526,G57527,G57528,G57529,G57530,G57531,G57532,G57533,G57534,G57535,G57536,G57537,G57538,G57539,G57540,
       G57541,G57542,G57543,G57544,G57545,G57546,G57547,G57548,G57549,G57550,G57551,G57552,G57553,G57554,G57555,G57556,G57557,G57558,G57559,G57560,
       G57561,G57562,G57563,G57564,G57565,G57566,G57567,G57568,G57569,G57570,G57571,G57572,G57573,G57574,G57575,G57576,G57577,G57578,G57579,G57580,
       G57581,G57582,G57583,G57584,G57585,G57586,G57587,G57588,G57589,G57590,G57591,G57592,G57593,G57594,G57595,G57596,G57597,G57598,G57599,G57600,
       G57601,G57602,G57603,G57604,G57605,G57606,G57607,G57608,G57609,G57610,G57611,G57612,G57613,G57614,G57615,G57616,G57617,G57618,G57619,G57620,
       G57621,G57622,G57623,G57624,G57625,G57626,G57627,G57628,G57629,G57630,G57631,G57632,G57633,G57634,G57635,G57636,G57637,G57638,G57639,G57640,
       G57641,G57642,G57643,G57644,G57645,G57646,G57647,G57648,G57649,G57650,G57651,G57652,G57653,G57654,G57655,G57656,G57657,G57658,G57659,G57660,
       G57661,G57662,G57663,G57664,G57665,G57666,G57667,G57668,G57669,G57670,G57671,G57672,G57673,G57674,G57675,G57676,G57677,G57678,G57679,G57680,
       G57681,G57682,G57683,G57684,G57685,G57686,G57687,G57688,G57689,G57690,G57691,G57692,G57693,G57694,G57695,G57696,G57697,G57698,G57699,G57700,
       G57701,G57702,G57703,G57704,G57705,G57706,G57707,G57708,G57709,G57710,G57711,G57712,G57713,G57714,G57715,G57716,G57717,G57718,G57719,G57720,
       G57721,G57722,G57723,G57724,G57725,G57726,G57727,G57728,G57729,G57730,G57731,G57732,G57733,G57734,G57735,G57736,G57737,G57738,G57739,G57740,
       G57741,G57742,G57743,G57744,G57745,G57746,G57747,G57748,G57749,G57750,G57751,G57752,G57753,G57754,G57755,G57756,G57757,G57758,G57759,G57760,
       G57761,G57762,G57763,G57764,G57765,G57766,G57767,G57768,G57769,G57770,G57771,G57772,G57773,G57774,G57775,G57776,G57777,G57778,G57779,G57780,
       G57781,G57782,G57783,G57784,G57785,G57786,G57787,G57788,G57789,G57790,G57791,G57792,G57793,G57794,G57795,G57796,G57797,G57798,G57799,G57800,
       G57801,G57802,G57803,G57804,G57805,G57806,G57807,G57808,G57809,G57810,G57811,G57812,G57813,G57814,G57815,G57816,G57817,G57818,G57819,G57820,
       G57821,G57822,G57823,G57824,G57825,G57826,G57827,G57828,G57829,G57830,G57831,G57832,G57833,G57834,G57835,G57836,G57837,G57838,G57839,G57840,
       G57841,G57842,G57843,G57844,G57845,G57846,G57847,G57848,G57849,G57850,G57851,G57852,G57853,G57854,G57855,G57856,G57857,G57858,G57859,G57860,
       G57861,G57862,G57863,G57864,G57865,G57866,G57867,G57868,G57869,G57870,G57871,G57872,G57873,G57874,G57875,G57876,G57877,G57878,G57879,G57880,
       G57881,G57882,G57883,G57884,G57885,G57886,G57887,G57888,G57889,G57890,G57891,G57892,G57893,G57894,G57895,G57896,G57897,G57898,G57899,G57900,
       G57901,G57902,G57903,G57904,G57905,G57906,G57907,G57908,G57909,G57910,G57911,G57912,G57913,G57914,G57915,G57916,G57917,G57918,G57919,G57920,
       G57921,G57922,G57923,G57924,G57925,G57926,G57927,G57928,G57929,G57930,G57931,G57932,G57933,G57934,G57935,G57936,G57937,G57938,G57939,G57940,
       G57941,G57942,G57943,G57944,G57945,G57946,G57947,G57948,G57949,G57950,G57951,G57952,G57953,G57954,G57955,G57956,G57957,G57958,G57959,G57960,
       G57961,G57962,G57963,G57964,G57965,G57966,G57967,G57968,G57969,G57970,G57971,G57972,G57973,G57974,G57975,G57976,G57977,G57978,G57979,G57980,
       G57981,G57982,G57983,G57984,G57985,G57986,G57987,G57988,G57989,G57990,G57991,G57992,G57993,G57994,G57995,G57996,G57997,G57998,G57999,G58000,
       G58001,G58002,G58003,G58004,G58005,G58006,G58007,G58008,G58009,G58010,G58011,G58012,G58013,G58014,G58015,G58016,G58017,G58018,G58019,G58020,
       G58021,G58022,G58023,G58024,G58025,G58026,G58027,G58028,G58029,G58030,G58031,G58032,G58033,G58034,G58035,G58036,G58037,G58038,G58039,G58040,
       G58041,G58042,G58043,G58044,G58045,G58046,G58047,G58048,G58049,G58050,G58051,G58052,G58053,G58054,G58055,G58056,G58057,G58058,G58059,G58060,
       G58061,G58062,G58063,G58064,G58065,G58066,G58067,G58068,G58069,G58070,G58071,G58072,G58073,G58074,G58075,G58076,G58077,G58078,G58079,G58080,
       G58081,G58082,G58083,G58084,G58085,G58086,G58087,G58088,G58089,G58090,G58091,G58092,G58093,G58094,G58095,G58096,G58097,G58098,G58099,G58100,
       G58101,G58102,G58103,G58104,G58105,G58106,G58107,G58108,G58109,G58110,G58111,G58112,G58113,G58114,G58115,G58116,G58117,G58118,G58119,G58120,
       G58121,G58122,G58123,G58124,G58125,G58126,G58127,G58128,G58129,G58130,G58131,G58132,G58133,G58134,G58135,G58136,G58137,G58138,G58139,G58140,
       G58141,G58142,G58143,G58144,G58145,G58146,G58147,G58148,G58149,G58150,G58151,G58152,G58153,G58154,G58155,G58156,G58157,G58158,G58159,G58160,
       G58161,G58162,G58163,G58164,G58165,G58166,G58167,G58168,G58169,G58170,G58171,G58172,G58173,G58174,G58175,G58176,G58177,G58178,G58179,G58180,
       G58181,G58182,G58183,G58184,G58185,G58186,G58187,G58188,G58189,G58190,G58191,G58192,G58193,G58194,G58195,G58196,G58197,G58198,G58199,G58200,
       G58201,G58202,G58203,G58204,G58205,G58206,G58207,G58208,G58209,G58210,G58211,G58212,G58213,G58214,G58215,G58216,G58217,G58218,G58219,G58220,
       G58221,G58222,G58223,G58224,G58225,G58226,G58227,G58228,G58229,G58230,G58231,G58232,G58233,G58234,G58235,G58236,G58237,G58238,G58239,G58240,
       G58241,G58242,G58243,G58244,G58245,G58246,G58247,G58248,G58249,G58250,G58251,G58252,G58253,G58254,G58255,G58256,G58257,G58258,G58259,G58260,
       G58261,G58262,G58263,G58264,G58265,G58266,G58267,G58268,G58269,G58270,G58271,G58272,G58273,G58274,G58275,G58276,G58277,G58278,G58279,G58280,
       G58281,G58282,G58283,G58284,G58285,G58286,G58287,G58288,G58289,G58290,G58291,G58292,G58293,G58294,G58295,G58296,G58297,G58298,G58299,G58300,
       G58301,G58302,G58303,G58304,G58305,G58306,G58307,G58308,G58309,G58310,G58311,G58312,G58313,G58314,G58315,G58316,G58317,G58318,G58319,G58320,
       G58321,G58322,G58323,G58324,G58325,G58326,G58327,G58328,G58329,G58330,G58331,G58332,G58333,G58334,G58335,G58336,G58337,G58338,G58339,G58340,
       G58341,G58342,G58343,G58344,G58345,G58346,G58347,G58348,G58349,G58350,G58351,G58352,G58353,G58354,G58355,G58356,G58357,G58358,G58359,G58360,
       G58361,G58362,G58363,G58364,G58365,G58366,G58367,G58368,G58369,G58370,G58371,G58372,G58373,G58374,G58375,G58376,G58377,G58378,G58379,G58380,
       G58381,G58382,G58383,G58384,G58385,G58386,G58387,G58388,G58389,G58390,G58391,G58392,G58393,G58394,G58395,G58396,G58397,G58398,G58399,G58400,
       G58401,G58402,G58403,G58404,G58405,G58406,G58407,G58408,G58409,G58410,G58411,G58412,G58413,G58414,G58415,G58416,G58417,G58418,G58419,G58420,
       G58421,G58422,G58423,G58424,G58425,G58426,G58427,G58428,G58429,G58430,G58431,G58432,G58433,G58434,G58435,G58436,G58437,G58438,G58439,G58440,
       G58441,G58442,G58443,G58444,G58445,G58446,G58447,G58448,G58449,G58450,G58451,G58452,G58453,G58454,G58455,G58456,G58457,G58458,G58459,G58460,
       G58461,G58462,G58463,G58464,G58465,G58466,G58467,G58468,G58469,G58470,G58471,G58472,G58473,G58474,G58475,G58476,G58477,G58478,G58479,G58480,
       G58481,G58482,G58483,G58484,G58485,G58486,G58487,G58488,G58489,G58490,G58491,G58492,G58493,G58494,G58495,G58496,G58497,G58498,G58499,G58500,
       G58501,G58502,G58503,G58504,G58505,G58506,G58507,G58508,G58509,G58510,G58511,G58512,G58513,G58514,G58515,G58516,G58517,G58518,G58519,G58520,
       G58521,G58522,G58523,G58524,G58525,G58526,G58527,G58528,G58529,G58530,G58531,G58532,G58533,G58534,G58535,G58536,G58537,G58538,G58539,G58540,
       G58541,G58542,G58543,G58544,G58545,G58546,G58547,G58548,G58549,G58550,G58551,G58552,G58553,G58554,G58555,G58556,G58557,G58558,G58559,G58560,
       G58561,G58562,G58563,G58564,G58565,G58566,G58567,G58568,G58569,G58570,G58571,G58572,G58573,G58574,G58575,G58576,G58577,G58578,G58579,G58580,
       G58581,G58582,G58583,G58584,G58585,G58586,G58587,G58588,G58589,G58590,G58591,G58592,G58593,G58594,G58595,G58596,G58597,G58598,G58599,G58600,
       G58601,G58602,G58603,G58604,G58605,G58606,G58607,G58608,G58609,G58610,G58611,G58612,G58613,G58614,G58615,G58616,G58617,G58618,G58619,G58620,
       G58621,G58622,G58623,G58624,G58625,G58626,G58627,G58628,G58629,G58630,G58631,G58632,G58633,G58634,G58635,G58636,G58637,G58638,G58639,G58640,
       G58641,G58642,G58643,G58644,G58645,G58646,G58647,G58648,G58649,G58650,G58651,G58652,G58653,G58654,G58655,G58656,G58657,G58658,G58659,G58660,
       G58661,G58662,G58663,G58664,G58665,G58666,G58667,G58668,G58669,G58670,G58671,G58672,G58673,G58674,G58675,G58676,G58677,G58678,G58679,G58680,
       G58681,G58682,G58683,G58684,G58685,G58686,G58687,G58688,G58689,G58690,G58691,G58692,G58693,G58694,G58695,G58696,G58697,G58698,G58699,G58700,
       G58701,G58702,G58703,G58704,G58705,G58706,G58707,G58708,G58709,G58710,G58711,G58712,G58713,G58714,G58715,G58716,G58717,G58718,G58719,G58720,
       G58721,G58722,G58723,G58724,G58725,G58726,G58727,G58728,G58729,G58730,G58731,G58732,G58733,G58734,G58735,G58736,G58737,G58738,G58739,G58740,
       G58741,G58742,G58743,G58744,G58745,G58746,G58747,G58748,G58749,G58750,G58751,G58752,G58753,G58754,G58755,G58756,G58757,G58758,G58759,G58760,
       G58761,G58762,G58763,G58764,G58765,G58766,G58767,G58768,G58769,G58770,G58771,G58772,G58773,G58774,G58775,G58776,G58777,G58778,G58779,G58780,
       G58781,G58782,G58783,G58784,G58785,G58786,G58787,G58788,G58789,G58790,G58791,G58792,G58793,G58794,G58795,G58796,G58797,G58798,G58799,G58800,
       G58801,G58802,G58803,G58804,G58805,G58806,G58807,G58808,G58809,G58810,G58811,G58812,G58813,G58814,G58815,G58816,G58817,G58818,G58819,G58820,
       G58821,G58822,G58823,G58824,G58825,G58826,G58827,G58828,G58829,G58830,G58831,G58832,G58833,G58834,G58835,G58836,G58837,G58838,G58839,G58840,
       G58841,G58842,G58843,G58844,G58845,G58846,G58847,G58848,G58849,G58850,G58851,G58852,G58853,G58854,G58855,G58856,G58857,G58858,G58859,G58860,
       G58861,G58862,G58863,G58864,G58865,G58866,G58867,G58868,G58869,G58870,G58871,G58872,G58873,G58874,G58875,G58876,G58877,G58878,G58879,G58880,
       G58881,G58882,G58883,G58884,G58885,G58886,G58887,G58888,G58889,G58890,G58891,G58892,G58893,G58894,G58895,G58896,G58897,G58898,G58899,G58900,
       G58901,G58902,G58903,G58904,G58905,G58906,G58907,G58908,G58909,G58910,G58911,G58912,G58913,G58914,G58915,G58916,G58917,G58918,G58919,G58920,
       G58921,G58922,G58923,G58924,G58925,G58926,G58927,G58928,G58929,G58930,G58931,G58932,G58933,G58934,G58935,G58936,G58937,G58938,G58939,G58940,
       G58941,G58942,G58943,G58944,G58945,G58946,G58947,G58948,G58949,G58950,G58951,G58952,G58953,G58954,G58955,G58956,G58957,G58958,G58959,G58960,
       G58961,G58962,G58963,G58964,G58965,G58966,G58967,G58968,G58969,G58970,G58971,G58972,G58973,G58974,G58975,G58976,G58977,G58978,G58979,G58980,
       G58981,G58982,G58983,G58984,G58985,G58986,G58987,G58988,G58989,G58990,G58991,G58992,G58993,G58994,G58995,G58996,G58997,G58998,G58999,G59000,
       G59001,G59002,G59003,G59004,G59005,G59006,G59007,G59008,G59009,G59010,G59011,G59012,G59013,G59014,G59015,G59016,G59017,G59018,G59019,G59020,
       G59021,G59022,G59023,G59024,G59025,G59026,G59027,G59028,G59029,G59030,G59031,G59032,G59033,G59034,G59035,G59036,G59037,G59038,G59039,G59040,
       G59041,G59042,G59043,G59044,G59045,G59046,G59047,G59048,G59049,G59050,G59051,G59052,G59053,G59054,G59055,G59056,G59057,G59058,G59059,G59060,
       G59061,G59062,G59063,G59064,G59065,G59066,G59067,G59068,G59069,G59070,G59071,G59072,G59073,G59074,G59075,G59076,G59077,G59078,G59079,G59080,
       G59081,G59082,G59083,G59084,G59085,G59086,G59087,G59088,G59089,G59090,G59091,G59092,G59093,G59094,G59095,G59096,G59097,G59098,G59099,G59100,
       G59101,G59102,G59103,G59104,G59105,G59106,G59107,G59108,G59109,G59110,G59111,G59112,G59113,G59114,G59115,G59116,G59117,G59118,G59119,G59120,
       G59121,G59122,G59123,G59124,G59125,G59126,G59127,G59128,G59129,G59130,G59131,G59132,G59133,G59134,G59135,G59136,G59137,G59138,G59139,G59140,
       G59141,G59142,G59143,G59144,G59145,G59146,G59147,G59148,G59149,G59150,G59151,G59152,G59153,G59154,G59155,G59156,G59157,G59158,G59159,G59160,
       G59161,G59162,G59163,G59164,G59165,G59166,G59167,G59168,G59169,G59170,G59171,G59172,G59173,G59174,G59175,G59176,G59177,G59178,G59179,G59180,
       G59181,G59182,G59183,G59184,G59185,G59186,G59187,G59188,G59189,G59190,G59191,G59192,G59193,G59194,G59195,G59196,G59197,G59198,G59199,G59200,
       G59201,G59202,G59203,G59204,G59205,G59206,G59207,G59208,G59209,G59210,G59211,G59212,G59213,G59214,G59215,G59216,G59217,G59218,G59219,G59220,
       G59221,G59222,G59223,G59224,G59225,G59226,G59227,G59228,G59229,G59230,G59231,G59232,G59233,G59234,G59235,G59236,G59237,G59238,G59239,G59240,
       G59241,G59242,G59243,G59244,G59245,G59246,G59247,G59248,G59249,G59250,G59251,G59252,G59253,G59254,G59255,G59256,G59257,G59258,G59259,G59260,
       G59261,G59262,G59263,G59264,G59265,G59266,G59267,G59268,G59269,G59270,G59271,G59272,G59273,G59274,G59275,G59276,G59277,G59278,G59279,G59280,
       G59281,G59282,G59283,G59284,G59285,G59286,G59287,G59288,G59289,G59290,G59291,G59292,G59293,G59294,G59295,G59296,G59297,G59298,G59299,G59300,
       G59301,G59302,G59303,G59304,G59305,G59306,G59307,G59308,G59309,G59310,G59311,G59312,G59313,G59314,G59315,G59316,G59317,G59318,G59319,G59320,
       G59321,G59322,G59323,G59324,G59325,G59326,G59327,G59328,G59329,G59330,G59331,G59332,G59333,G59334,G59335,G59336,G59337,G59338,G59339,G59340,
       G59341,G59342,G59343,G59344,G59345,G59346,G59347,G59348,G59349,G59350,G59351,G59352,G59353,G59354,G59355,G59356,G59357,G59358,G59359,G59360,
       G59361,G59362,G59363,G59364,G59365,G59366,G59367,G59368,G59369,G59370,G59371,G59372,G59373,G59374,G59375,G59376,G59377,G59378,G59379,G59380,
       G59381,G59382,G59383,G59384,G59385,G59386,G59387,G59388,G59389,G59390,G59391,G59392,G59393,G59394,G59395,G59396,G59397,G59398,G59399,G59400,
       G59401,G59402,G59403,G59404,G59405,G59406,G59407,G59408,G59409,G59410,G59411,G59412,G59413,G59414,G59415,G59416,G59417,G59418,G59419,G59420,
       G59421,G59422,G59423,G59424,G59425,G59426,G59427,G59428,G59429,G59430,G59431,G59432,G59433,G59434,G59435,G59436,G59437,G59438,G59439,G59440,
       G59441,G59442,G59443,G59444,G59445,G59446,G59447,G59448,G59449,G59450,G59451,G59452,G59453,G59454,G59455,G59456,G59457,G59458,G59459,G59460,
       G59461,G59462,G59463,G59464,G59465,G59466,G59467,G59468,G59469,G59470,G59471,G59472,G59473,G59474,G59475,G59476,G59477,G59478,G59479,G59480,
       G59481,G59482,G59483,G59484,G59485,G59486,G59487,G59488,G59489,G59490,G59491,G59492,G59493,G59494,G59495,G59496,G59497,G59498,G59499,G59500,
       G59501,G59502,G59503,G59504,G59505,G59506,G59507,G59508,G59509,G59510,G59511,G59512,G59513,G59514,G59515,G59516,G59517,G59518,G59519,G59520,
       G59521,G59522,G59523,G59524,G59525,G59526,G59527,G59528,G59529,G59530,G59531,G59532,G59533,G59534,G59535,G59536,G59537,G59538,G59539,G59540,
       G59541,G59542,G59543,G59544,G59545,G59546,G59547,G59548,G59549,G59550,G59551,G59552,G59553,G59554,G59555,G59556,G59557,G59558,G59559,G59560,
       G59561,G59562,G59563,G59564,G59565,G59566,G59567,G59568,G59569,G59570,G59571,G59572,G59573,G59574,G59575,G59576,G59577,G59578,G59579,G59580,
       G59581,G59582,G59583,G59584,G59585,G59586,G59587,G59588,G59589,G59590,G59591,G59592,G59593,G59594,G59595,G59596,G59597,G59598,G59599,G59600,
       G59601,G59602,G59603,G59604,G59605,G59606,G59607,G59608,G59609,G59610,G59611,G59612,G59613,G59614,G59615,G59616,G59617,G59618,G59619,G59620,
       G59621,G59622,G59623,G59624,G59625,G59626,G59627,G59628,G59629,G59630,G59631,G59632,G59633,G59634,G59635,G59636,G59637,G59638,G59639,G59640,
       G59641,G59642,G59643,G59644,G59645,G59646,G59647,G59648,G59649,G59650,G59651,G59652,G59653,G59654,G59655,G59656,G59657,G59658,G59659,G59660,
       G59661,G59662,G59663,G59664,G59665,G59666,G59667,G59668,G59669,G59670,G59671,G59672,G59673,G59674,G59675,G59676,G59677,G59678,G59679,G59680,
       G59681,G59682,G59683,G59684,G59685,G59686,G59687,G59688,G59689,G59690,G59691,G59692,G59693,G59694,G59695,G59696,G59697,G59698,G59699,G59700,
       G59701,G59702,G59703,G59704,G59705,G59706,G59707,G59708,G59709,G59710,G59711,G59712,G59713,G59714,G59715,G59716,G59717,G59718,G59719,G59720,
       G59721,G59722,G59723,G59724,G59725,G59726,G59727,G59728,G59729,G59730,G59731,G59732,G59733,G59734,G59735,G59736,G59737,G59738,G59739,G59740,
       G59741,G59742,G59743,G59744,G59745,G59746,G59747,G59748,G59749,G59750,G59751,G59752,G59753,G59754,G59755,G59756,G59757,G59758,G59759,G59760,
       G59761,G59762,G59763,G59764,G59765,G59766,G59767,G59768,G59769,G59770,G59771,G59772,G59773,G59774,G59775,G59776,G59777,G59778,G59779,G59780,
       G59781,G59782,G59783,G59784,G59785,G59786,G59787,G59788,G59789,G59790,G59791,G59792,G59793,G59794,G59795,G59796,G59797,G59798,G59799,G59800,
       G59801,G59802,G59803,G59804,G59805,G59806,G59807,G59808,G59809,G59810,G59811,G59812,G59813,G59814,G59815,G59816,G59817,G59818,G59819,G59820,
       G59821,G59822,G59823,G59824,G59825,G59826,G59827,G59828,G59829,G59830,G59831,G59832,G59833,G59834,G59835,G59836,G59837,G59838,G59839,G59840,
       G59841,G59842,G59843,G59844,G59845,G59846,G59847,G59848,G59849,G59850,G59851,G59852,G59853,G59854,G59855,G59856,G59857,G59858,G59859,G59860,
       G59861,G59862,G59863,G59864,G59865,G59866,G59867,G59868,G59869,G59870,G59871,G59872,G59873,G59874,G59875,G59876,G59877,G59878,G59879,G59880,
       G59881,G59882,G59883,G59884,G59885,G59886,G59887,G59888,G59889,G59890,G59891,G59892,G59893,G59894,G59895,G59896,G59897,G59898,G59899,G59900,
       G59901,G59902,G59903,G59904,G59905,G59906,G59907,G59908,G59909,G59910,G59911,G59912,G59913,G59914,G59915,G59916,G59917,G59918,G59919,G59920,
       G59921,G59922,G59923,G59924,G59925,G59926,G59927,G59928,G59929,G59930,G59931,G59932,G59933,G59934,G59935,G59936,G59937,G59938,G59939,G59940,
       G59941,G59942,G59943,G59944,G59945,G59946,G59947,G59948,G59949,G59950,G59951,G59952,G59953,G59954,G59955,G59956,G59957,G59958,G59959,G59960,
       G59961,G59962,G59963,G59964,G59965,G59966,G59967,G59968,G59969,G59970,G59971,G59972,G59973,G59974,G59975,G59976,G59977,G59978,G59979,G59980,
       G59981,G59982,G59983,G59984,G59985,G59986,G59987,G59988,G59989,G59990,G59991,G59992,G59993,G59994,G59995,G59996,G59997,G59998,G59999,G60000,
       G60001,G60002,G60003,G60004,G60005,G60006,G60007,G60008,G60009,G60010,G60011,G60012,G60013,G60014,G60015,G60016,G60017,G60018,G60019,G60020,
       G60021,G60022,G60023,G60024,G60025,G60026,G60027,G60028,G60029,G60030,G60031,G60032,G60033,G60034,G60035,G60036,G60037,G60038,G60039,G60040,
       G60041,G60042,G60043,G60044,G60045,G60046,G60047,G60048,G60049,G60050,G60051,G60052,G60053,G60054,G60055,G60056,G60057,G60058,G60059,G60060,
       G60061,G60062,G60063,G60064,G60065,G60066,G60067,G60068,G60069,G60070,G60071,G60072,G60073,G60074,G60075,G60076,G60077,G60078,G60079,G60080,
       G60081,G60082,G60083,G60084,G60085,G60086,G60087,G60088,G60089,G60090,G60091,G60092,G60093,G60094,G60095,G60096,G60097,G60098,G60099,G60100,
       G60101,G60102,G60103,G60104,G60105,G60106,G60107,G60108,G60109,G60110,G60111,G60112,G60113,G60114,G60115,G60116,G60117,G60118,G60119,G60120,
       G60121,G60122,G60123,G60124,G60125,G60126,G60127,G60128,G60129,G60130,G60131,G60132,G60133,G60134,G60135,G60136,G60137,G60138,G60139,G60140,
       G60141,G60142,G60143,G60144,G60145,G60146,G60147,G60148,G60149,G60150,G60151,G60152,G60153,G60154,G60155,G60156,G60157,G60158,G60159,G60160,
       G60161,G60162,G60163,G60164,G60165,G60166,G60167,G60168,G60169,G60170,G60171,G60172,G60173,G60174,G60175,G60176,G60177,G60178,G60179,G60180,
       G60181,G60182,G60183,G60184,G60185,G60186,G60187,G60188,G60189,G60190,G60191,G60192,G60193,G60194,G60195,G60196,G60197,G60198,G60199,G60200,
       G60201,G60202,G60203,G60204,G60205,G60206,G60207,G60208,G60209,G60210,G60211,G60212,G60213,G60214,G60215,G60216,G60217,G60218,G60219,G60220,
       G60221,G60222,G60223,G60224,G60225,G60226,G60227,G60228,G60229,G60230,G60231,G60232,G60233,G60234,G60235,G60236,G60237,G60238,G60239,G60240,
       G60241,G60242,G60243,G60244,G60245,G60246,G60247,G60248,G60249,G60250,G60251,G60252,G60253;

  dff DFF_135(CK,G58839,G1556);
  dff DFF_136(CK,G58840,G1557);
  dff DFF_137(CK,G58841,G1558);
  dff DFF_138(CK,G58842,G1559);
  dff DFF_139(CK,G58843,G1560);
  dff DFF_140(CK,G58844,G1561);
  dff DFF_141(CK,G58845,G1562);
  dff DFF_142(CK,G58846,G1563);
  dff DFF_143(CK,G58847,G1564);
  dff DFF_144(CK,G58848,G1565);
  dff DFF_145(CK,G58849,G1566);
  dff DFF_146(CK,G58850,G1567);
  dff DFF_147(CK,G58851,G1568);
  dff DFF_148(CK,G58852,G1569);
  dff DFF_149(CK,G58853,G1570);
  dff DFF_150(CK,G58854,G1571);
  dff DFF_151(CK,G58855,G1572);
  dff DFF_152(CK,G58856,G1573);
  dff DFF_153(CK,G58857,G1574);
  dff DFF_154(CK,G58858,G1575);
  dff DFF_155(CK,G58859,G1576);
  dff DFF_156(CK,G58860,G1577);
  dff DFF_157(CK,G58861,G1578);
  dff DFF_158(CK,G58862,G1579);
  dff DFF_159(CK,G58863,G1580);
  dff DFF_160(CK,G58864,G1581);
  dff DFF_161(CK,G58865,G1582);
  dff DFF_162(CK,G58866,G1583);
  dff DFF_163(CK,G58867,G1584);
  dff DFF_164(CK,G58868,G1585);
  dff DFF_165(CK,G58869,G1586);
  dff DFF_166(CK,G58870,G1587);
  dff DFF_167(CK,G58871,G1596);
  dff DFF_168(CK,G58872,G1597);
  dff DFF_169(CK,G58873,G1598);
  dff DFF_170(CK,G58874,G1599);
  dff DFF_171(CK,G58875,G1600);
  dff DFF_172(CK,G58876,G1601);
  dff DFF_173(CK,G58877,G1602);
  dff DFF_174(CK,G58878,G1603);
  dff DFF_175(CK,G58879,G1604);
  dff DFF_176(CK,G58880,G1605);
  dff DFF_177(CK,G58881,G1606);
  dff DFF_178(CK,G58882,G1607);
  dff DFF_179(CK,G58883,G1608);
  dff DFF_180(CK,G58884,G1609);
  dff DFF_181(CK,G58885,G1610);
  dff DFF_182(CK,G58886,G1611);
  dff DFF_183(CK,G58887,G1612);
  dff DFF_184(CK,G58888,G1613);
  dff DFF_185(CK,G58889,G1614);
  dff DFF_186(CK,G58890,G1615);
  dff DFF_187(CK,G58891,G1616);
  dff DFF_188(CK,G58892,G1617);
  dff DFF_189(CK,G58893,G1618);
  dff DFF_190(CK,G58894,G1619);
  dff DFF_191(CK,G58895,G1620);
  dff DFF_192(CK,G58896,G1621);
  dff DFF_193(CK,G58897,G1622);
  dff DFF_194(CK,G58898,G1623);
  dff DFF_195(CK,G58899,G1624);
  dff DFF_196(CK,G58900,G1625);
  dff DFF_197(CK,G58901,G1626);
  dff DFF_198(CK,G58902,G1627);
  dff DFF_199(CK,G58903,G1552);
  dff DFF_200(CK,G58904,G1731);
  dff DFF_201(CK,G58905,G1553);
  dff DFF_202(CK,G58906,G1730);
  dff DFF_203(CK,G58907,G3276);
  dff DFF_204(CK,G58908,G3275);
  dff DFF_205(CK,G58909,G3274);
  dff DFF_206(CK,G58910,G3273);
  dff DFF_207(CK,G58911,G2314);
  dff DFF_208(CK,G58912,G2315);
  dff DFF_209(CK,G58913,G2316);
  dff DFF_210(CK,G58914,G2317);
  dff DFF_211(CK,G58915,G2318);
  dff DFF_212(CK,G58916,G2319);
  dff DFF_213(CK,G58917,G2320);
  dff DFF_214(CK,G58918,G2321);
  dff DFF_215(CK,G58919,G2322);
  dff DFF_216(CK,G58920,G2323);
  dff DFF_217(CK,G58921,G2324);
  dff DFF_218(CK,G58922,G2325);
  dff DFF_219(CK,G58923,G2326);
  dff DFF_220(CK,G58924,G2327);
  dff DFF_221(CK,G58925,G2328);
  dff DFF_222(CK,G58926,G2329);
  dff DFF_223(CK,G58927,G2330);
  dff DFF_224(CK,G58928,G2331);
  dff DFF_225(CK,G58929,G2332);
  dff DFF_226(CK,G58930,G2333);
  dff DFF_227(CK,G58931,G2334);
  dff DFF_228(CK,G58932,G2335);
  dff DFF_229(CK,G58933,G2336);
  dff DFF_230(CK,G58934,G2337);
  dff DFF_231(CK,G58935,G2338);
  dff DFF_232(CK,G58936,G2339);
  dff DFF_233(CK,G58937,G2340);
  dff DFF_234(CK,G58938,G2341);
  dff DFF_235(CK,G58939,G2342);
  dff DFF_236(CK,G58940,G2343);
  dff DFF_237(CK,G58941,G2344);
  dff DFF_238(CK,G58942,G2345);
  dff DFF_239(CK,G58943,G2346);
  dff DFF_240(CK,G58944,G3272);
  dff DFF_241(CK,G58945,G3271);
  dff DFF_242(CK,G58946,G2347);
  dff DFF_243(CK,G58947,G2348);
  dff DFF_244(CK,G58948,G2349);
  dff DFF_245(CK,G58949,G2350);
  dff DFF_246(CK,G58950,G2351);
  dff DFF_247(CK,G58951,G2352);
  dff DFF_248(CK,G58952,G2353);
  dff DFF_249(CK,G58953,G2354);
  dff DFF_250(CK,G58954,G2355);
  dff DFF_251(CK,G58955,G2356);
  dff DFF_252(CK,G58956,G2357);
  dff DFF_253(CK,G58957,G2358);
  dff DFF_254(CK,G58958,G2359);
  dff DFF_255(CK,G58959,G2360);
  dff DFF_256(CK,G58960,G2361);
  dff DFF_257(CK,G58961,G2362);
  dff DFF_258(CK,G58962,G2363);
  dff DFF_259(CK,G58963,G2364);
  dff DFF_260(CK,G58964,G2365);
  dff DFF_261(CK,G58965,G2366);
  dff DFF_262(CK,G58966,G2367);
  dff DFF_263(CK,G58967,G2368);
  dff DFF_264(CK,G58968,G2369);
  dff DFF_265(CK,G58969,G2370);
  dff DFF_266(CK,G58970,G2371);
  dff DFF_267(CK,G58971,G2372);
  dff DFF_268(CK,G58972,G2373);
  dff DFF_269(CK,G58973,G2374);
  dff DFF_270(CK,G58974,G2375);
  dff DFF_271(CK,G58975,G2376);
  dff DFF_272(CK,G58976,G2377);
  dff DFF_273(CK,G58977,G2378);
  dff DFF_274(CK,G58978,G2379);
  dff DFF_275(CK,G58979,G2380);
  dff DFF_276(CK,G58980,G2381);
  dff DFF_277(CK,G58981,G2382);
  dff DFF_278(CK,G58982,G2383);
  dff DFF_279(CK,G58983,G2384);
  dff DFF_280(CK,G58984,G2385);
  dff DFF_281(CK,G58985,G2386);
  dff DFF_282(CK,G58986,G2387);
  dff DFF_283(CK,G58987,G2388);
  dff DFF_284(CK,G58988,G2389);
  dff DFF_285(CK,G58989,G2390);
  dff DFF_286(CK,G58990,G2391);
  dff DFF_287(CK,G58991,G2392);
  dff DFF_288(CK,G58992,G2393);
  dff DFF_289(CK,G58993,G2394);
  dff DFF_290(CK,G58994,G2395);
  dff DFF_291(CK,G58995,G2396);
  dff DFF_292(CK,G58996,G2397);
  dff DFF_293(CK,G58997,G2398);
  dff DFF_294(CK,G58998,G2399);
  dff DFF_295(CK,G58999,G2400);
  dff DFF_296(CK,G59000,G2401);
  dff DFF_297(CK,G59001,G2402);
  dff DFF_298(CK,G59002,G2403);
  dff DFF_299(CK,G59003,G2404);
  dff DFF_300(CK,G59004,G2405);
  dff DFF_301(CK,G59005,G2406);
  dff DFF_302(CK,G59006,G2407);
  dff DFF_303(CK,G59007,G2408);
  dff DFF_304(CK,G59008,G2409);
  dff DFF_305(CK,G59009,G2410);
  dff DFF_306(CK,G59010,G2411);
  dff DFF_307(CK,G59011,G2412);
  dff DFF_308(CK,G59012,G2413);
  dff DFF_309(CK,G59013,G2414);
  dff DFF_310(CK,G59014,G2415);
  dff DFF_311(CK,G59015,G2416);
  dff DFF_312(CK,G59016,G2417);
  dff DFF_313(CK,G59017,G2418);
  dff DFF_314(CK,G59018,G2419);
  dff DFF_315(CK,G59019,G2420);
  dff DFF_316(CK,G59020,G2421);
  dff DFF_317(CK,G59021,G2422);
  dff DFF_318(CK,G59022,G2423);
  dff DFF_319(CK,G59023,G2424);
  dff DFF_320(CK,G59024,G2425);
  dff DFF_321(CK,G59025,G2426);
  dff DFF_322(CK,G59026,G2427);
  dff DFF_323(CK,G59027,G2428);
  dff DFF_324(CK,G59028,G2429);
  dff DFF_325(CK,G59029,G2430);
  dff DFF_326(CK,G59030,G2431);
  dff DFF_327(CK,G59031,G2432);
  dff DFF_328(CK,G59032,G2433);
  dff DFF_329(CK,G59033,G2434);
  dff DFF_330(CK,G59034,G2435);
  dff DFF_331(CK,G59035,G2436);
  dff DFF_332(CK,G59036,G2437);
  dff DFF_333(CK,G59037,G2438);
  dff DFF_334(CK,G59038,G2439);
  dff DFF_335(CK,G59039,G2440);
  dff DFF_336(CK,G59040,G2441);
  dff DFF_337(CK,G59041,G2442);
  dff DFF_338(CK,G59042,G2443);
  dff DFF_339(CK,G59043,G2444);
  dff DFF_340(CK,G59044,G2445);
  dff DFF_341(CK,G59045,G2446);
  dff DFF_342(CK,G59046,G2447);
  dff DFF_343(CK,G59047,G2448);
  dff DFF_344(CK,G59048,G2449);
  dff DFF_345(CK,G59049,G2450);
  dff DFF_346(CK,G59050,G2451);
  dff DFF_347(CK,G59051,G2452);
  dff DFF_348(CK,G59052,G2453);
  dff DFF_349(CK,G59053,G2454);
  dff DFF_350(CK,G59054,G2455);
  dff DFF_351(CK,G59055,G2456);
  dff DFF_352(CK,G59056,G2457);
  dff DFF_353(CK,G59057,G2458);
  dff DFF_354(CK,G59058,G2459);
  dff DFF_355(CK,G59059,G2460);
  dff DFF_356(CK,G59060,G2461);
  dff DFF_357(CK,G59061,G2462);
  dff DFF_358(CK,G59062,G2463);
  dff DFF_359(CK,G59063,G2464);
  dff DFF_360(CK,G59064,G2465);
  dff DFF_361(CK,G59065,G2466);
  dff DFF_362(CK,G59066,G2467);
  dff DFF_363(CK,G59067,G2468);
  dff DFF_364(CK,G59068,G2469);
  dff DFF_365(CK,G59069,G2470);
  dff DFF_366(CK,G59070,G2471);
  dff DFF_367(CK,G59071,G2472);
  dff DFF_368(CK,G59072,G2473);
  dff DFF_369(CK,G59073,G2474);
  dff DFF_370(CK,G59074,G2475);
  dff DFF_371(CK,G59075,G2476);
  dff DFF_372(CK,G59076,G2477);
  dff DFF_373(CK,G59077,G2478);
  dff DFF_374(CK,G59078,G2479);
  dff DFF_375(CK,G59079,G2480);
  dff DFF_376(CK,G59080,G2481);
  dff DFF_377(CK,G59081,G2482);
  dff DFF_378(CK,G59082,G2483);
  dff DFF_379(CK,G59083,G2484);
  dff DFF_380(CK,G59084,G2485);
  dff DFF_381(CK,G59085,G2486);
  dff DFF_382(CK,G59086,G2487);
  dff DFF_383(CK,G59087,G2488);
  dff DFF_384(CK,G59088,G2489);
  dff DFF_385(CK,G59089,G2490);
  dff DFF_386(CK,G59090,G2491);
  dff DFF_387(CK,G59091,G2492);
  dff DFF_388(CK,G59092,G2493);
  dff DFF_389(CK,G59093,G2494);
  dff DFF_390(CK,G59094,G2495);
  dff DFF_391(CK,G59095,G2496);
  dff DFF_392(CK,G59096,G2497);
  dff DFF_393(CK,G59097,G2498);
  dff DFF_394(CK,G59098,G2499);
  dff DFF_395(CK,G59099,G2500);
  dff DFF_396(CK,G59100,G2501);
  dff DFF_397(CK,G59101,G2502);
  dff DFF_398(CK,G59102,G2503);
  dff DFF_399(CK,G59103,G2504);
  dff DFF_400(CK,G59104,G2505);
  dff DFF_401(CK,G59105,G2506);
  dff DFF_402(CK,G59106,G2507);
  dff DFF_403(CK,G59107,G2508);
  dff DFF_404(CK,G59108,G3270);
  dff DFF_405(CK,G59109,G3269);
  dff DFF_406(CK,G59110,G3268);
  dff DFF_407(CK,G59111,G3266);
  dff DFF_408(CK,G59112,G3265);
  dff DFF_409(CK,G59113,G2509);
  dff DFF_410(CK,G59114,G2510);
  dff DFF_411(CK,G59115,G2511);
  dff DFF_412(CK,G59116,G2512);
  dff DFF_413(CK,G59117,G2747);
  dff DFF_414(CK,G59118,G2513);
  dff DFF_415(CK,G59119,G2514);
  dff DFF_416(CK,G59120,G2515);
  dff DFF_417(CK,G59121,G2516);
  dff DFF_418(CK,G59122,G2517);
  dff DFF_419(CK,G59123,G2518);
  dff DFF_420(CK,G59124,G2519);
  dff DFF_421(CK,G59125,G2520);
  dff DFF_422(CK,G59126,G2521);
  dff DFF_423(CK,G59127,G2522);
  dff DFF_424(CK,G59128,G2523);
  dff DFF_425(CK,G59129,G2524);
  dff DFF_426(CK,G59130,G2525);
  dff DFF_427(CK,G59131,G2526);
  dff DFF_428(CK,G59132,G2527);
  dff DFF_429(CK,G59133,G2528);
  dff DFF_430(CK,G59134,G2529);
  dff DFF_431(CK,G59135,G2530);
  dff DFF_432(CK,G59136,G2531);
  dff DFF_433(CK,G59137,G2532);
  dff DFF_434(CK,G59138,G2533);
  dff DFF_435(CK,G59139,G2534);
  dff DFF_436(CK,G59140,G2535);
  dff DFF_437(CK,G59141,G2536);
  dff DFF_438(CK,G59142,G2537);
  dff DFF_439(CK,G59143,G2538);
  dff DFF_440(CK,G59144,G2539);
  dff DFF_441(CK,G59145,G2540);
  dff DFF_442(CK,G59146,G2541);
  dff DFF_443(CK,G59147,G2542);
  dff DFF_444(CK,G59148,G2543);
  dff DFF_445(CK,G59149,G2544);
  dff DFF_446(CK,G59150,G2545);
  dff DFF_447(CK,G59151,G2546);
  dff DFF_448(CK,G59152,G2547);
  dff DFF_449(CK,G59153,G2548);
  dff DFF_450(CK,G59154,G2549);
  dff DFF_451(CK,G59155,G2550);
  dff DFF_452(CK,G59156,G2551);
  dff DFF_453(CK,G59157,G2552);
  dff DFF_454(CK,G59158,G2553);
  dff DFF_455(CK,G59159,G2554);
  dff DFF_456(CK,G59160,G2555);
  dff DFF_457(CK,G59161,G2556);
  dff DFF_458(CK,G59162,G2557);
  dff DFF_459(CK,G59163,G2558);
  dff DFF_460(CK,G59164,G2559);
  dff DFF_461(CK,G59165,G2560);
  dff DFF_462(CK,G59166,G2561);
  dff DFF_463(CK,G59167,G2562);
  dff DFF_464(CK,G59168,G2563);
  dff DFF_465(CK,G59169,G2564);
  dff DFF_466(CK,G59170,G2565);
  dff DFF_467(CK,G59171,G2566);
  dff DFF_468(CK,G59172,G2567);
  dff DFF_469(CK,G59173,G2568);
  dff DFF_470(CK,G59174,G2569);
  dff DFF_471(CK,G59175,G2570);
  dff DFF_472(CK,G59176,G2571);
  dff DFF_473(CK,G59177,G2572);
  dff DFF_474(CK,G59178,G2573);
  dff DFF_475(CK,G59179,G2574);
  dff DFF_476(CK,G59180,G2575);
  dff DFF_477(CK,G59181,G2576);
  dff DFF_478(CK,G59182,G2577);
  dff DFF_479(CK,G59183,G2578);
  dff DFF_480(CK,G59184,G2579);
  dff DFF_481(CK,G59185,G2580);
  dff DFF_482(CK,G59186,G2581);
  dff DFF_483(CK,G59187,G2582);
  dff DFF_484(CK,G59188,G2583);
  dff DFF_485(CK,G59189,G2584);
  dff DFF_486(CK,G59190,G2585);
  dff DFF_487(CK,G59191,G2586);
  dff DFF_488(CK,G59192,G2587);
  dff DFF_489(CK,G59193,G2588);
  dff DFF_490(CK,G59194,G2589);
  dff DFF_491(CK,G59195,G2590);
  dff DFF_492(CK,G59196,G2591);
  dff DFF_493(CK,G59197,G2592);
  dff DFF_494(CK,G59198,G2593);
  dff DFF_495(CK,G59199,G2594);
  dff DFF_496(CK,G59200,G2595);
  dff DFF_497(CK,G59201,G2596);
  dff DFF_498(CK,G59202,G2597);
  dff DFF_499(CK,G59203,G2598);
  dff DFF_500(CK,G59204,G2599);
  dff DFF_501(CK,G59205,G2600);
  dff DFF_502(CK,G59206,G2601);
  dff DFF_503(CK,G59207,G2602);
  dff DFF_504(CK,G59208,G2603);
  dff DFF_505(CK,G59209,G2604);
  dff DFF_506(CK,G59210,G2605);
  dff DFF_507(CK,G59211,G2606);
  dff DFF_508(CK,G59212,G2607);
  dff DFF_509(CK,G59213,G2608);
  dff DFF_510(CK,G59214,G2609);
  dff DFF_511(CK,G59215,G2610);
  dff DFF_512(CK,G59216,G2611);
  dff DFF_513(CK,G59217,G2612);
  dff DFF_514(CK,G59218,G2613);
  dff DFF_515(CK,G59219,G2614);
  dff DFF_516(CK,G59220,G2615);
  dff DFF_517(CK,G59221,G2616);
  dff DFF_518(CK,G59222,G2617);
  dff DFF_519(CK,G59223,G2618);
  dff DFF_520(CK,G59224,G2619);
  dff DFF_521(CK,G59225,G2620);
  dff DFF_522(CK,G59226,G2621);
  dff DFF_523(CK,G59227,G2622);
  dff DFF_524(CK,G59228,G2623);
  dff DFF_525(CK,G59229,G2624);
  dff DFF_526(CK,G59230,G2625);
  dff DFF_527(CK,G59231,G2626);
  dff DFF_528(CK,G59232,G2627);
  dff DFF_529(CK,G59233,G2628);
  dff DFF_530(CK,G59234,G2629);
  dff DFF_531(CK,G59235,G2630);
  dff DFF_532(CK,G59236,G2631);
  dff DFF_533(CK,G59237,G2632);
  dff DFF_534(CK,G59238,G2633);
  dff DFF_535(CK,G59239,G2634);
  dff DFF_536(CK,G59240,G2635);
  dff DFF_537(CK,G59241,G2636);
  dff DFF_538(CK,G59242,G2637);
  dff DFF_539(CK,G59243,G2638);
  dff DFF_540(CK,G59244,G2639);
  dff DFF_541(CK,G59245,G2640);
  dff DFF_542(CK,G59246,G2641);
  dff DFF_543(CK,G59247,G2642);
  dff DFF_544(CK,G59248,G2643);
  dff DFF_545(CK,G59249,G2644);
  dff DFF_546(CK,G59250,G2645);
  dff DFF_547(CK,G59251,G2646);
  dff DFF_548(CK,G59252,G2647);
  dff DFF_549(CK,G59253,G2648);
  dff DFF_550(CK,G59254,G2649);
  dff DFF_551(CK,G59255,G2650);
  dff DFF_552(CK,G59256,G2651);
  dff DFF_553(CK,G59257,G2652);
  dff DFF_554(CK,G59258,G2653);
  dff DFF_555(CK,G59259,G2654);
  dff DFF_556(CK,G59260,G2655);
  dff DFF_557(CK,G59261,G2656);
  dff DFF_558(CK,G59262,G2657);
  dff DFF_559(CK,G59263,G2658);
  dff DFF_560(CK,G59264,G2659);
  dff DFF_561(CK,G59265,G2660);
  dff DFF_562(CK,G59266,G2661);
  dff DFF_563(CK,G59267,G2662);
  dff DFF_564(CK,G59268,G2663);
  dff DFF_565(CK,G59269,G2664);
  dff DFF_566(CK,G59270,G2665);
  dff DFF_567(CK,G59271,G2666);
  dff DFF_568(CK,G59272,G2667);
  dff DFF_569(CK,G59273,G2668);
  dff DFF_570(CK,G59274,G2669);
  dff DFF_571(CK,G59275,G2670);
  dff DFF_572(CK,G59276,G2671);
  dff DFF_573(CK,G59277,G2672);
  dff DFF_574(CK,G59278,G2673);
  dff DFF_575(CK,G59279,G2674);
  dff DFF_576(CK,G59280,G2675);
  dff DFF_577(CK,G59281,G2676);
  dff DFF_578(CK,G59282,G2677);
  dff DFF_579(CK,G59283,G2678);
  dff DFF_580(CK,G59284,G2679);
  dff DFF_581(CK,G59285,G2680);
  dff DFF_582(CK,G59286,G2681);
  dff DFF_583(CK,G59287,G2682);
  dff DFF_584(CK,G59288,G2683);
  dff DFF_585(CK,G59289,G2684);
  dff DFF_586(CK,G59290,G2685);
  dff DFF_587(CK,G59291,G2686);
  dff DFF_588(CK,G59292,G2687);
  dff DFF_589(CK,G59293,G2688);
  dff DFF_590(CK,G59294,G2689);
  dff DFF_591(CK,G59295,G2690);
  dff DFF_592(CK,G59296,G2691);
  dff DFF_593(CK,G59297,G2692);
  dff DFF_594(CK,G59298,G2693);
  dff DFF_595(CK,G59299,G2694);
  dff DFF_596(CK,G59300,G2695);
  dff DFF_597(CK,G59301,G2696);
  dff DFF_598(CK,G59302,G2697);
  dff DFF_599(CK,G59303,G2698);
  dff DFF_600(CK,G59304,G2699);
  dff DFF_601(CK,G59305,G2700);
  dff DFF_602(CK,G59306,G2701);
  dff DFF_603(CK,G59307,G2702);
  dff DFF_604(CK,G59308,G2703);
  dff DFF_605(CK,G59309,G2704);
  dff DFF_606(CK,G59310,G2705);
  dff DFF_607(CK,G59311,G2706);
  dff DFF_608(CK,G59312,G2707);
  dff DFF_609(CK,G59313,G2708);
  dff DFF_610(CK,G59314,G2709);
  dff DFF_611(CK,G59315,G2710);
  dff DFF_612(CK,G59316,G2711);
  dff DFF_613(CK,G59317,G2712);
  dff DFF_614(CK,G59318,G2713);
  dff DFF_615(CK,G59319,G2714);
  dff DFF_616(CK,G59320,G2715);
  dff DFF_617(CK,G59321,G2716);
  dff DFF_618(CK,G59322,G2717);
  dff DFF_619(CK,G59323,G2718);
  dff DFF_620(CK,G59324,G2719);
  dff DFF_621(CK,G59325,G2720);
  dff DFF_622(CK,G59326,G2721);
  dff DFF_623(CK,G59327,G2722);
  dff DFF_624(CK,G59328,G2723);
  dff DFF_625(CK,G59329,G2724);
  dff DFF_626(CK,G59330,G2725);
  dff DFF_627(CK,G59331,G2726);
  dff DFF_628(CK,G59332,G2727);
  dff DFF_629(CK,G59333,G2728);
  dff DFF_630(CK,G59334,G2729);
  dff DFF_631(CK,G59335,G2730);
  dff DFF_632(CK,G59336,G2731);
  dff DFF_633(CK,G59337,G2732);
  dff DFF_634(CK,G59338,G2733);
  dff DFF_635(CK,G59339,G2734);
  dff DFF_636(CK,G59340,G2735);
  dff DFF_637(CK,G59341,G2736);
  dff DFF_638(CK,G59342,G2737);
  dff DFF_639(CK,G59343,G2738);
  dff DFF_640(CK,G59344,G2739);
  dff DFF_641(CK,G59345,G3264);
  dff DFF_642(CK,G59346,G2740);
  dff DFF_643(CK,G59347,G2741);
  dff DFF_644(CK,G59348,G2742);
  dff DFF_645(CK,G59349,G3263);
  dff DFF_646(CK,G59350,G2743);
  dff DFF_647(CK,G59351,G3262);
  dff DFF_648(CK,G59352,G2744);
  dff DFF_649(CK,G59353,G2745);
  dff DFF_650(CK,G59354,G3261);
  dff DFF_651(CK,G59355,G3260);
  dff DFF_652(CK,G59356,G9273);
  dff DFF_653(CK,G59357,G9272);
  dff DFF_654(CK,G59358,G9271);
  dff DFF_655(CK,G59359,G9270);
  dff DFF_656(CK,G59360,G8311);
  dff DFF_657(CK,G59361,G8312);
  dff DFF_658(CK,G59362,G8313);
  dff DFF_659(CK,G59363,G8314);
  dff DFF_660(CK,G59364,G8315);
  dff DFF_661(CK,G59365,G8316);
  dff DFF_662(CK,G59366,G8317);
  dff DFF_663(CK,G59367,G8318);
  dff DFF_664(CK,G59368,G8319);
  dff DFF_665(CK,G59369,G8320);
  dff DFF_666(CK,G59370,G8321);
  dff DFF_667(CK,G59371,G8322);
  dff DFF_668(CK,G59372,G8323);
  dff DFF_669(CK,G59373,G8324);
  dff DFF_670(CK,G59374,G8325);
  dff DFF_671(CK,G59375,G8326);
  dff DFF_672(CK,G59376,G8327);
  dff DFF_673(CK,G59377,G8328);
  dff DFF_674(CK,G59378,G8329);
  dff DFF_675(CK,G59379,G8330);
  dff DFF_676(CK,G59380,G8331);
  dff DFF_677(CK,G59381,G8332);
  dff DFF_678(CK,G59382,G8333);
  dff DFF_679(CK,G59383,G8334);
  dff DFF_680(CK,G59384,G8335);
  dff DFF_681(CK,G59385,G8336);
  dff DFF_682(CK,G59386,G8337);
  dff DFF_683(CK,G59387,G8338);
  dff DFF_684(CK,G59388,G8339);
  dff DFF_685(CK,G59389,G8340);
  dff DFF_686(CK,G59390,G8341);
  dff DFF_687(CK,G59391,G8342);
  dff DFF_688(CK,G59392,G8343);
  dff DFF_689(CK,G59393,G9269);
  dff DFF_690(CK,G59394,G9268);
  dff DFF_691(CK,G59395,G8344);
  dff DFF_692(CK,G59396,G8345);
  dff DFF_693(CK,G59397,G8346);
  dff DFF_694(CK,G59398,G8347);
  dff DFF_695(CK,G59399,G8348);
  dff DFF_696(CK,G59400,G8349);
  dff DFF_697(CK,G59401,G8350);
  dff DFF_698(CK,G59402,G8351);
  dff DFF_699(CK,G59403,G8352);
  dff DFF_700(CK,G59404,G8353);
  dff DFF_701(CK,G59405,G8354);
  dff DFF_702(CK,G59406,G8355);
  dff DFF_703(CK,G59407,G8356);
  dff DFF_704(CK,G59408,G8357);
  dff DFF_705(CK,G59409,G8358);
  dff DFF_706(CK,G59410,G8359);
  dff DFF_707(CK,G59411,G8360);
  dff DFF_708(CK,G59412,G8361);
  dff DFF_709(CK,G59413,G8362);
  dff DFF_710(CK,G59414,G8363);
  dff DFF_711(CK,G59415,G8364);
  dff DFF_712(CK,G59416,G8365);
  dff DFF_713(CK,G59417,G8366);
  dff DFF_714(CK,G59418,G8367);
  dff DFF_715(CK,G59419,G8368);
  dff DFF_716(CK,G59420,G8369);
  dff DFF_717(CK,G59421,G8370);
  dff DFF_718(CK,G59422,G8371);
  dff DFF_719(CK,G59423,G8372);
  dff DFF_720(CK,G59424,G8373);
  dff DFF_721(CK,G59425,G8374);
  dff DFF_722(CK,G59426,G8375);
  dff DFF_723(CK,G59427,G8376);
  dff DFF_724(CK,G59428,G8377);
  dff DFF_725(CK,G59429,G8378);
  dff DFF_726(CK,G59430,G8379);
  dff DFF_727(CK,G59431,G8380);
  dff DFF_728(CK,G59432,G8381);
  dff DFF_729(CK,G59433,G8382);
  dff DFF_730(CK,G59434,G8383);
  dff DFF_731(CK,G59435,G8384);
  dff DFF_732(CK,G59436,G8385);
  dff DFF_733(CK,G59437,G8386);
  dff DFF_734(CK,G59438,G8387);
  dff DFF_735(CK,G59439,G8388);
  dff DFF_736(CK,G59440,G8389);
  dff DFF_737(CK,G59441,G8390);
  dff DFF_738(CK,G59442,G8391);
  dff DFF_739(CK,G59443,G8392);
  dff DFF_740(CK,G59444,G8393);
  dff DFF_741(CK,G59445,G8394);
  dff DFF_742(CK,G59446,G8395);
  dff DFF_743(CK,G59447,G8396);
  dff DFF_744(CK,G59448,G8397);
  dff DFF_745(CK,G59449,G8398);
  dff DFF_746(CK,G59450,G8399);
  dff DFF_747(CK,G59451,G8400);
  dff DFF_748(CK,G59452,G8401);
  dff DFF_749(CK,G59453,G8402);
  dff DFF_750(CK,G59454,G8403);
  dff DFF_751(CK,G59455,G8404);
  dff DFF_752(CK,G59456,G8405);
  dff DFF_753(CK,G59457,G8406);
  dff DFF_754(CK,G59458,G8407);
  dff DFF_755(CK,G59459,G8408);
  dff DFF_756(CK,G59460,G8409);
  dff DFF_757(CK,G59461,G8410);
  dff DFF_758(CK,G59462,G8411);
  dff DFF_759(CK,G59463,G8412);
  dff DFF_760(CK,G59464,G8413);
  dff DFF_761(CK,G59465,G8414);
  dff DFF_762(CK,G59466,G8415);
  dff DFF_763(CK,G59467,G8416);
  dff DFF_764(CK,G59468,G8417);
  dff DFF_765(CK,G59469,G8418);
  dff DFF_766(CK,G59470,G8419);
  dff DFF_767(CK,G59471,G8420);
  dff DFF_768(CK,G59472,G8421);
  dff DFF_769(CK,G59473,G8422);
  dff DFF_770(CK,G59474,G8423);
  dff DFF_771(CK,G59475,G8424);
  dff DFF_772(CK,G59476,G8425);
  dff DFF_773(CK,G59477,G8426);
  dff DFF_774(CK,G59478,G8427);
  dff DFF_775(CK,G59479,G8428);
  dff DFF_776(CK,G59480,G8429);
  dff DFF_777(CK,G59481,G8430);
  dff DFF_778(CK,G59482,G8431);
  dff DFF_779(CK,G59483,G8432);
  dff DFF_780(CK,G59484,G8433);
  dff DFF_781(CK,G59485,G8434);
  dff DFF_782(CK,G59486,G8435);
  dff DFF_783(CK,G59487,G8436);
  dff DFF_784(CK,G59488,G8437);
  dff DFF_785(CK,G59489,G8438);
  dff DFF_786(CK,G59490,G8439);
  dff DFF_787(CK,G59491,G8440);
  dff DFF_788(CK,G59492,G8441);
  dff DFF_789(CK,G59493,G8442);
  dff DFF_790(CK,G59494,G8443);
  dff DFF_791(CK,G59495,G8444);
  dff DFF_792(CK,G59496,G8445);
  dff DFF_793(CK,G59497,G8446);
  dff DFF_794(CK,G59498,G8447);
  dff DFF_795(CK,G59499,G8448);
  dff DFF_796(CK,G59500,G8449);
  dff DFF_797(CK,G59501,G8450);
  dff DFF_798(CK,G59502,G8451);
  dff DFF_799(CK,G59503,G8452);
  dff DFF_800(CK,G59504,G8453);
  dff DFF_801(CK,G59505,G8454);
  dff DFF_802(CK,G59506,G8455);
  dff DFF_803(CK,G59507,G8456);
  dff DFF_804(CK,G59508,G8457);
  dff DFF_805(CK,G59509,G8458);
  dff DFF_806(CK,G59510,G8459);
  dff DFF_807(CK,G59511,G8460);
  dff DFF_808(CK,G59512,G8461);
  dff DFF_809(CK,G59513,G8462);
  dff DFF_810(CK,G59514,G8463);
  dff DFF_811(CK,G59515,G8464);
  dff DFF_812(CK,G59516,G8465);
  dff DFF_813(CK,G59517,G8466);
  dff DFF_814(CK,G59518,G8467);
  dff DFF_815(CK,G59519,G8468);
  dff DFF_816(CK,G59520,G8469);
  dff DFF_817(CK,G59521,G8470);
  dff DFF_818(CK,G59522,G8471);
  dff DFF_819(CK,G59523,G8472);
  dff DFF_820(CK,G59524,G8473);
  dff DFF_821(CK,G59525,G8474);
  dff DFF_822(CK,G59526,G8475);
  dff DFF_823(CK,G59527,G8476);
  dff DFF_824(CK,G59528,G8477);
  dff DFF_825(CK,G59529,G8478);
  dff DFF_826(CK,G59530,G8479);
  dff DFF_827(CK,G59531,G8480);
  dff DFF_828(CK,G59532,G8481);
  dff DFF_829(CK,G59533,G8482);
  dff DFF_830(CK,G59534,G8483);
  dff DFF_831(CK,G59535,G8484);
  dff DFF_832(CK,G59536,G8485);
  dff DFF_833(CK,G59537,G8486);
  dff DFF_834(CK,G59538,G8487);
  dff DFF_835(CK,G59539,G8488);
  dff DFF_836(CK,G59540,G8489);
  dff DFF_837(CK,G59541,G8490);
  dff DFF_838(CK,G59542,G8491);
  dff DFF_839(CK,G59543,G8492);
  dff DFF_840(CK,G59544,G8493);
  dff DFF_841(CK,G59545,G8494);
  dff DFF_842(CK,G59546,G8495);
  dff DFF_843(CK,G59547,G8496);
  dff DFF_844(CK,G59548,G8497);
  dff DFF_845(CK,G59549,G8498);
  dff DFF_846(CK,G59550,G8499);
  dff DFF_847(CK,G59551,G8500);
  dff DFF_848(CK,G59552,G8501);
  dff DFF_849(CK,G59553,G8502);
  dff DFF_850(CK,G59554,G8503);
  dff DFF_851(CK,G59555,G8504);
  dff DFF_852(CK,G59556,G8505);
  dff DFF_853(CK,G59557,G9267);
  dff DFF_854(CK,G59558,G9266);
  dff DFF_855(CK,G59559,G9265);
  dff DFF_856(CK,G59560,G9263);
  dff DFF_857(CK,G59561,G9262);
  dff DFF_858(CK,G59562,G8506);
  dff DFF_859(CK,G59563,G8507);
  dff DFF_860(CK,G59564,G8508);
  dff DFF_861(CK,G59565,G8509);
  dff DFF_862(CK,G59566,G8744);
  dff DFF_863(CK,G59567,G8510);
  dff DFF_864(CK,G59568,G8511);
  dff DFF_865(CK,G59569,G8512);
  dff DFF_866(CK,G59570,G8513);
  dff DFF_867(CK,G59571,G8514);
  dff DFF_868(CK,G59572,G8515);
  dff DFF_869(CK,G59573,G8516);
  dff DFF_870(CK,G59574,G8517);
  dff DFF_871(CK,G59575,G8518);
  dff DFF_872(CK,G59576,G8519);
  dff DFF_873(CK,G59577,G8520);
  dff DFF_874(CK,G59578,G8521);
  dff DFF_875(CK,G59579,G8522);
  dff DFF_876(CK,G59580,G8523);
  dff DFF_877(CK,G59581,G8524);
  dff DFF_878(CK,G59582,G8525);
  dff DFF_879(CK,G59583,G8526);
  dff DFF_880(CK,G59584,G8527);
  dff DFF_881(CK,G59585,G8528);
  dff DFF_882(CK,G59586,G8529);
  dff DFF_883(CK,G59587,G8530);
  dff DFF_884(CK,G59588,G8531);
  dff DFF_885(CK,G59589,G8532);
  dff DFF_886(CK,G59590,G8533);
  dff DFF_887(CK,G59591,G8534);
  dff DFF_888(CK,G59592,G8535);
  dff DFF_889(CK,G59593,G8536);
  dff DFF_890(CK,G59594,G8537);
  dff DFF_891(CK,G59595,G8538);
  dff DFF_892(CK,G59596,G8539);
  dff DFF_893(CK,G59597,G8540);
  dff DFF_894(CK,G59598,G8541);
  dff DFF_895(CK,G59599,G8542);
  dff DFF_896(CK,G59600,G8543);
  dff DFF_897(CK,G59601,G8544);
  dff DFF_898(CK,G59602,G8545);
  dff DFF_899(CK,G59603,G8546);
  dff DFF_900(CK,G59604,G8547);
  dff DFF_901(CK,G59605,G8548);
  dff DFF_902(CK,G59606,G8549);
  dff DFF_903(CK,G59607,G8550);
  dff DFF_904(CK,G59608,G8551);
  dff DFF_905(CK,G59609,G8552);
  dff DFF_906(CK,G59610,G8553);
  dff DFF_907(CK,G59611,G8554);
  dff DFF_908(CK,G59612,G8555);
  dff DFF_909(CK,G59613,G8556);
  dff DFF_910(CK,G59614,G8557);
  dff DFF_911(CK,G59615,G8558);
  dff DFF_912(CK,G59616,G8559);
  dff DFF_913(CK,G59617,G8560);
  dff DFF_914(CK,G59618,G8561);
  dff DFF_915(CK,G59619,G8562);
  dff DFF_916(CK,G59620,G8563);
  dff DFF_917(CK,G59621,G8564);
  dff DFF_918(CK,G59622,G8565);
  dff DFF_919(CK,G59623,G8566);
  dff DFF_920(CK,G59624,G8567);
  dff DFF_921(CK,G59625,G8568);
  dff DFF_922(CK,G59626,G8569);
  dff DFF_923(CK,G59627,G8570);
  dff DFF_924(CK,G59628,G8571);
  dff DFF_925(CK,G59629,G8572);
  dff DFF_926(CK,G59630,G8573);
  dff DFF_927(CK,G59631,G8574);
  dff DFF_928(CK,G59632,G8575);
  dff DFF_929(CK,G59633,G8576);
  dff DFF_930(CK,G59634,G8577);
  dff DFF_931(CK,G59635,G8578);
  dff DFF_932(CK,G59636,G8579);
  dff DFF_933(CK,G59637,G8580);
  dff DFF_934(CK,G59638,G8581);
  dff DFF_935(CK,G59639,G8582);
  dff DFF_936(CK,G59640,G8583);
  dff DFF_937(CK,G59641,G8584);
  dff DFF_938(CK,G59642,G8585);
  dff DFF_939(CK,G59643,G8586);
  dff DFF_940(CK,G59644,G8587);
  dff DFF_941(CK,G59645,G8588);
  dff DFF_942(CK,G59646,G8589);
  dff DFF_943(CK,G59647,G8590);
  dff DFF_944(CK,G59648,G8591);
  dff DFF_945(CK,G59649,G8592);
  dff DFF_946(CK,G59650,G8593);
  dff DFF_947(CK,G59651,G8594);
  dff DFF_948(CK,G59652,G8595);
  dff DFF_949(CK,G59653,G8596);
  dff DFF_950(CK,G59654,G8597);
  dff DFF_951(CK,G59655,G8598);
  dff DFF_952(CK,G59656,G8599);
  dff DFF_953(CK,G59657,G8600);
  dff DFF_954(CK,G59658,G8601);
  dff DFF_955(CK,G59659,G8602);
  dff DFF_956(CK,G59660,G8603);
  dff DFF_957(CK,G59661,G8604);
  dff DFF_958(CK,G59662,G8605);
  dff DFF_959(CK,G59663,G8606);
  dff DFF_960(CK,G59664,G8607);
  dff DFF_961(CK,G59665,G8608);
  dff DFF_962(CK,G59666,G8609);
  dff DFF_963(CK,G59667,G8610);
  dff DFF_964(CK,G59668,G8611);
  dff DFF_965(CK,G59669,G8612);
  dff DFF_966(CK,G59670,G8613);
  dff DFF_967(CK,G59671,G8614);
  dff DFF_968(CK,G59672,G8615);
  dff DFF_969(CK,G59673,G8616);
  dff DFF_970(CK,G59674,G8617);
  dff DFF_971(CK,G59675,G8618);
  dff DFF_972(CK,G59676,G8619);
  dff DFF_973(CK,G59677,G8620);
  dff DFF_974(CK,G59678,G8621);
  dff DFF_975(CK,G59679,G8622);
  dff DFF_976(CK,G59680,G8623);
  dff DFF_977(CK,G59681,G8624);
  dff DFF_978(CK,G59682,G8625);
  dff DFF_979(CK,G59683,G8626);
  dff DFF_980(CK,G59684,G8627);
  dff DFF_981(CK,G59685,G8628);
  dff DFF_982(CK,G59686,G8629);
  dff DFF_983(CK,G59687,G8630);
  dff DFF_984(CK,G59688,G8631);
  dff DFF_985(CK,G59689,G8632);
  dff DFF_986(CK,G59690,G8633);
  dff DFF_987(CK,G59691,G8634);
  dff DFF_988(CK,G59692,G8635);
  dff DFF_989(CK,G59693,G8636);
  dff DFF_990(CK,G59694,G8637);
  dff DFF_991(CK,G59695,G8638);
  dff DFF_992(CK,G59696,G8639);
  dff DFF_993(CK,G59697,G8640);
  dff DFF_994(CK,G59698,G8641);
  dff DFF_995(CK,G59699,G8642);
  dff DFF_996(CK,G59700,G8643);
  dff DFF_997(CK,G59701,G8644);
  dff DFF_998(CK,G59702,G8645);
  dff DFF_999(CK,G59703,G8646);
  dff DFF_1000(CK,G59704,G8647);
  dff DFF_1001(CK,G59705,G8648);
  dff DFF_1002(CK,G59706,G8649);
  dff DFF_1003(CK,G59707,G8650);
  dff DFF_1004(CK,G59708,G8651);
  dff DFF_1005(CK,G59709,G8652);
  dff DFF_1006(CK,G59710,G8653);
  dff DFF_1007(CK,G59711,G8654);
  dff DFF_1008(CK,G59712,G8655);
  dff DFF_1009(CK,G59713,G8656);
  dff DFF_1010(CK,G59714,G8657);
  dff DFF_1011(CK,G59715,G8658);
  dff DFF_1012(CK,G59716,G8659);
  dff DFF_1013(CK,G59717,G8660);
  dff DFF_1014(CK,G59718,G8661);
  dff DFF_1015(CK,G59719,G8662);
  dff DFF_1016(CK,G59720,G8663);
  dff DFF_1017(CK,G59721,G8664);
  dff DFF_1018(CK,G59722,G8665);
  dff DFF_1019(CK,G59723,G8666);
  dff DFF_1020(CK,G59724,G8667);
  dff DFF_1021(CK,G59725,G8668);
  dff DFF_1022(CK,G59726,G8669);
  dff DFF_1023(CK,G59727,G8670);
  dff DFF_1024(CK,G59728,G8671);
  dff DFF_1025(CK,G59729,G8672);
  dff DFF_1026(CK,G59730,G8673);
  dff DFF_1027(CK,G59731,G8674);
  dff DFF_1028(CK,G59732,G8675);
  dff DFF_1029(CK,G59733,G8676);
  dff DFF_1030(CK,G59734,G8677);
  dff DFF_1031(CK,G59735,G8678);
  dff DFF_1032(CK,G59736,G8679);
  dff DFF_1033(CK,G59737,G8680);
  dff DFF_1034(CK,G59738,G8681);
  dff DFF_1035(CK,G59739,G8682);
  dff DFF_1036(CK,G59740,G8683);
  dff DFF_1037(CK,G59741,G8684);
  dff DFF_1038(CK,G59742,G8685);
  dff DFF_1039(CK,G59743,G8686);
  dff DFF_1040(CK,G59744,G8687);
  dff DFF_1041(CK,G59745,G8688);
  dff DFF_1042(CK,G59746,G8689);
  dff DFF_1043(CK,G59747,G8690);
  dff DFF_1044(CK,G59748,G8691);
  dff DFF_1045(CK,G59749,G8692);
  dff DFF_1046(CK,G59750,G8693);
  dff DFF_1047(CK,G59751,G8694);
  dff DFF_1048(CK,G59752,G8695);
  dff DFF_1049(CK,G59753,G8696);
  dff DFF_1050(CK,G59754,G8697);
  dff DFF_1051(CK,G59755,G8698);
  dff DFF_1052(CK,G59756,G8699);
  dff DFF_1053(CK,G59757,G8700);
  dff DFF_1054(CK,G59758,G8701);
  dff DFF_1055(CK,G59759,G8702);
  dff DFF_1056(CK,G59760,G8703);
  dff DFF_1057(CK,G59761,G8704);
  dff DFF_1058(CK,G59762,G8705);
  dff DFF_1059(CK,G59763,G8706);
  dff DFF_1060(CK,G59764,G8707);
  dff DFF_1061(CK,G59765,G8708);
  dff DFF_1062(CK,G59766,G8709);
  dff DFF_1063(CK,G59767,G8710);
  dff DFF_1064(CK,G59768,G8711);
  dff DFF_1065(CK,G59769,G8712);
  dff DFF_1066(CK,G59770,G8713);
  dff DFF_1067(CK,G59771,G8714);
  dff DFF_1068(CK,G59772,G8715);
  dff DFF_1069(CK,G59773,G8716);
  dff DFF_1070(CK,G59774,G8717);
  dff DFF_1071(CK,G59775,G8718);
  dff DFF_1072(CK,G59776,G8719);
  dff DFF_1073(CK,G59777,G8720);
  dff DFF_1074(CK,G59778,G8721);
  dff DFF_1075(CK,G59779,G8722);
  dff DFF_1076(CK,G59780,G8723);
  dff DFF_1077(CK,G59781,G8724);
  dff DFF_1078(CK,G59782,G8725);
  dff DFF_1079(CK,G59783,G8726);
  dff DFF_1080(CK,G59784,G8727);
  dff DFF_1081(CK,G59785,G8728);
  dff DFF_1082(CK,G59786,G8729);
  dff DFF_1083(CK,G59787,G8730);
  dff DFF_1084(CK,G59788,G8731);
  dff DFF_1085(CK,G59789,G8732);
  dff DFF_1086(CK,G59790,G8733);
  dff DFF_1087(CK,G59791,G8734);
  dff DFF_1088(CK,G59792,G8735);
  dff DFF_1089(CK,G59793,G8736);
  dff DFF_1090(CK,G59794,G9261);
  dff DFF_1091(CK,G59795,G8737);
  dff DFF_1092(CK,G59796,G8738);
  dff DFF_1093(CK,G59797,G8739);
  dff DFF_1094(CK,G59798,G9260);
  dff DFF_1095(CK,G59799,G8740);
  dff DFF_1096(CK,G59800,G9259);
  dff DFF_1097(CK,G59801,G8741);
  dff DFF_1098(CK,G59802,G8742);
  dff DFF_1099(CK,G59803,G9258);
  dff DFF_1100(CK,G59804,G9257);
  dff DFF_1101(CK,G59805,G15270);
  dff DFF_1102(CK,G59806,G15269);
  dff DFF_1103(CK,G59807,G15268);
  dff DFF_1104(CK,G59808,G15267);
  dff DFF_1105(CK,G59809,G14308);
  dff DFF_1106(CK,G59810,G14309);
  dff DFF_1107(CK,G59811,G14310);
  dff DFF_1108(CK,G59812,G14311);
  dff DFF_1109(CK,G59813,G14312);
  dff DFF_1110(CK,G59814,G14313);
  dff DFF_1111(CK,G59815,G14314);
  dff DFF_1112(CK,G59816,G14315);
  dff DFF_1113(CK,G59817,G14316);
  dff DFF_1114(CK,G59818,G14317);
  dff DFF_1115(CK,G59819,G14318);
  dff DFF_1116(CK,G59820,G14319);
  dff DFF_1117(CK,G59821,G14320);
  dff DFF_1118(CK,G59822,G14321);
  dff DFF_1119(CK,G59823,G14322);
  dff DFF_1120(CK,G59824,G14323);
  dff DFF_1121(CK,G59825,G14324);
  dff DFF_1122(CK,G59826,G14325);
  dff DFF_1123(CK,G59827,G14326);
  dff DFF_1124(CK,G59828,G14327);
  dff DFF_1125(CK,G59829,G14328);
  dff DFF_1126(CK,G59830,G14329);
  dff DFF_1127(CK,G59831,G14330);
  dff DFF_1128(CK,G59832,G14331);
  dff DFF_1129(CK,G59833,G14332);
  dff DFF_1130(CK,G59834,G14333);
  dff DFF_1131(CK,G59835,G14334);
  dff DFF_1132(CK,G59836,G14335);
  dff DFF_1133(CK,G59837,G14336);
  dff DFF_1134(CK,G59838,G14337);
  dff DFF_1135(CK,G59839,G14338);
  dff DFF_1136(CK,G59840,G14339);
  dff DFF_1137(CK,G59841,G14340);
  dff DFF_1138(CK,G59842,G15266);
  dff DFF_1139(CK,G59843,G15265);
  dff DFF_1140(CK,G59844,G14341);
  dff DFF_1141(CK,G59845,G14342);
  dff DFF_1142(CK,G59846,G14343);
  dff DFF_1143(CK,G59847,G14344);
  dff DFF_1144(CK,G59848,G14345);
  dff DFF_1145(CK,G59849,G14346);
  dff DFF_1146(CK,G59850,G14347);
  dff DFF_1147(CK,G59851,G14348);
  dff DFF_1148(CK,G59852,G14349);
  dff DFF_1149(CK,G59853,G14350);
  dff DFF_1150(CK,G59854,G14351);
  dff DFF_1151(CK,G59855,G14352);
  dff DFF_1152(CK,G59856,G14353);
  dff DFF_1153(CK,G59857,G14354);
  dff DFF_1154(CK,G59858,G14355);
  dff DFF_1155(CK,G59859,G14356);
  dff DFF_1156(CK,G59860,G14357);
  dff DFF_1157(CK,G59861,G14358);
  dff DFF_1158(CK,G59862,G14359);
  dff DFF_1159(CK,G59863,G14360);
  dff DFF_1160(CK,G59864,G14361);
  dff DFF_1161(CK,G59865,G14362);
  dff DFF_1162(CK,G59866,G14363);
  dff DFF_1163(CK,G59867,G14364);
  dff DFF_1164(CK,G59868,G14365);
  dff DFF_1165(CK,G59869,G14366);
  dff DFF_1166(CK,G59870,G14367);
  dff DFF_1167(CK,G59871,G14368);
  dff DFF_1168(CK,G59872,G14369);
  dff DFF_1169(CK,G59873,G14370);
  dff DFF_1170(CK,G59874,G14371);
  dff DFF_1171(CK,G59875,G14372);
  dff DFF_1172(CK,G59876,G14373);
  dff DFF_1173(CK,G59877,G14374);
  dff DFF_1174(CK,G59878,G14375);
  dff DFF_1175(CK,G59879,G14376);
  dff DFF_1176(CK,G59880,G14377);
  dff DFF_1177(CK,G59881,G14378);
  dff DFF_1178(CK,G59882,G14379);
  dff DFF_1179(CK,G59883,G14380);
  dff DFF_1180(CK,G59884,G14381);
  dff DFF_1181(CK,G59885,G14382);
  dff DFF_1182(CK,G59886,G14383);
  dff DFF_1183(CK,G59887,G14384);
  dff DFF_1184(CK,G59888,G14385);
  dff DFF_1185(CK,G59889,G14386);
  dff DFF_1186(CK,G59890,G14387);
  dff DFF_1187(CK,G59891,G14388);
  dff DFF_1188(CK,G59892,G14389);
  dff DFF_1189(CK,G59893,G14390);
  dff DFF_1190(CK,G59894,G14391);
  dff DFF_1191(CK,G59895,G14392);
  dff DFF_1192(CK,G59896,G14393);
  dff DFF_1193(CK,G59897,G14394);
  dff DFF_1194(CK,G59898,G14395);
  dff DFF_1195(CK,G59899,G14396);
  dff DFF_1196(CK,G59900,G14397);
  dff DFF_1197(CK,G59901,G14398);
  dff DFF_1198(CK,G59902,G14399);
  dff DFF_1199(CK,G59903,G14400);
  dff DFF_1200(CK,G59904,G14401);
  dff DFF_1201(CK,G59905,G14402);
  dff DFF_1202(CK,G59906,G14403);
  dff DFF_1203(CK,G59907,G14404);
  dff DFF_1204(CK,G59908,G14405);
  dff DFF_1205(CK,G59909,G14406);
  dff DFF_1206(CK,G59910,G14407);
  dff DFF_1207(CK,G59911,G14408);
  dff DFF_1208(CK,G59912,G14409);
  dff DFF_1209(CK,G59913,G14410);
  dff DFF_1210(CK,G59914,G14411);
  dff DFF_1211(CK,G59915,G14412);
  dff DFF_1212(CK,G59916,G14413);
  dff DFF_1213(CK,G59917,G14414);
  dff DFF_1214(CK,G59918,G14415);
  dff DFF_1215(CK,G59919,G14416);
  dff DFF_1216(CK,G59920,G14417);
  dff DFF_1217(CK,G59921,G14418);
  dff DFF_1218(CK,G59922,G14419);
  dff DFF_1219(CK,G59923,G14420);
  dff DFF_1220(CK,G59924,G14421);
  dff DFF_1221(CK,G59925,G14422);
  dff DFF_1222(CK,G59926,G14423);
  dff DFF_1223(CK,G59927,G14424);
  dff DFF_1224(CK,G59928,G14425);
  dff DFF_1225(CK,G59929,G14426);
  dff DFF_1226(CK,G59930,G14427);
  dff DFF_1227(CK,G59931,G14428);
  dff DFF_1228(CK,G59932,G14429);
  dff DFF_1229(CK,G59933,G14430);
  dff DFF_1230(CK,G59934,G14431);
  dff DFF_1231(CK,G59935,G14432);
  dff DFF_1232(CK,G59936,G14433);
  dff DFF_1233(CK,G59937,G14434);
  dff DFF_1234(CK,G59938,G14435);
  dff DFF_1235(CK,G59939,G14436);
  dff DFF_1236(CK,G59940,G14437);
  dff DFF_1237(CK,G59941,G14438);
  dff DFF_1238(CK,G59942,G14439);
  dff DFF_1239(CK,G59943,G14440);
  dff DFF_1240(CK,G59944,G14441);
  dff DFF_1241(CK,G59945,G14442);
  dff DFF_1242(CK,G59946,G14443);
  dff DFF_1243(CK,G59947,G14444);
  dff DFF_1244(CK,G59948,G14445);
  dff DFF_1245(CK,G59949,G14446);
  dff DFF_1246(CK,G59950,G14447);
  dff DFF_1247(CK,G59951,G14448);
  dff DFF_1248(CK,G59952,G14449);
  dff DFF_1249(CK,G59953,G14450);
  dff DFF_1250(CK,G59954,G14451);
  dff DFF_1251(CK,G59955,G14452);
  dff DFF_1252(CK,G59956,G14453);
  dff DFF_1253(CK,G59957,G14454);
  dff DFF_1254(CK,G59958,G14455);
  dff DFF_1255(CK,G59959,G14456);
  dff DFF_1256(CK,G59960,G14457);
  dff DFF_1257(CK,G59961,G14458);
  dff DFF_1258(CK,G59962,G14459);
  dff DFF_1259(CK,G59963,G14460);
  dff DFF_1260(CK,G59964,G14461);
  dff DFF_1261(CK,G59965,G14462);
  dff DFF_1262(CK,G59966,G14463);
  dff DFF_1263(CK,G59967,G14464);
  dff DFF_1264(CK,G59968,G14465);
  dff DFF_1265(CK,G59969,G14466);
  dff DFF_1266(CK,G59970,G14467);
  dff DFF_1267(CK,G59971,G14468);
  dff DFF_1268(CK,G59972,G14469);
  dff DFF_1269(CK,G59973,G14470);
  dff DFF_1270(CK,G59974,G14471);
  dff DFF_1271(CK,G59975,G14472);
  dff DFF_1272(CK,G59976,G14473);
  dff DFF_1273(CK,G59977,G14474);
  dff DFF_1274(CK,G59978,G14475);
  dff DFF_1275(CK,G59979,G14476);
  dff DFF_1276(CK,G59980,G14477);
  dff DFF_1277(CK,G59981,G14478);
  dff DFF_1278(CK,G59982,G14479);
  dff DFF_1279(CK,G59983,G14480);
  dff DFF_1280(CK,G59984,G14481);
  dff DFF_1281(CK,G59985,G14482);
  dff DFF_1282(CK,G59986,G14483);
  dff DFF_1283(CK,G59987,G14484);
  dff DFF_1284(CK,G59988,G14485);
  dff DFF_1285(CK,G59989,G14486);
  dff DFF_1286(CK,G59990,G14487);
  dff DFF_1287(CK,G59991,G14488);
  dff DFF_1288(CK,G59992,G14489);
  dff DFF_1289(CK,G59993,G14490);
  dff DFF_1290(CK,G59994,G14491);
  dff DFF_1291(CK,G59995,G14492);
  dff DFF_1292(CK,G59996,G14493);
  dff DFF_1293(CK,G59997,G14494);
  dff DFF_1294(CK,G59998,G14495);
  dff DFF_1295(CK,G59999,G14496);
  dff DFF_1296(CK,G60000,G14497);
  dff DFF_1297(CK,G60001,G14498);
  dff DFF_1298(CK,G60002,G14499);
  dff DFF_1299(CK,G60003,G14500);
  dff DFF_1300(CK,G60004,G14501);
  dff DFF_1301(CK,G60005,G14502);
  dff DFF_1302(CK,G60006,G15264);
  dff DFF_1303(CK,G60007,G15263);
  dff DFF_1304(CK,G60008,G15262);
  dff DFF_1305(CK,G60009,G15260);
  dff DFF_1306(CK,G60010,G15259);
  dff DFF_1307(CK,G60011,G14503);
  dff DFF_1308(CK,G60012,G14504);
  dff DFF_1309(CK,G60013,G14505);
  dff DFF_1310(CK,G60014,G14506);
  dff DFF_1311(CK,G60015,G14741);
  dff DFF_1312(CK,G60016,G14507);
  dff DFF_1313(CK,G60017,G14508);
  dff DFF_1314(CK,G60018,G14509);
  dff DFF_1315(CK,G60019,G14510);
  dff DFF_1316(CK,G60020,G14511);
  dff DFF_1317(CK,G60021,G14512);
  dff DFF_1318(CK,G60022,G14513);
  dff DFF_1319(CK,G60023,G14514);
  dff DFF_1320(CK,G60024,G14515);
  dff DFF_1321(CK,G60025,G14516);
  dff DFF_1322(CK,G60026,G14517);
  dff DFF_1323(CK,G60027,G14518);
  dff DFF_1324(CK,G60028,G14519);
  dff DFF_1325(CK,G60029,G14520);
  dff DFF_1326(CK,G60030,G14521);
  dff DFF_1327(CK,G60031,G14522);
  dff DFF_1328(CK,G60032,G14523);
  dff DFF_1329(CK,G60033,G14524);
  dff DFF_1330(CK,G60034,G14525);
  dff DFF_1331(CK,G60035,G14526);
  dff DFF_1332(CK,G60036,G14527);
  dff DFF_1333(CK,G60037,G14528);
  dff DFF_1334(CK,G60038,G14529);
  dff DFF_1335(CK,G60039,G14530);
  dff DFF_1336(CK,G60040,G14531);
  dff DFF_1337(CK,G60041,G14532);
  dff DFF_1338(CK,G60042,G14533);
  dff DFF_1339(CK,G60043,G14534);
  dff DFF_1340(CK,G60044,G14535);
  dff DFF_1341(CK,G60045,G14536);
  dff DFF_1342(CK,G60046,G14537);
  dff DFF_1343(CK,G60047,G14538);
  dff DFF_1344(CK,G60048,G14539);
  dff DFF_1345(CK,G60049,G14540);
  dff DFF_1346(CK,G60050,G14541);
  dff DFF_1347(CK,G60051,G14542);
  dff DFF_1348(CK,G60052,G14543);
  dff DFF_1349(CK,G60053,G14544);
  dff DFF_1350(CK,G60054,G14545);
  dff DFF_1351(CK,G60055,G14546);
  dff DFF_1352(CK,G60056,G14547);
  dff DFF_1353(CK,G60057,G14548);
  dff DFF_1354(CK,G60058,G14549);
  dff DFF_1355(CK,G60059,G14550);
  dff DFF_1356(CK,G60060,G14551);
  dff DFF_1357(CK,G60061,G14552);
  dff DFF_1358(CK,G60062,G14553);
  dff DFF_1359(CK,G60063,G14554);
  dff DFF_1360(CK,G60064,G14555);
  dff DFF_1361(CK,G60065,G14556);
  dff DFF_1362(CK,G60066,G14557);
  dff DFF_1363(CK,G60067,G14558);
  dff DFF_1364(CK,G60068,G14559);
  dff DFF_1365(CK,G60069,G14560);
  dff DFF_1366(CK,G60070,G14561);
  dff DFF_1367(CK,G60071,G14562);
  dff DFF_1368(CK,G60072,G14563);
  dff DFF_1369(CK,G60073,G14564);
  dff DFF_1370(CK,G60074,G14565);
  dff DFF_1371(CK,G60075,G14566);
  dff DFF_1372(CK,G60076,G14567);
  dff DFF_1373(CK,G60077,G14568);
  dff DFF_1374(CK,G60078,G14569);
  dff DFF_1375(CK,G60079,G14570);
  dff DFF_1376(CK,G60080,G14571);
  dff DFF_1377(CK,G60081,G14572);
  dff DFF_1378(CK,G60082,G14573);
  dff DFF_1379(CK,G60083,G14574);
  dff DFF_1380(CK,G60084,G14575);
  dff DFF_1381(CK,G60085,G14576);
  dff DFF_1382(CK,G60086,G14577);
  dff DFF_1383(CK,G60087,G14578);
  dff DFF_1384(CK,G60088,G14579);
  dff DFF_1385(CK,G60089,G14580);
  dff DFF_1386(CK,G60090,G14581);
  dff DFF_1387(CK,G60091,G14582);
  dff DFF_1388(CK,G60092,G14583);
  dff DFF_1389(CK,G60093,G14584);
  dff DFF_1390(CK,G60094,G14585);
  dff DFF_1391(CK,G60095,G14586);
  dff DFF_1392(CK,G60096,G14587);
  dff DFF_1393(CK,G60097,G14588);
  dff DFF_1394(CK,G60098,G14589);
  dff DFF_1395(CK,G60099,G14590);
  dff DFF_1396(CK,G60100,G14591);
  dff DFF_1397(CK,G60101,G14592);
  dff DFF_1398(CK,G60102,G14593);
  dff DFF_1399(CK,G60103,G14594);
  dff DFF_1400(CK,G60104,G14595);
  dff DFF_1401(CK,G60105,G14596);
  dff DFF_1402(CK,G60106,G14597);
  dff DFF_1403(CK,G60107,G14598);
  dff DFF_1404(CK,G60108,G14599);
  dff DFF_1405(CK,G60109,G14600);
  dff DFF_1406(CK,G60110,G14601);
  dff DFF_1407(CK,G60111,G14602);
  dff DFF_1408(CK,G60112,G14603);
  dff DFF_1409(CK,G60113,G14604);
  dff DFF_1410(CK,G60114,G14605);
  dff DFF_1411(CK,G60115,G14606);
  dff DFF_1412(CK,G60116,G14607);
  dff DFF_1413(CK,G60117,G14608);
  dff DFF_1414(CK,G60118,G14609);
  dff DFF_1415(CK,G60119,G14610);
  dff DFF_1416(CK,G60120,G14611);
  dff DFF_1417(CK,G60121,G14612);
  dff DFF_1418(CK,G60122,G14613);
  dff DFF_1419(CK,G60123,G14614);
  dff DFF_1420(CK,G60124,G14615);
  dff DFF_1421(CK,G60125,G14616);
  dff DFF_1422(CK,G60126,G14617);
  dff DFF_1423(CK,G60127,G14618);
  dff DFF_1424(CK,G60128,G14619);
  dff DFF_1425(CK,G60129,G14620);
  dff DFF_1426(CK,G60130,G14621);
  dff DFF_1427(CK,G60131,G14622);
  dff DFF_1428(CK,G60132,G14623);
  dff DFF_1429(CK,G60133,G14624);
  dff DFF_1430(CK,G60134,G14625);
  dff DFF_1431(CK,G60135,G14626);
  dff DFF_1432(CK,G60136,G14627);
  dff DFF_1433(CK,G60137,G14628);
  dff DFF_1434(CK,G60138,G14629);
  dff DFF_1435(CK,G60139,G14630);
  dff DFF_1436(CK,G60140,G14631);
  dff DFF_1437(CK,G60141,G14632);
  dff DFF_1438(CK,G60142,G14633);
  dff DFF_1439(CK,G60143,G14634);
  dff DFF_1440(CK,G60144,G14635);
  dff DFF_1441(CK,G60145,G14636);
  dff DFF_1442(CK,G60146,G14637);
  dff DFF_1443(CK,G60147,G14638);
  dff DFF_1444(CK,G60148,G14639);
  dff DFF_1445(CK,G60149,G14640);
  dff DFF_1446(CK,G60150,G14641);
  dff DFF_1447(CK,G60151,G14642);
  dff DFF_1448(CK,G60152,G14643);
  dff DFF_1449(CK,G60153,G14644);
  dff DFF_1450(CK,G60154,G14645);
  dff DFF_1451(CK,G60155,G14646);
  dff DFF_1452(CK,G60156,G14647);
  dff DFF_1453(CK,G60157,G14648);
  dff DFF_1454(CK,G60158,G14649);
  dff DFF_1455(CK,G60159,G14650);
  dff DFF_1456(CK,G60160,G14651);
  dff DFF_1457(CK,G60161,G14652);
  dff DFF_1458(CK,G60162,G14653);
  dff DFF_1459(CK,G60163,G14654);
  dff DFF_1460(CK,G60164,G14655);
  dff DFF_1461(CK,G60165,G14656);
  dff DFF_1462(CK,G60166,G14657);
  dff DFF_1463(CK,G60167,G14658);
  dff DFF_1464(CK,G60168,G14659);
  dff DFF_1465(CK,G60169,G14660);
  dff DFF_1466(CK,G60170,G14661);
  dff DFF_1467(CK,G60171,G14662);
  dff DFF_1468(CK,G60172,G14663);
  dff DFF_1469(CK,G60173,G14664);
  dff DFF_1470(CK,G60174,G14665);
  dff DFF_1471(CK,G60175,G14666);
  dff DFF_1472(CK,G60176,G14667);
  dff DFF_1473(CK,G60177,G14668);
  dff DFF_1474(CK,G60178,G14669);
  dff DFF_1475(CK,G60179,G14670);
  dff DFF_1476(CK,G60180,G14671);
  dff DFF_1477(CK,G60181,G14672);
  dff DFF_1478(CK,G60182,G14673);
  dff DFF_1479(CK,G60183,G14674);
  dff DFF_1480(CK,G60184,G14675);
  dff DFF_1481(CK,G60185,G14676);
  dff DFF_1482(CK,G60186,G14677);
  dff DFF_1483(CK,G60187,G14678);
  dff DFF_1484(CK,G60188,G14679);
  dff DFF_1485(CK,G60189,G14680);
  dff DFF_1486(CK,G60190,G14681);
  dff DFF_1487(CK,G60191,G14682);
  dff DFF_1488(CK,G60192,G14683);
  dff DFF_1489(CK,G60193,G14684);
  dff DFF_1490(CK,G60194,G14685);
  dff DFF_1491(CK,G60195,G14686);
  dff DFF_1492(CK,G60196,G14687);
  dff DFF_1493(CK,G60197,G14688);
  dff DFF_1494(CK,G60198,G14689);
  dff DFF_1495(CK,G60199,G14690);
  dff DFF_1496(CK,G60200,G14691);
  dff DFF_1497(CK,G60201,G14692);
  dff DFF_1498(CK,G60202,G14693);
  dff DFF_1499(CK,G60203,G14694);
  dff DFF_1500(CK,G60204,G14695);
  dff DFF_1501(CK,G60205,G14696);
  dff DFF_1502(CK,G60206,G14697);
  dff DFF_1503(CK,G60207,G14698);
  dff DFF_1504(CK,G60208,G14699);
  dff DFF_1505(CK,G60209,G14700);
  dff DFF_1506(CK,G60210,G14701);
  dff DFF_1507(CK,G60211,G14702);
  dff DFF_1508(CK,G60212,G14703);
  dff DFF_1509(CK,G60213,G14704);
  dff DFF_1510(CK,G60214,G14705);
  dff DFF_1511(CK,G60215,G14706);
  dff DFF_1512(CK,G60216,G14707);
  dff DFF_1513(CK,G60217,G14708);
  dff DFF_1514(CK,G60218,G14709);
  dff DFF_1515(CK,G60219,G14710);
  dff DFF_1516(CK,G60220,G14711);
  dff DFF_1517(CK,G60221,G14712);
  dff DFF_1518(CK,G60222,G14713);
  dff DFF_1519(CK,G60223,G14714);
  dff DFF_1520(CK,G60224,G14715);
  dff DFF_1521(CK,G60225,G14716);
  dff DFF_1522(CK,G60226,G14717);
  dff DFF_1523(CK,G60227,G14718);
  dff DFF_1524(CK,G60228,G14719);
  dff DFF_1525(CK,G60229,G14720);
  dff DFF_1526(CK,G60230,G14721);
  dff DFF_1527(CK,G60231,G14722);
  dff DFF_1528(CK,G60232,G14723);
  dff DFF_1529(CK,G60233,G14724);
  dff DFF_1530(CK,G60234,G14725);
  dff DFF_1531(CK,G60235,G14726);
  dff DFF_1532(CK,G60236,G14727);
  dff DFF_1533(CK,G60237,G14728);
  dff DFF_1534(CK,G60238,G14729);
  dff DFF_1535(CK,G60239,G14730);
  dff DFF_1536(CK,G60240,G14731);
  dff DFF_1537(CK,G60241,G14732);
  dff DFF_1538(CK,G60242,G14733);
  dff DFF_1539(CK,G60243,G15258);
  dff DFF_1540(CK,G60244,G14734);
  dff DFF_1541(CK,G60245,G14735);
  dff DFF_1542(CK,G60246,G14736);
  dff DFF_1543(CK,G60247,G15257);
  dff DFF_1544(CK,G60248,G14737);
  dff DFF_1545(CK,G60249,G15256);
  dff DFF_1546(CK,G60250,G14738);
  dff DFF_1547(CK,G60251,G14739);
  dff DFF_1548(CK,G60252,G15255);
  dff DFF_1549(CK,G60253,G15254);
  not GNAME1550(G1550,G15276);
  not GNAME1551(G1551,G15275);
  nand GNAME1552(G1552,G20096,G1730,G1591);
  nand GNAME1553(G1553,G1724,G1725,G1731,G59351);
  nor GNAME1554(G1554,G1726,G1727,G1592,G60251);
  and GNAME1555(G1555,G1591,G20083);
  nand GNAME1556(G1556,G1735,G1733,G1734);
  nand GNAME1557(G1557,G1738,G1736,G1737);
  nand GNAME1558(G1558,G1741,G1739,G1740);
  nand GNAME1559(G1559,G1744,G1742,G1743);
  nand GNAME1560(G1560,G1747,G1745,G1746);
  nand GNAME1561(G1561,G1750,G1748,G1749);
  nand GNAME1562(G1562,G1753,G1751,G1752);
  nand GNAME1563(G1563,G1756,G1754,G1755);
  nand GNAME1564(G1564,G1759,G1757,G1758);
  nand GNAME1565(G1565,G1762,G1760,G1761);
  nand GNAME1566(G1566,G1765,G1763,G1764);
  nand GNAME1567(G1567,G1768,G1766,G1767);
  nand GNAME1568(G1568,G1771,G1769,G1770);
  nand GNAME1569(G1569,G1774,G1772,G1773);
  nand GNAME1570(G1570,G1777,G1775,G1776);
  nand GNAME1571(G1571,G1780,G1778,G1779);
  nand GNAME1572(G1572,G1783,G1781,G1782);
  nand GNAME1573(G1573,G1786,G1784,G1785);
  nand GNAME1574(G1574,G1789,G1787,G1788);
  nand GNAME1575(G1575,G1792,G1790,G1791);
  nand GNAME1576(G1576,G1795,G1793,G1794);
  nand GNAME1577(G1577,G1798,G1796,G1797);
  nand GNAME1578(G1578,G1801,G1799,G1800);
  nand GNAME1579(G1579,G1804,G1802,G1803);
  nand GNAME1580(G1580,G1807,G1805,G1806);
  nand GNAME1581(G1581,G1810,G1808,G1809);
  nand GNAME1582(G1582,G1813,G1811,G1812);
  nand GNAME1583(G1583,G1816,G1814,G1815);
  nand GNAME1584(G1584,G1819,G1817,G1818);
  nand GNAME1585(G1585,G1822,G1820,G1821);
  nand GNAME1586(G1586,G1825,G1823,G1824);
  nand GNAME1587(G1587,G1828,G1826,G1827);
  and GNAME1588(G1588,G58904,G58903);
  and GNAME1589(G1589,G36,G58906);
  and GNAME1590(G1590,G37,G58905);
  and GNAME1591(G1591,G1722,G1723,G59800,G59794);
  not GNAME1592(G1592,G20086);
  not GNAME1593(G1593,G20096);
  nor GNAME1594(G1594,G1554,G1595);
  and GNAME1595(G1595,G1732,G1730);
  nand GNAME1596(G1596,G1829,G1830);
  nand GNAME1597(G1597,G1831,G1832);
  nand GNAME1598(G1598,G1833,G1834);
  nand GNAME1599(G1599,G1835,G1836);
  nand GNAME1600(G1600,G1837,G1838);
  nand GNAME1601(G1601,G1839,G1840);
  nand GNAME1602(G1602,G1841,G1842);
  nand GNAME1603(G1603,G1843,G1844);
  nand GNAME1604(G1604,G1845,G1846);
  nand GNAME1605(G1605,G1847,G1848);
  nand GNAME1606(G1606,G1849,G1850);
  nand GNAME1607(G1607,G1851,G1852);
  nand GNAME1608(G1608,G1853,G1854);
  nand GNAME1609(G1609,G1855,G1856);
  nand GNAME1610(G1610,G1857,G1858);
  nand GNAME1611(G1611,G1859,G1860);
  nand GNAME1612(G1612,G1861,G1862);
  nand GNAME1613(G1613,G1863,G1864);
  nand GNAME1614(G1614,G1865,G1866);
  nand GNAME1615(G1615,G1867,G1868);
  nand GNAME1616(G1616,G1869,G1870);
  nand GNAME1617(G1617,G1871,G1872);
  nand GNAME1618(G1618,G1873,G1874);
  nand GNAME1619(G1619,G1875,G1876);
  nand GNAME1620(G1620,G1877,G1878);
  nand GNAME1621(G1621,G1879,G1880);
  nand GNAME1622(G1622,G1881,G1882);
  nand GNAME1623(G1623,G1883,G1884);
  nand GNAME1624(G1624,G1885,G1886);
  nand GNAME1625(G1625,G1887,G1888);
  nand GNAME1626(G1626,G1889,G1890);
  nand GNAME1627(G1627,G1891,G1892);
  nand GNAME1628(G1628,G1893,G1894);
  nand GNAME1629(G1629,G1895,G1896);
  nand GNAME1630(G1630,G1897,G1898);
  nand GNAME1631(G1631,G1899,G1900);
  nand GNAME1632(G1632,G1901,G1902);
  nand GNAME1633(G1633,G1903,G1904);
  nand GNAME1634(G1634,G1905,G1906);
  nand GNAME1635(G1635,G1907,G1908);
  nand GNAME1636(G1636,G1909,G1910);
  nand GNAME1637(G1637,G1911,G1912);
  nand GNAME1638(G1638,G1913,G1914);
  nand GNAME1639(G1639,G1915,G1916);
  nand GNAME1640(G1640,G1917,G1918);
  nand GNAME1641(G1641,G1919,G1920);
  nand GNAME1642(G1642,G1921,G1922);
  nand GNAME1643(G1643,G1923,G1924);
  nand GNAME1644(G1644,G1925,G1926);
  nand GNAME1645(G1645,G1927,G1928);
  nand GNAME1646(G1646,G1929,G1930);
  nand GNAME1647(G1647,G1931,G1932);
  nand GNAME1648(G1648,G1933,G1934);
  nand GNAME1649(G1649,G1935,G1936);
  nand GNAME1650(G1650,G1937,G1938);
  nand GNAME1651(G1651,G1939,G1940);
  nand GNAME1652(G1652,G1941,G1942);
  nand GNAME1653(G1653,G1943,G1944);
  nand GNAME1654(G1654,G1945,G1946);
  nand GNAME1655(G1655,G1947,G1948);
  nand GNAME1656(G1656,G1949,G1950);
  nand GNAME1657(G1657,G1951,G1952);
  nand GNAME1658(G1658,G1953,G1954);
  nand GNAME1659(G1659,G1955,G1956);
  nand GNAME1660(G1660,G1957,G1958);
  nand GNAME1661(G1661,G1959,G1960);
  nand GNAME1662(G1662,G1961,G1962);
  nand GNAME1663(G1663,G1963,G1964);
  nand GNAME1664(G1664,G1965,G1966);
  nand GNAME1665(G1665,G1967,G1968);
  nand GNAME1666(G1666,G1969,G1970);
  nand GNAME1667(G1667,G1971,G1972);
  nand GNAME1668(G1668,G1973,G1974);
  nand GNAME1669(G1669,G1975,G1976);
  nand GNAME1670(G1670,G1977,G1978);
  nand GNAME1671(G1671,G1979,G1980);
  nand GNAME1672(G1672,G1981,G1982);
  nand GNAME1673(G1673,G1983,G1984);
  nand GNAME1674(G1674,G1985,G1986);
  nand GNAME1675(G1675,G1987,G1988);
  nand GNAME1676(G1676,G1989,G1990);
  nand GNAME1677(G1677,G1991,G1992);
  nand GNAME1678(G1678,G1993,G1994);
  nand GNAME1679(G1679,G1995,G1996);
  nand GNAME1680(G1680,G1997,G1998);
  nand GNAME1681(G1681,G1999,G2000);
  nand GNAME1682(G1682,G2001,G2002);
  nand GNAME1683(G1683,G2003,G2004);
  nand GNAME1684(G1684,G2005,G2006);
  nand GNAME1685(G1685,G2007,G2008);
  nand GNAME1686(G1686,G2009,G2010);
  nand GNAME1687(G1687,G2011,G2012);
  nand GNAME1688(G1688,G2013,G2014);
  nand GNAME1689(G1689,G2015,G2016);
  nand GNAME1690(G1690,G2017,G2018);
  nand GNAME1691(G1691,G2019,G2020);
  nand GNAME1692(G1692,G2021,G2022);
  nand GNAME1693(G1693,G2023,G2024);
  nand GNAME1694(G1694,G2025,G2026);
  nand GNAME1695(G1695,G2027,G2028);
  nand GNAME1696(G1696,G2029,G2030);
  nand GNAME1697(G1697,G2031,G2032);
  nand GNAME1698(G1698,G2033,G2034);
  nand GNAME1699(G1699,G2035,G2036);
  nand GNAME1700(G1700,G2037,G2038);
  nand GNAME1701(G1701,G2039,G2040);
  nand GNAME1702(G1702,G2041,G2042);
  nand GNAME1703(G1703,G2043,G2044);
  nand GNAME1704(G1704,G2045,G2046);
  nand GNAME1705(G1705,G2047,G2048);
  nand GNAME1706(G1706,G2049,G2050);
  nand GNAME1707(G1707,G2051,G2052);
  nand GNAME1708(G1708,G2053,G2054);
  nand GNAME1709(G1709,G2055,G2056);
  nand GNAME1710(G1710,G2057,G2058);
  nand GNAME1711(G1711,G2059,G2060);
  nand GNAME1712(G1712,G2061,G2062);
  nand GNAME1713(G1713,G2063,G2064);
  nand GNAME1714(G1714,G2065,G2066);
  nand GNAME1715(G1715,G2067,G2068);
  nand GNAME1716(G1716,G2069,G2070);
  nand GNAME1717(G1717,G2071,G2072);
  nand GNAME1718(G1718,G2073,G2074);
  nand GNAME1719(G1719,G2075,G2076);
  nand GNAME1720(G1720,G2077,G2078);
  nand GNAME1721(G1721,G2079,G2080);
  nor GNAME1722(G1722,G59358,G59357,G59356,G59799);
  nor GNAME1723(G1723,G59802,G59359);
  nor GNAME1724(G1724,G58908,G58907,G58909,G59345,G58910);
  nor GNAME1725(G1725,G59350,G59353);
  or GNAME1726(G1726,G60248,G59808,G59807,G59806,G59805);
  nand GNAME1727(G1727,G60249,G60243);
  and GNAME1728(G1728,G20106,G20081,G20084);
  not GNAME1729(G1729,G1728);
  not GNAME1730(G1730,G1554);
  not GNAME1731(G1731,G1555);
  nand GNAME1732(G1732,G1591,G20096);
  nand GNAME1733(G1733,G1594,G59662);
  nand GNAME1734(G1734,G1554,G60111);
  nand GNAME1735(G1735,G1595,G58839);
  nand GNAME1736(G1736,G1594,G59663);
  nand GNAME1737(G1737,G1554,G60112);
  nand GNAME1738(G1738,G1595,G58840);
  nand GNAME1739(G1739,G1594,G59664);
  nand GNAME1740(G1740,G1554,G60113);
  nand GNAME1741(G1741,G1595,G58841);
  nand GNAME1742(G1742,G1594,G59665);
  nand GNAME1743(G1743,G1554,G60114);
  nand GNAME1744(G1744,G1595,G58842);
  nand GNAME1745(G1745,G1594,G59666);
  nand GNAME1746(G1746,G1554,G60115);
  nand GNAME1747(G1747,G1595,G58843);
  nand GNAME1748(G1748,G1594,G59667);
  nand GNAME1749(G1749,G1554,G60116);
  nand GNAME1750(G1750,G1595,G58844);
  nand GNAME1751(G1751,G1594,G59668);
  nand GNAME1752(G1752,G1554,G60117);
  nand GNAME1753(G1753,G1595,G58845);
  nand GNAME1754(G1754,G1594,G59669);
  nand GNAME1755(G1755,G1554,G60118);
  nand GNAME1756(G1756,G1595,G58846);
  nand GNAME1757(G1757,G1594,G59670);
  nand GNAME1758(G1758,G1554,G60119);
  nand GNAME1759(G1759,G1595,G58847);
  nand GNAME1760(G1760,G1594,G59671);
  nand GNAME1761(G1761,G1554,G60120);
  nand GNAME1762(G1762,G1595,G58848);
  nand GNAME1763(G1763,G1594,G59672);
  nand GNAME1764(G1764,G1554,G60121);
  nand GNAME1765(G1765,G1595,G58849);
  nand GNAME1766(G1766,G1594,G59673);
  nand GNAME1767(G1767,G1554,G60122);
  nand GNAME1768(G1768,G1595,G58850);
  nand GNAME1769(G1769,G1594,G59674);
  nand GNAME1770(G1770,G1554,G60123);
  nand GNAME1771(G1771,G1595,G58851);
  nand GNAME1772(G1772,G1594,G59675);
  nand GNAME1773(G1773,G1554,G60124);
  nand GNAME1774(G1774,G1595,G58852);
  nand GNAME1775(G1775,G1594,G59676);
  nand GNAME1776(G1776,G1554,G60125);
  nand GNAME1777(G1777,G1595,G58853);
  nand GNAME1778(G1778,G1594,G59677);
  nand GNAME1779(G1779,G1554,G60126);
  nand GNAME1780(G1780,G1595,G58854);
  nand GNAME1781(G1781,G1594,G59678);
  nand GNAME1782(G1782,G1554,G60127);
  nand GNAME1783(G1783,G1595,G58855);
  nand GNAME1784(G1784,G1594,G59679);
  nand GNAME1785(G1785,G1554,G60128);
  nand GNAME1786(G1786,G1595,G58856);
  nand GNAME1787(G1787,G1594,G59680);
  nand GNAME1788(G1788,G1554,G60129);
  nand GNAME1789(G1789,G1595,G58857);
  nand GNAME1790(G1790,G1594,G59681);
  nand GNAME1791(G1791,G1554,G60130);
  nand GNAME1792(G1792,G1595,G58858);
  nand GNAME1793(G1793,G1594,G59682);
  nand GNAME1794(G1794,G1554,G60131);
  nand GNAME1795(G1795,G1595,G58859);
  nand GNAME1796(G1796,G1594,G59683);
  nand GNAME1797(G1797,G1554,G60132);
  nand GNAME1798(G1798,G1595,G58860);
  nand GNAME1799(G1799,G1594,G59684);
  nand GNAME1800(G1800,G1554,G60133);
  nand GNAME1801(G1801,G1595,G58861);
  nand GNAME1802(G1802,G1594,G59685);
  nand GNAME1803(G1803,G1554,G60134);
  nand GNAME1804(G1804,G1595,G58862);
  nand GNAME1805(G1805,G1594,G59686);
  nand GNAME1806(G1806,G1554,G60135);
  nand GNAME1807(G1807,G1595,G58863);
  nand GNAME1808(G1808,G1594,G59687);
  nand GNAME1809(G1809,G1554,G60136);
  nand GNAME1810(G1810,G1595,G58864);
  nand GNAME1811(G1811,G1594,G59688);
  nand GNAME1812(G1812,G1554,G60137);
  nand GNAME1813(G1813,G1595,G58865);
  nand GNAME1814(G1814,G1594,G59689);
  nand GNAME1815(G1815,G1554,G60138);
  nand GNAME1816(G1816,G1595,G58866);
  nand GNAME1817(G1817,G1594,G59690);
  nand GNAME1818(G1818,G1554,G60139);
  nand GNAME1819(G1819,G1595,G58867);
  nand GNAME1820(G1820,G1594,G59691);
  nand GNAME1821(G1821,G1554,G60140);
  nand GNAME1822(G1822,G1595,G58868);
  nand GNAME1823(G1823,G1594,G59692);
  nand GNAME1824(G1824,G1554,G60141);
  nand GNAME1825(G1825,G1595,G58869);
  nand GNAME1826(G1826,G1594,G59693);
  nand GNAME1827(G1827,G1554,G60142);
  nand GNAME1828(G1828,G1595,G58870);
  nand GNAME1829(G1829,G1731,G58871);
  nand GNAME1830(G1830,G1555,G59662);
  nand GNAME1831(G1831,G1731,G58872);
  nand GNAME1832(G1832,G1555,G59663);
  nand GNAME1833(G1833,G1731,G58873);
  nand GNAME1834(G1834,G1555,G59664);
  nand GNAME1835(G1835,G1731,G58874);
  nand GNAME1836(G1836,G1555,G59665);
  nand GNAME1837(G1837,G1731,G58875);
  nand GNAME1838(G1838,G1555,G59666);
  nand GNAME1839(G1839,G1731,G58876);
  nand GNAME1840(G1840,G1555,G59667);
  nand GNAME1841(G1841,G1731,G58877);
  nand GNAME1842(G1842,G1555,G59668);
  nand GNAME1843(G1843,G1731,G58878);
  nand GNAME1844(G1844,G1555,G59669);
  nand GNAME1845(G1845,G1731,G58879);
  nand GNAME1846(G1846,G1555,G59670);
  nand GNAME1847(G1847,G1731,G58880);
  nand GNAME1848(G1848,G1555,G59671);
  nand GNAME1849(G1849,G1731,G58881);
  nand GNAME1850(G1850,G1555,G59672);
  nand GNAME1851(G1851,G1731,G58882);
  nand GNAME1852(G1852,G1555,G59673);
  nand GNAME1853(G1853,G1731,G58883);
  nand GNAME1854(G1854,G1555,G59674);
  nand GNAME1855(G1855,G1731,G58884);
  nand GNAME1856(G1856,G1555,G59675);
  nand GNAME1857(G1857,G1731,G58885);
  nand GNAME1858(G1858,G1555,G59676);
  nand GNAME1859(G1859,G1731,G58886);
  nand GNAME1860(G1860,G1555,G59677);
  nand GNAME1861(G1861,G1731,G58887);
  nand GNAME1862(G1862,G1555,G59678);
  nand GNAME1863(G1863,G1731,G58888);
  nand GNAME1864(G1864,G1555,G59679);
  nand GNAME1865(G1865,G1731,G58889);
  nand GNAME1866(G1866,G1555,G59680);
  nand GNAME1867(G1867,G1731,G58890);
  nand GNAME1868(G1868,G1555,G59681);
  nand GNAME1869(G1869,G1731,G58891);
  nand GNAME1870(G1870,G1555,G59682);
  nand GNAME1871(G1871,G1731,G58892);
  nand GNAME1872(G1872,G1555,G59683);
  nand GNAME1873(G1873,G1731,G58893);
  nand GNAME1874(G1874,G1555,G59684);
  nand GNAME1875(G1875,G1731,G58894);
  nand GNAME1876(G1876,G1555,G59685);
  nand GNAME1877(G1877,G1731,G58895);
  nand GNAME1878(G1878,G1555,G59686);
  nand GNAME1879(G1879,G1731,G58896);
  nand GNAME1880(G1880,G1555,G59687);
  nand GNAME1881(G1881,G1731,G58897);
  nand GNAME1882(G1882,G1555,G59688);
  nand GNAME1883(G1883,G1731,G58898);
  nand GNAME1884(G1884,G1555,G59689);
  nand GNAME1885(G1885,G1731,G58899);
  nand GNAME1886(G1886,G1555,G59690);
  nand GNAME1887(G1887,G1731,G58900);
  nand GNAME1888(G1888,G1555,G59691);
  nand GNAME1889(G1889,G1731,G58901);
  nand GNAME1890(G1890,G1555,G59692);
  nand GNAME1891(G1891,G1731,G58902);
  nand GNAME1892(G1892,G1555,G59693);
  nand GNAME1893(G1893,G1593,G58880);
  nand GNAME1894(G1894,G20096,G58848);
  nand GNAME1895(G1895,G1593,G58879);
  nand GNAME1896(G1896,G20096,G58847);
  nand GNAME1897(G1897,G1593,G58878);
  nand GNAME1898(G1898,G20096,G58846);
  nand GNAME1899(G1899,G1593,G58877);
  nand GNAME1900(G1900,G20096,G58845);
  nand GNAME1901(G1901,G1593,G58876);
  nand GNAME1902(G1902,G20096,G58844);
  nand GNAME1903(G1903,G1593,G58875);
  nand GNAME1904(G1904,G20096,G58843);
  nand GNAME1905(G1905,G1593,G58874);
  nand GNAME1906(G1906,G20096,G58842);
  nand GNAME1907(G1907,G1593,G58902);
  nand GNAME1908(G1908,G20096,G58870);
  nand GNAME1909(G1909,G1593,G58901);
  nand GNAME1910(G1910,G20096,G58869);
  nand GNAME1911(G1911,G1593,G58873);
  nand GNAME1912(G1912,G20096,G58841);
  nand GNAME1913(G1913,G1593,G58900);
  nand GNAME1914(G1914,G20096,G58868);
  nand GNAME1915(G1915,G1593,G58899);
  nand GNAME1916(G1916,G20096,G58867);
  nand GNAME1917(G1917,G1593,G58898);
  nand GNAME1918(G1918,G20096,G58866);
  nand GNAME1919(G1919,G1593,G58897);
  nand GNAME1920(G1920,G20096,G58865);
  nand GNAME1921(G1921,G1593,G58896);
  nand GNAME1922(G1922,G20096,G58864);
  nand GNAME1923(G1923,G1593,G58895);
  nand GNAME1924(G1924,G20096,G58863);
  nand GNAME1925(G1925,G1593,G58894);
  nand GNAME1926(G1926,G20096,G58862);
  nand GNAME1927(G1927,G1593,G58893);
  nand GNAME1928(G1928,G20096,G58861);
  nand GNAME1929(G1929,G1593,G58892);
  nand GNAME1930(G1930,G20096,G58860);
  nand GNAME1931(G1931,G1593,G58891);
  nand GNAME1932(G1932,G20096,G58859);
  nand GNAME1933(G1933,G1593,G58872);
  nand GNAME1934(G1934,G20096,G58840);
  nand GNAME1935(G1935,G1593,G58890);
  nand GNAME1936(G1936,G20096,G58858);
  nand GNAME1937(G1937,G1593,G58889);
  nand GNAME1938(G1938,G20096,G58857);
  nand GNAME1939(G1939,G1593,G58888);
  nand GNAME1940(G1940,G20096,G58856);
  nand GNAME1941(G1941,G1593,G58887);
  nand GNAME1942(G1942,G20096,G58855);
  nand GNAME1943(G1943,G1593,G58886);
  nand GNAME1944(G1944,G20096,G58854);
  nand GNAME1945(G1945,G1593,G58885);
  nand GNAME1946(G1946,G20096,G58853);
  nand GNAME1947(G1947,G1593,G58884);
  nand GNAME1948(G1948,G20096,G58852);
  nand GNAME1949(G1949,G1593,G58883);
  nand GNAME1950(G1950,G20096,G58851);
  nand GNAME1951(G1951,G1593,G58882);
  nand GNAME1952(G1952,G20096,G58850);
  nand GNAME1953(G1953,G1593,G58881);
  nand GNAME1954(G1954,G20096,G58849);
  nand GNAME1955(G1955,G1593,G58871);
  nand GNAME1956(G1956,G20096,G58839);
  nand GNAME1957(G1957,G1592,G23);
  nand GNAME1958(G1958,G20086,G58848);
  nand GNAME1959(G1959,G1592,G24);
  nand GNAME1960(G1960,G20086,G58847);
  nand GNAME1961(G1961,G1592,G25);
  nand GNAME1962(G1962,G20086,G58846);
  nand GNAME1963(G1963,G1592,G26);
  nand GNAME1964(G1964,G20086,G58845);
  nand GNAME1965(G1965,G1592,G27);
  nand GNAME1966(G1966,G20086,G58844);
  nand GNAME1967(G1967,G1592,G28);
  nand GNAME1968(G1968,G20086,G58843);
  nand GNAME1969(G1969,G1592,G29);
  nand GNAME1970(G1970,G20086,G58842);
  nand GNAME1971(G1971,G1592,G1);
  nand GNAME1972(G1972,G20086,G58870);
  nand GNAME1973(G1973,G1592,G2);
  nand GNAME1974(G1974,G20086,G58869);
  nand GNAME1975(G1975,G1592,G30);
  nand GNAME1976(G1976,G20086,G58841);
  nand GNAME1977(G1977,G1592,G3);
  nand GNAME1978(G1978,G20086,G58868);
  nand GNAME1979(G1979,G1592,G4);
  nand GNAME1980(G1980,G20086,G58867);
  nand GNAME1981(G1981,G1592,G5);
  nand GNAME1982(G1982,G20086,G58866);
  nand GNAME1983(G1983,G1592,G6);
  nand GNAME1984(G1984,G20086,G58865);
  nand GNAME1985(G1985,G1592,G7);
  nand GNAME1986(G1986,G20086,G58864);
  nand GNAME1987(G1987,G1592,G8);
  nand GNAME1988(G1988,G20086,G58863);
  nand GNAME1989(G1989,G1592,G9);
  nand GNAME1990(G1990,G20086,G58862);
  nand GNAME1991(G1991,G1592,G10);
  nand GNAME1992(G1992,G20086,G58861);
  nand GNAME1993(G1993,G1592,G11);
  nand GNAME1994(G1994,G20086,G58860);
  nand GNAME1995(G1995,G1592,G12);
  nand GNAME1996(G1996,G20086,G58859);
  nand GNAME1997(G1997,G1592,G31);
  nand GNAME1998(G1998,G20086,G58840);
  nand GNAME1999(G1999,G1592,G13);
  nand GNAME2000(G2000,G20086,G58858);
  nand GNAME2001(G2001,G1592,G14);
  nand GNAME2002(G2002,G20086,G58857);
  nand GNAME2003(G2003,G1592,G15);
  nand GNAME2004(G2004,G20086,G58856);
  nand GNAME2005(G2005,G1592,G16);
  nand GNAME2006(G2006,G20086,G58855);
  nand GNAME2007(G2007,G1592,G17);
  nand GNAME2008(G2008,G20086,G58854);
  nand GNAME2009(G2009,G1592,G18);
  nand GNAME2010(G2010,G20086,G58853);
  nand GNAME2011(G2011,G1592,G19);
  nand GNAME2012(G2012,G20086,G58852);
  nand GNAME2013(G2013,G1592,G20);
  nand GNAME2014(G2014,G20086,G58851);
  nand GNAME2015(G2015,G1592,G21);
  nand GNAME2016(G2016,G20086,G58850);
  nand GNAME2017(G2017,G1592,G22);
  nand GNAME2018(G2018,G20086,G58849);
  nand GNAME2019(G2019,G1592,G32);
  nand GNAME2020(G2020,G20086,G58839);
  nand GNAME2021(G2021,G1729,G59380);
  nand GNAME2022(G2022,G1728,G58931);
  nand GNAME2023(G2023,G1729,G59381);
  nand GNAME2024(G2024,G1728,G58932);
  nand GNAME2025(G2025,G1729,G59382);
  nand GNAME2026(G2026,G1728,G58933);
  nand GNAME2027(G2027,G1729,G59383);
  nand GNAME2028(G2028,G1728,G58934);
  nand GNAME2029(G2029,G1729,G59384);
  nand GNAME2030(G2030,G1728,G58935);
  nand GNAME2031(G2031,G1729,G59385);
  nand GNAME2032(G2032,G1728,G58936);
  nand GNAME2033(G2033,G1729,G59386);
  nand GNAME2034(G2034,G1728,G58937);
  nand GNAME2035(G2035,G1729,G59387);
  nand GNAME2036(G2036,G1728,G58938);
  nand GNAME2037(G2037,G1729,G59360);
  nand GNAME2038(G2038,G1728,G58911);
  nand GNAME2039(G2039,G1729,G59361);
  nand GNAME2040(G2040,G1728,G58912);
  nand GNAME2041(G2041,G1729,G59362);
  nand GNAME2042(G2042,G1728,G58913);
  nand GNAME2043(G2043,G1729,G59363);
  nand GNAME2044(G2044,G1728,G58914);
  nand GNAME2045(G2045,G1729,G59364);
  nand GNAME2046(G2046,G1728,G58915);
  nand GNAME2047(G2047,G1729,G59365);
  nand GNAME2048(G2048,G1728,G58916);
  nand GNAME2049(G2049,G1729,G59366);
  nand GNAME2050(G2050,G1728,G58917);
  nand GNAME2051(G2051,G1729,G59367);
  nand GNAME2052(G2052,G1728,G58918);
  nand GNAME2053(G2053,G1729,G59368);
  nand GNAME2054(G2054,G1728,G58919);
  nand GNAME2055(G2055,G1729,G59369);
  nand GNAME2056(G2056,G1728,G58920);
  nand GNAME2057(G2057,G1729,G59388);
  nand GNAME2058(G2058,G1728,G58939);
  nand GNAME2059(G2059,G1729,G59370);
  nand GNAME2060(G2060,G1728,G58921);
  nand GNAME2061(G2061,G1729,G59371);
  nand GNAME2062(G2062,G1728,G58922);
  nand GNAME2063(G2063,G1729,G59372);
  nand GNAME2064(G2064,G1728,G58923);
  nand GNAME2065(G2065,G1729,G59373);
  nand GNAME2066(G2066,G1728,G58924);
  nand GNAME2067(G2067,G1729,G59374);
  nand GNAME2068(G2068,G1728,G58925);
  nand GNAME2069(G2069,G1729,G59375);
  nand GNAME2070(G2070,G1728,G58926);
  nand GNAME2071(G2071,G1729,G59376);
  nand GNAME2072(G2072,G1728,G58927);
  nand GNAME2073(G2073,G1729,G59377);
  nand GNAME2074(G2074,G1728,G58928);
  nand GNAME2075(G2075,G1729,G59378);
  nand GNAME2076(G2076,G1728,G58929);
  nand GNAME2077(G2077,G1729,G59379);
  nand GNAME2078(G2078,G1728,G58930);
  nand GNAME2079(G2079,G1729,G59389);
  nand GNAME2080(G2080,G1728,G58940);
  or GNAME2081(G2081,G60017,G2083);
  nand GNAME2082(G2082,G2083,G60017);
  not GNAME2083(G2083,G60016);
  nand GNAME2084(G2084,G2082,G2081);
  not GNAME2085(G2085,G13989);
  not GNAME2086(G2086,G14021);
  nand GNAME2087(G2087,G14026,G15863);
  or GNAME2088(G2088,G15863,G14026);
  nand GNAME2089(G2089,G14014,G8063);
  nand GNAME2090(G2090,G14015,G14289);
  nand GNAME2091(G2091,G14013,G8070);
  or GNAME2092(G2092,G8070,G14013);
  nand GNAME2093(G2093,G8068,G14287);
  or GNAME2094(G2094,G14287,G8068);
  nand GNAME2095(G2095,G14011,G8071);
  or GNAME2096(G2096,G8071,G14011);
  nand GNAME2097(G2097,G8067,G14285);
  or GNAME2098(G2098,G14285,G8067);
  nand GNAME2099(G2099,G14009,G8072);
  or GNAME2100(G2100,G8072,G14009);
  or GNAME2101(G2101,G14307,G8088);
  nand GNAME2102(G2102,G14307,G8088);
  or GNAME2103(G2103,G14008,G14007);
  nand GNAME2104(G2104,G14007,G14008);
  or GNAME2105(G2105,G14006,G8089);
  nand GNAME2106(G2106,G14006,G8089);
  or GNAME2107(G2107,G14282,G14005);
  nand GNAME2108(G2108,G14005,G14282);
  or GNAME2109(G2109,G14004,G8090);
  nand GNAME2110(G2110,G14004,G8090);
  or GNAME2111(G2111,G14281,G14003);
  nand GNAME2112(G2112,G14003,G14281);
  or GNAME2113(G2113,G14002,G8091);
  nand GNAME2114(G2114,G14002,G8091);
  or GNAME2115(G2115,G14280,G14001);
  nand GNAME2116(G2116,G14001,G14280);
  nand GNAME2117(G2117,G14027,G8076);
  nor GNAME2118(G2118,G59346,G7985);
  nor GNAME2119(G2119,G59346,G2771);
  nand GNAME2120(G2120,G3536,G3537,G3538,G3539);
  nand GNAME2121(G2121,G3540,G3541,G3542,G3543);
  nand GNAME2122(G2122,G3544,G3545,G3546,G3547);
  nand GNAME2123(G2123,G3548,G3549,G3550,G3551);
  nand GNAME2124(G2124,G3552,G3553,G3554,G3555);
  nand GNAME2125(G2125,G3556,G3557,G3558,G3559);
  nand GNAME2126(G2126,G3560,G3561,G3562,G3563);
  nand GNAME2127(G2127,G3564,G3565,G3566,G3567);
  nand GNAME2128(G2128,G3568,G3569,G3570,G3571);
  nand GNAME2129(G2129,G3572,G3573,G3574,G3575);
  nand GNAME2130(G2130,G3576,G3577,G3578,G3579);
  nand GNAME2131(G2131,G3580,G3581,G3582,G3583);
  nand GNAME2132(G2132,G3584,G3585,G3586,G3587);
  nand GNAME2133(G2133,G3588,G3589,G3590,G3591);
  nand GNAME2134(G2134,G3592,G3593,G3594,G3595);
  nand GNAME2135(G2135,G3596,G3597,G3598,G3599);
  nand GNAME2136(G2136,G7831,G2817);
  nand GNAME2137(G2137,G7819,G7820);
  or GNAME2138(G2138,G2137,G7805);
  nand GNAME2139(G2139,G7821,G3248,G7820);
  nand GNAME2140(G2140,G3251,G7822,G7823);
  nand GNAME2141(G2141,G3251,G7824,G7825);
  nand GNAME2142(G2142,G3251,G7826,G7827);
  nand GNAME2143(G2143,G3251,G7828,G7829);
  and GNAME2144(G2144,G7015,G7805);
  and GNAME2145(G2145,G7070,G7805);
  and GNAME2146(G2146,G7125,G7805);
  nand GNAME2147(G2147,G7806,G7807);
  nand GNAME2148(G2148,G7808,G7809);
  nand GNAME2149(G2149,G7814,G7812,G7813);
  nand GNAME2150(G2150,G7979,G7980,G2817,G7816);
  nand GNAME2151(G2151,G7981,G7982,G2817,G7817);
  nand GNAME2152(G2152,G7658,G7659,G7660,G7661);
  nand GNAME2153(G2153,G7665,G7666,G7664,G7662,G7663);
  nand GNAME2154(G2154,G7681,G7682,G7680,G7678,G7679);
  nand GNAME2155(G2155,G7686,G7687,G7685,G7683,G7684);
  nand GNAME2156(G2156,G7691,G7692,G7690,G7688,G7689);
  nand GNAME2157(G2157,G7696,G7697,G7695,G7693,G7694);
  nand GNAME2158(G2158,G7701,G7702,G7700,G7698,G7699);
  nand GNAME2159(G2159,G7706,G7707,G7705,G7703,G7704);
  nand GNAME2160(G2160,G7711,G7712,G7710,G7708,G7709);
  nand GNAME2161(G2161,G7716,G7717,G7715,G7713,G7714);
  nand GNAME2162(G2162,G7721,G7722,G7720,G7718,G7719);
  nand GNAME2163(G2163,G7726,G7727,G7725,G7723,G7724);
  nand GNAME2164(G2164,G7740,G7741,G7739,G7737,G7738);
  nand GNAME2165(G2165,G7745,G7746,G7744,G7742,G7743);
  nand GNAME2166(G2166,G7750,G7751,G7749,G7747,G7748);
  nand GNAME2167(G2167,G7755,G7756,G7754,G7752,G7753);
  nand GNAME2168(G2168,G7760,G7761,G7759,G7757,G7758);
  nand GNAME2169(G2169,G7765,G7766,G7764,G7762,G7763);
  nand GNAME2170(G2170,G7770,G7771,G7769,G7767,G7768);
  nand GNAME2171(G2171,G7775,G7776,G7774,G7772,G7773);
  nand GNAME2172(G2172,G7780,G7781,G7779,G7777,G7778);
  nand GNAME2173(G2173,G7785,G7786,G7784,G7782,G7783);
  nand GNAME2174(G2174,G7631,G7632,G7630,G7628,G7629);
  nand GNAME2175(G2175,G7636,G7637,G7635,G7633,G7634);
  nand GNAME2176(G2176,G7641,G7642,G7640,G7638,G7639);
  nand GNAME2177(G2177,G7646,G7647,G7645,G7643,G7644);
  nand GNAME2178(G2178,G7651,G7652,G7650,G7648,G7649);
  nand GNAME2179(G2179,G7656,G7657,G7655,G7653,G7654);
  nand GNAME2180(G2180,G3768,G7669,G7675,G7676,G7671);
  nand GNAME2181(G2181,G3769,G7728,G7734,G7735,G7730);
  nand GNAME2182(G2182,G3770,G7787,G7793,G7794,G7789);
  nand GNAME2183(G2183,G3771,G7796,G7802,G7803,G7798);
  and GNAME2184(G2184,G2128,G2859);
  and GNAME2185(G2185,G2129,G2859);
  and GNAME2186(G2186,G2130,G2859);
  and GNAME2187(G2187,G2131,G2859);
  and GNAME2188(G2188,G2132,G2859);
  and GNAME2189(G2189,G2133,G2859);
  and GNAME2190(G2190,G2134,G2859);
  and GNAME2191(G2191,G2135,G2859);
  nand GNAME2192(G2192,G2875,G3242,G3994,G3799,G3812);
  nand GNAME2193(G2193,G3800,G3994,G7623,G3246);
  nand GNAME2194(G2194,G7498,G7499,G7500,G7501);
  nand GNAME2195(G2195,G7505,G7506,G7504,G7502,G7503);
  nand GNAME2196(G2196,G7520,G7521,G7519,G7517,G7518);
  nand GNAME2197(G2197,G7525,G7526,G7524,G7522,G7523);
  nand GNAME2198(G2198,G7530,G7531,G7529,G7527,G7528);
  nand GNAME2199(G2199,G7535,G7536,G7534,G7532,G7533);
  nand GNAME2200(G2200,G7540,G7541,G7539,G7537,G7538);
  nand GNAME2201(G2201,G7545,G7546,G7544,G7542,G7543);
  nand GNAME2202(G2202,G7550,G7551,G7549,G7547,G7548);
  nand GNAME2203(G2203,G7552,G7553,G7554,G7555);
  nand GNAME2204(G2204,G7556,G7557,G7558,G7559);
  nand GNAME2205(G2205,G7560,G7561,G7562,G7563);
  nand GNAME2206(G2206,G7569,G7570,G7571,G7572);
  nand GNAME2207(G2207,G7573,G7574,G7575,G7576);
  nand GNAME2208(G2208,G7577,G7578,G7579,G7580);
  nand GNAME2209(G2209,G7581,G7582,G7583,G7584);
  nand GNAME2210(G2210,G7585,G7586,G7587,G7588);
  nand GNAME2211(G2211,G7589,G7590,G7591,G7592);
  nand GNAME2212(G2212,G7593,G7594,G7595,G7596);
  nand GNAME2213(G2213,G7597,G7598,G7599,G7600);
  nand GNAME2214(G2214,G7601,G7602,G7603,G7604);
  nand GNAME2215(G2215,G7605,G7606,G7607,G7608);
  nand GNAME2216(G2216,G7471,G7472,G7473,G7474);
  nand GNAME2217(G2217,G7475,G7476,G7477,G7478);
  nand GNAME2218(G2218,G7479,G7480,G7481,G7482);
  nand GNAME2219(G2219,G7483,G7484,G7485,G7486);
  nand GNAME2220(G2220,G7487,G7488,G7489,G7490);
  nand GNAME2221(G2221,G7496,G7497,G7495,G7493,G7494);
  nand GNAME2222(G2222,G7515,G7516,G7514,G7512,G7513);
  nand GNAME2223(G2223,G7567,G7568,G7566,G7564,G7565);
  nand GNAME2224(G2224,G7612,G7613,G7611,G7609,G7610);
  nand GNAME2225(G2225,G7617,G7618,G7616,G7614,G7615);
  and GNAME2226(G2226,G7032,G2867);
  and GNAME2227(G2227,G7087,G2867);
  and GNAME2228(G2228,G7142,G2867);
  and GNAME2229(G2229,G7180,G2867);
  and GNAME2230(G2230,G7236,G2867);
  and GNAME2231(G2231,G7292,G2867);
  and GNAME2232(G2232,G7348,G2867);
  and GNAME2233(G2233,G7404,G2867);
  and GNAME2234(G2234,G59100,G2859);
  and GNAME2235(G2235,G59101,G2859);
  and GNAME2236(G2236,G59102,G2859);
  and GNAME2237(G2237,G59103,G2859);
  and GNAME2238(G2238,G59104,G2859);
  nand GNAME2239(G2239,G7445,G3798,G7444);
  nand GNAME2240(G2240,G3242,G3764,G3956,G3802,G3810);
  nand GNAME2241(G2241,G3800,G7444,G7452,G7453);
  nand GNAME2242(G2242,G7050,G7051,G7052,G7053);
  nand GNAME2243(G2243,G7105,G7106,G7107,G7108);
  nand GNAME2244(G2244,G7160,G7161,G7162,G7163);
  nand GNAME2245(G2245,G7218,G7219,G7217,G7215,G7216);
  nand GNAME2246(G2246,G7274,G7275,G7273,G7271,G7272);
  nand GNAME2247(G2247,G3737,G7328,G3794,G7327);
  nand GNAME2248(G2248,G3750,G3785,G3188,G7383,G7384);
  nand GNAME2249(G2249,G3763,G3794,G3808,G7439,G7440);
  nand GNAME2250(G2250,G6870,G6871,G6872,G6873);
  nand GNAME2251(G2251,G6877,G6878,G6876,G6874,G6875);
  nand GNAME2252(G2252,G6887,G6888,G6886,G6884,G6885);
  nand GNAME2253(G2253,G6892,G6893,G6891,G6889,G6890);
  nand GNAME2254(G2254,G6897,G6898,G6896,G6894,G6895);
  nand GNAME2255(G2255,G6902,G6903,G6901,G6899,G6900);
  nand GNAME2256(G2256,G6907,G6908,G6906,G6904,G6905);
  nand GNAME2257(G2257,G6912,G6913,G6911,G6909,G6910);
  nand GNAME2258(G2258,G6917,G6918,G6916,G6914,G6915);
  nand GNAME2259(G2259,G6922,G6923,G6921,G6919,G6920);
  nand GNAME2260(G2260,G6927,G6928,G6926,G6924,G6925);
  nand GNAME2261(G2261,G6932,G6933,G6931,G6929,G6930);
  nand GNAME2262(G2262,G6942,G6943,G6941,G6939,G6940);
  nand GNAME2263(G2263,G6947,G6948,G6946,G6944,G6945);
  nand GNAME2264(G2264,G6952,G6953,G6951,G6949,G6950);
  nand GNAME2265(G2265,G6957,G6958,G6956,G6954,G6955);
  nand GNAME2266(G2266,G6962,G6963,G6961,G6959,G6960);
  nand GNAME2267(G2267,G6967,G6968,G6966,G6964,G6965);
  nand GNAME2268(G2268,G6972,G6973,G6971,G6969,G6970);
  nand GNAME2269(G2269,G6977,G6978,G6976,G6974,G6975);
  nand GNAME2270(G2270,G6982,G6983,G6981,G6979,G6980);
  nand GNAME2271(G2271,G6987,G6988,G6986,G6984,G6985);
  nand GNAME2272(G2272,G6843,G6844,G6842,G6840,G6841);
  nand GNAME2273(G2273,G6848,G6849,G6847,G6845,G6846);
  nand GNAME2274(G2274,G6853,G6854,G6852,G6850,G6851);
  nand GNAME2275(G2275,G6858,G6859,G6857,G6855,G6856);
  nand GNAME2276(G2276,G6863,G6864,G6862,G6860,G6861);
  nand GNAME2277(G2277,G6868,G6869,G6867,G6865,G6866);
  nand GNAME2278(G2278,G6882,G6883,G6881,G6879,G6880);
  nand GNAME2279(G2279,G6937,G6938,G6936,G6934,G6935);
  nand GNAME2280(G2280,G6992,G6993,G6991,G6989,G6990);
  nand GNAME2281(G2281,G3664,G6996,G6994,G6995);
  and GNAME2282(G2282,G3869,G59149);
  and GNAME2283(G2283,G3869,G59140);
  and GNAME2284(G2284,G3869,G59139);
  and GNAME2285(G2285,G3869,G59138);
  and GNAME2286(G2286,G3869,G59137);
  and GNAME2287(G2287,G3869,G59136);
  and GNAME2288(G2288,G3869,G59135);
  and GNAME2289(G2289,G3869,G59134);
  and GNAME2290(G2290,G3869,G59133);
  and GNAME2291(G2291,G3869,G59132);
  and GNAME2292(G2292,G3869,G59131);
  and GNAME2293(G2293,G3869,G59130);
  and GNAME2294(G2294,G3869,G59129);
  and GNAME2295(G2295,G3869,G59128);
  and GNAME2296(G2296,G3869,G59127);
  and GNAME2297(G2297,G3869,G59126);
  and GNAME2298(G2298,G3869,G59125);
  and GNAME2299(G2299,G3869,G59124);
  and GNAME2300(G2300,G3869,G59123);
  and GNAME2301(G2301,G3869,G59122);
  and GNAME2302(G2302,G3869,G59121);
  and GNAME2303(G2303,G3869,G59120);
  and GNAME2304(G2304,G3869,G59119);
  and GNAME2305(G2305,G3869,G59118);
  and GNAME2306(G2306,G2795,G6582);
  and GNAME2307(G2307,G2795,G6599);
  and GNAME2308(G2308,G2795,G6616);
  and GNAME2309(G2309,G2795,G6633);
  and GNAME2310(G2310,G2795,G6650);
  and GNAME2311(G2311,G2795,G6667);
  and GNAME2312(G2312,G2795,G6684);
  and GNAME2313(G2313,G2795,G6701);
  nand GNAME2314(G2314,G6308,G6306,G6307);
  nand GNAME2315(G2315,G6305,G6303,G6304);
  nand GNAME2316(G2316,G6302,G6300,G6301);
  nand GNAME2317(G2317,G6299,G6297,G6298);
  nand GNAME2318(G2318,G6296,G6294,G6295);
  nand GNAME2319(G2319,G6293,G6291,G6292);
  nand GNAME2320(G2320,G6290,G6288,G6289);
  nand GNAME2321(G2321,G6287,G6285,G6286);
  nand GNAME2322(G2322,G6284,G6282,G6283);
  nand GNAME2323(G2323,G6281,G6279,G6280);
  nand GNAME2324(G2324,G6278,G6276,G6277);
  nand GNAME2325(G2325,G6275,G6273,G6274);
  nand GNAME2326(G2326,G6272,G6270,G6271);
  nand GNAME2327(G2327,G6269,G6267,G6268);
  nand GNAME2328(G2328,G6266,G6264,G6265);
  nand GNAME2329(G2329,G6263,G6261,G6262);
  nand GNAME2330(G2330,G6260,G6258,G6259);
  nand GNAME2331(G2331,G6257,G6255,G6256);
  nand GNAME2332(G2332,G6254,G6252,G6253);
  nand GNAME2333(G2333,G6251,G6249,G6250);
  nand GNAME2334(G2334,G6248,G6246,G6247);
  nand GNAME2335(G2335,G6245,G6243,G6244);
  nand GNAME2336(G2336,G6242,G6240,G6241);
  nand GNAME2337(G2337,G6239,G6237,G6238);
  nand GNAME2338(G2338,G6236,G6234,G6235);
  nand GNAME2339(G2339,G6233,G6231,G6232);
  nand GNAME2340(G2340,G6230,G6228,G6229);
  nand GNAME2341(G2341,G6227,G6225,G6226);
  nand GNAME2342(G2342,G6224,G6222,G6223);
  nand GNAME2343(G2343,G6221,G6219,G6220);
  nand GNAME2344(G2344,G3789,G6218,G7834,G7920,G7921);
  nand GNAME2345(G2345,G3788,G6214,G7832,G7833);
  nand GNAME2346(G2346,G7918,G7919,G6206,G6211);
  and GNAME2347(G2347,G3964,G58946);
  and GNAME2348(G2348,G3964,G58947);
  and GNAME2349(G2349,G3964,G58948);
  and GNAME2350(G2350,G3964,G58949);
  and GNAME2351(G2351,G3964,G58950);
  and GNAME2352(G2352,G3964,G58951);
  and GNAME2353(G2353,G3964,G58952);
  and GNAME2354(G2354,G3964,G58953);
  and GNAME2355(G2355,G3964,G58954);
  and GNAME2356(G2356,G3964,G58955);
  and GNAME2357(G2357,G3964,G58956);
  and GNAME2358(G2358,G3964,G58957);
  and GNAME2359(G2359,G3964,G58958);
  and GNAME2360(G2360,G3964,G58959);
  and GNAME2361(G2361,G3964,G58960);
  and GNAME2362(G2362,G3964,G58961);
  and GNAME2363(G2363,G3964,G58962);
  and GNAME2364(G2364,G3964,G58963);
  and GNAME2365(G2365,G3964,G58964);
  and GNAME2366(G2366,G3964,G58965);
  and GNAME2367(G2367,G3964,G58966);
  and GNAME2368(G2368,G3964,G58967);
  and GNAME2369(G2369,G3964,G58968);
  and GNAME2370(G2370,G3964,G58969);
  and GNAME2371(G2371,G3964,G58970);
  and GNAME2372(G2372,G3964,G58971);
  and GNAME2373(G2373,G3964,G58972);
  and GNAME2374(G2374,G3964,G58973);
  and GNAME2375(G2375,G3964,G58974);
  and GNAME2376(G2376,G3964,G58975);
  nand GNAME2377(G2377,G6205,G2912,G7987);
  nand GNAME2378(G2378,G3801,G3802,G6203,G6204);
  nand GNAME2379(G2379,G6202,G3814,G6201);
  nand GNAME2380(G2380,G7912,G7913,G3813,G3815);
  nand GNAME2381(G2381,G3534,G6182,G6180,G6181);
  nand GNAME2382(G2382,G3533,G6176,G6174,G6175);
  nand GNAME2383(G2383,G3532,G6170,G6168,G6169);
  nand GNAME2384(G2384,G3531,G6164,G6162,G6163);
  nand GNAME2385(G2385,G3530,G6158,G6156,G6157);
  nand GNAME2386(G2386,G3529,G6152,G6150,G6151);
  nand GNAME2387(G2387,G3528,G6146,G6144,G6145);
  nand GNAME2388(G2388,G3527,G6140,G6138,G6139);
  nand GNAME2389(G2389,G3526,G6121,G6119,G6120);
  nand GNAME2390(G2390,G3525,G6115,G6113,G6114);
  nand GNAME2391(G2391,G3524,G6109,G6107,G6108);
  nand GNAME2392(G2392,G3523,G6103,G6101,G6102);
  nand GNAME2393(G2393,G3522,G6097,G6095,G6096);
  nand GNAME2394(G2394,G3521,G6091,G6089,G6090);
  nand GNAME2395(G2395,G3520,G6085,G6083,G6084);
  nand GNAME2396(G2396,G3519,G6079,G6077,G6078);
  nand GNAME2397(G2397,G3518,G6060,G6058,G6059);
  nand GNAME2398(G2398,G3517,G6054,G6052,G6053);
  nand GNAME2399(G2399,G3516,G6048,G6046,G6047);
  nand GNAME2400(G2400,G3515,G6042,G6040,G6041);
  nand GNAME2401(G2401,G3514,G6036,G6034,G6035);
  nand GNAME2402(G2402,G3513,G6030,G6028,G6029);
  nand GNAME2403(G2403,G3512,G6024,G6022,G6023);
  nand GNAME2404(G2404,G3511,G6018,G6016,G6017);
  nand GNAME2405(G2405,G3510,G5999,G5997,G5998);
  nand GNAME2406(G2406,G3509,G5993,G5991,G5992);
  nand GNAME2407(G2407,G3508,G5987,G5985,G5986);
  nand GNAME2408(G2408,G3507,G5981,G5979,G5980);
  nand GNAME2409(G2409,G3506,G5975,G5973,G5974);
  nand GNAME2410(G2410,G3505,G5969,G5967,G5968);
  nand GNAME2411(G2411,G3504,G5963,G5961,G5962);
  nand GNAME2412(G2412,G3503,G5957,G5955,G5956);
  nand GNAME2413(G2413,G3502,G5938,G5936,G5937);
  nand GNAME2414(G2414,G3501,G5932,G5930,G5931);
  nand GNAME2415(G2415,G3500,G5926,G5924,G5925);
  nand GNAME2416(G2416,G3499,G5920,G5918,G5919);
  nand GNAME2417(G2417,G3498,G5914,G5912,G5913);
  nand GNAME2418(G2418,G3497,G5908,G5906,G5907);
  nand GNAME2419(G2419,G3496,G5902,G5900,G5901);
  nand GNAME2420(G2420,G3495,G5896,G5894,G5895);
  nand GNAME2421(G2421,G3494,G5877,G5875,G5876);
  nand GNAME2422(G2422,G3493,G5871,G5869,G5870);
  nand GNAME2423(G2423,G3492,G5865,G5863,G5864);
  nand GNAME2424(G2424,G3491,G5859,G5857,G5858);
  nand GNAME2425(G2425,G3490,G5853,G5851,G5852);
  nand GNAME2426(G2426,G3489,G5847,G5845,G5846);
  nand GNAME2427(G2427,G3488,G5841,G5839,G5840);
  nand GNAME2428(G2428,G3487,G5835,G5833,G5834);
  nand GNAME2429(G2429,G3486,G5816,G5814,G5815);
  nand GNAME2430(G2430,G3485,G5810,G5808,G5809);
  nand GNAME2431(G2431,G3484,G5804,G5802,G5803);
  nand GNAME2432(G2432,G3483,G5798,G5796,G5797);
  nand GNAME2433(G2433,G3482,G5792,G5790,G5791);
  nand GNAME2434(G2434,G3481,G5786,G5784,G5785);
  nand GNAME2435(G2435,G3480,G5780,G5778,G5779);
  nand GNAME2436(G2436,G3479,G5774,G5772,G5773);
  nand GNAME2437(G2437,G3478,G5755,G5753,G5754);
  nand GNAME2438(G2438,G3477,G5749,G5747,G5748);
  nand GNAME2439(G2439,G3476,G5743,G5741,G5742);
  nand GNAME2440(G2440,G3475,G5737,G5735,G5736);
  nand GNAME2441(G2441,G3474,G5731,G5729,G5730);
  nand GNAME2442(G2442,G3473,G5725,G5723,G5724);
  nand GNAME2443(G2443,G3472,G5719,G5717,G5718);
  nand GNAME2444(G2444,G3471,G5713,G5711,G5712);
  nand GNAME2445(G2445,G3470,G5694,G5692,G5693);
  nand GNAME2446(G2446,G3469,G5688,G5686,G5687);
  nand GNAME2447(G2447,G3468,G5682,G5680,G5681);
  nand GNAME2448(G2448,G3467,G5676,G5674,G5675);
  nand GNAME2449(G2449,G3466,G5670,G5668,G5669);
  nand GNAME2450(G2450,G3465,G5664,G5662,G5663);
  nand GNAME2451(G2451,G3464,G5658,G5656,G5657);
  nand GNAME2452(G2452,G3463,G5652,G5650,G5651);
  nand GNAME2453(G2453,G3462,G5633,G5631,G5632);
  nand GNAME2454(G2454,G3461,G5627,G5625,G5626);
  nand GNAME2455(G2455,G3460,G5621,G5619,G5620);
  nand GNAME2456(G2456,G3459,G5615,G5613,G5614);
  nand GNAME2457(G2457,G3458,G5609,G5607,G5608);
  nand GNAME2458(G2458,G3457,G5603,G5601,G5602);
  nand GNAME2459(G2459,G3456,G5597,G5595,G5596);
  nand GNAME2460(G2460,G3455,G5591,G5589,G5590);
  nand GNAME2461(G2461,G3454,G5572,G5570,G5571);
  nand GNAME2462(G2462,G3453,G5566,G5564,G5565);
  nand GNAME2463(G2463,G3452,G5560,G5558,G5559);
  nand GNAME2464(G2464,G3451,G5554,G5552,G5553);
  nand GNAME2465(G2465,G3450,G5548,G5546,G5547);
  nand GNAME2466(G2466,G3449,G5542,G5540,G5541);
  nand GNAME2467(G2467,G3448,G5536,G5534,G5535);
  nand GNAME2468(G2468,G3447,G5530,G5528,G5529);
  nand GNAME2469(G2469,G3446,G5511,G5509,G5510);
  nand GNAME2470(G2470,G3445,G5505,G5503,G5504);
  nand GNAME2471(G2471,G3444,G5499,G5497,G5498);
  nand GNAME2472(G2472,G3443,G5493,G5491,G5492);
  nand GNAME2473(G2473,G3442,G5487,G5485,G5486);
  nand GNAME2474(G2474,G3441,G5481,G5479,G5480);
  nand GNAME2475(G2475,G3440,G5475,G5473,G5474);
  nand GNAME2476(G2476,G3439,G5469,G5467,G5468);
  nand GNAME2477(G2477,G3438,G5450,G5448,G5449);
  nand GNAME2478(G2478,G3437,G5444,G5442,G5443);
  nand GNAME2479(G2479,G3436,G5438,G5436,G5437);
  nand GNAME2480(G2480,G3435,G5432,G5430,G5431);
  nand GNAME2481(G2481,G3434,G5426,G5424,G5425);
  nand GNAME2482(G2482,G3433,G5420,G5418,G5419);
  nand GNAME2483(G2483,G3432,G5414,G5412,G5413);
  nand GNAME2484(G2484,G3431,G5408,G5406,G5407);
  nand GNAME2485(G2485,G3430,G5389,G5387,G5388);
  nand GNAME2486(G2486,G3429,G5383,G5381,G5382);
  nand GNAME2487(G2487,G3428,G5377,G5375,G5376);
  nand GNAME2488(G2488,G3427,G5371,G5369,G5370);
  nand GNAME2489(G2489,G3426,G5365,G5363,G5364);
  nand GNAME2490(G2490,G3425,G5359,G5357,G5358);
  nand GNAME2491(G2491,G3424,G5353,G5351,G5352);
  nand GNAME2492(G2492,G3423,G5347,G5345,G5346);
  nand GNAME2493(G2493,G3422,G5328,G5326,G5327);
  nand GNAME2494(G2494,G3421,G5322,G5320,G5321);
  nand GNAME2495(G2495,G3420,G5316,G5314,G5315);
  nand GNAME2496(G2496,G3419,G5310,G5308,G5309);
  nand GNAME2497(G2497,G3418,G5304,G5302,G5303);
  nand GNAME2498(G2498,G3417,G5298,G5296,G5297);
  nand GNAME2499(G2499,G3416,G5292,G5290,G5291);
  nand GNAME2500(G2500,G3415,G5286,G5284,G5285);
  nand GNAME2501(G2501,G3414,G5267,G5265,G5266);
  nand GNAME2502(G2502,G3413,G5258,G5256,G5257);
  nand GNAME2503(G2503,G3412,G5249,G5247,G5248);
  nand GNAME2504(G2504,G3411,G5240,G5238,G5239);
  nand GNAME2505(G2505,G3410,G5231,G5229,G5230);
  nand GNAME2506(G2506,G3409,G5222,G5220,G5221);
  nand GNAME2507(G2507,G3408,G5213,G5211,G5212);
  nand GNAME2508(G2508,G3407,G5204,G5202,G5203);
  and GNAME2509(G2509,G5043,G59113);
  nand GNAME2510(G2510,G5079,G5077,G5078);
  nand GNAME2511(G2511,G5072,G5070,G5071);
  nand GNAME2512(G2512,G5061,G5059,G5060);
  nand GNAME2513(G2513,G3401,G5035,G5037,G5038);
  nand GNAME2514(G2514,G3400,G5029,G5031,G5032);
  nand GNAME2515(G2515,G3399,G5023,G5025,G5026);
  nand GNAME2516(G2516,G3398,G5017,G5019,G5020);
  nand GNAME2517(G2517,G3397,G5015,G5013,G5014);
  nand GNAME2518(G2518,G3396,G5009,G5007,G5008);
  nand GNAME2519(G2519,G3395,G5003,G5001,G5002);
  nand GNAME2520(G2520,G3394,G4997,G4995,G4996);
  nand GNAME2521(G2521,G3393,G4991,G4989,G4990);
  nand GNAME2522(G2522,G3392,G4985,G4983,G4984);
  nand GNAME2523(G2523,G3391,G4979,G4977,G4978);
  nand GNAME2524(G2524,G3390,G4973,G4971,G4972);
  nand GNAME2525(G2525,G3389,G4967,G4965,G4966);
  nand GNAME2526(G2526,G3388,G4961,G4959,G4960);
  nand GNAME2527(G2527,G3387,G4955,G4953,G4954);
  nand GNAME2528(G2528,G3386,G4949,G4947,G4948);
  nand GNAME2529(G2529,G3385,G4943,G4941,G4942);
  nand GNAME2530(G2530,G3384,G4937,G4935,G4936);
  nand GNAME2531(G2531,G3383,G4931,G4929,G4930);
  nand GNAME2532(G2532,G3382,G4925,G4923,G4924);
  nand GNAME2533(G2533,G3381,G4919,G4917,G4918);
  nand GNAME2534(G2534,G3380,G4913,G4911,G4912);
  nand GNAME2535(G2535,G3379,G4907,G4905,G4906);
  nand GNAME2536(G2536,G3378,G4901,G4899,G4900);
  nand GNAME2537(G2537,G3377,G4895,G4893,G4894);
  nand GNAME2538(G2538,G3376,G4889,G4887,G4888);
  nand GNAME2539(G2539,G3375,G4883,G4881,G4882);
  nand GNAME2540(G2540,G3374,G4877,G4875,G4876);
  nand GNAME2541(G2541,G3373,G4871,G4869,G4870);
  nand GNAME2542(G2542,G3372,G4865,G4863,G4864);
  nand GNAME2543(G2543,G3371,G4859,G4857,G4858);
  nand GNAME2544(G2544,G3370,G4853,G4851,G4852);
  nand GNAME2545(G2545,G4810,G4811,G4809,G4807,G4808);
  nand GNAME2546(G2546,G4805,G4806,G4804,G4802,G4803);
  nand GNAME2547(G2547,G4800,G4801,G4799,G4797,G4798);
  nand GNAME2548(G2548,G4795,G4796,G4794,G4792,G4793);
  nand GNAME2549(G2549,G4790,G4791,G4789,G4787,G4788);
  nand GNAME2550(G2550,G4785,G4786,G4784,G4782,G4783);
  nand GNAME2551(G2551,G4780,G4781,G4779,G4777,G4778);
  nand GNAME2552(G2552,G4775,G4776,G4774,G4772,G4773);
  nand GNAME2553(G2553,G4770,G4771,G4769,G4767,G4768);
  nand GNAME2554(G2554,G4765,G4766,G4764,G4762,G4763);
  nand GNAME2555(G2555,G4760,G4761,G4759,G4757,G4758);
  nand GNAME2556(G2556,G4755,G4756,G4754,G4752,G4753);
  nand GNAME2557(G2557,G4750,G4751,G4749,G4747,G4748);
  nand GNAME2558(G2558,G4745,G4746,G4744,G4742,G4743);
  nand GNAME2559(G2559,G4740,G4741,G4739,G4737,G4738);
  nand GNAME2560(G2560,G4735,G4736,G4734,G4732,G4733);
  nand GNAME2561(G2561,G4730,G4731,G4729,G4727,G4728);
  nand GNAME2562(G2562,G4725,G4726,G4724,G4722,G4723);
  nand GNAME2563(G2563,G4720,G4721,G4719,G4717,G4718);
  nand GNAME2564(G2564,G4715,G4716,G4714,G4712,G4713);
  nand GNAME2565(G2565,G4710,G4711,G4709,G4707,G4708);
  nand GNAME2566(G2566,G4705,G4706,G4704,G4702,G4703);
  nand GNAME2567(G2567,G4700,G4701,G4699,G4697,G4698);
  nand GNAME2568(G2568,G4695,G4696,G4694,G4692,G4693);
  nand GNAME2569(G2569,G4690,G4691,G4689,G4687,G4688);
  nand GNAME2570(G2570,G4685,G4686,G4684,G4682,G4683);
  nand GNAME2571(G2571,G4680,G4681,G4679,G4677,G4678);
  nand GNAME2572(G2572,G4675,G4676,G4674,G4672,G4673);
  nand GNAME2573(G2573,G4670,G4671,G4669,G4667,G4668);
  nand GNAME2574(G2574,G4665,G4666,G4664,G4662,G4663);
  nand GNAME2575(G2575,G4660,G4661,G4659,G4657,G4658);
  nand GNAME2576(G2576,G4655,G4656,G4654,G4652,G4653);
  nand GNAME2577(G2577,G4650,G4648,G4649);
  nand GNAME2578(G2578,G4647,G4645,G4646);
  nand GNAME2579(G2579,G4644,G4642,G4643);
  nand GNAME2580(G2580,G4641,G4639,G4640);
  nand GNAME2581(G2581,G4638,G4636,G4637);
  nand GNAME2582(G2582,G4635,G4633,G4634);
  nand GNAME2583(G2583,G4632,G4630,G4631);
  nand GNAME2584(G2584,G4629,G4627,G4628);
  nand GNAME2585(G2585,G4626,G4624,G4625);
  nand GNAME2586(G2586,G4623,G4621,G4622);
  nand GNAME2587(G2587,G4620,G4618,G4619);
  nand GNAME2588(G2588,G4617,G4615,G4616);
  nand GNAME2589(G2589,G4614,G4612,G4613);
  nand GNAME2590(G2590,G4611,G4609,G4610);
  nand GNAME2591(G2591,G4608,G4606,G4607);
  nand GNAME2592(G2592,G4605,G4603,G4604);
  nand GNAME2593(G2593,G4602,G4601,G4645);
  nand GNAME2594(G2594,G4600,G4599,G4642);
  nand GNAME2595(G2595,G4598,G4597,G4639);
  nand GNAME2596(G2596,G4596,G4595,G4636);
  nand GNAME2597(G2597,G4594,G4593,G4633);
  nand GNAME2598(G2598,G4592,G4591,G4630);
  nand GNAME2599(G2599,G4590,G4589,G4627);
  nand GNAME2600(G2600,G4626,G4587,G4588);
  nand GNAME2601(G2601,G4623,G4585,G4586);
  nand GNAME2602(G2602,G4620,G4583,G4584);
  nand GNAME2603(G2603,G4617,G4581,G4582);
  nand GNAME2604(G2604,G4614,G4579,G4580);
  nand GNAME2605(G2605,G4611,G4577,G4578);
  nand GNAME2606(G2606,G4608,G4575,G4576);
  nand GNAME2607(G2607,G4605,G4573,G4574);
  nand GNAME2608(G2608,G4570,G4568,G4569);
  nand GNAME2609(G2609,G4567,G4565,G4566);
  nand GNAME2610(G2610,G4564,G4562,G4563);
  nand GNAME2611(G2611,G4561,G4559,G4560);
  nand GNAME2612(G2612,G4558,G4556,G4557);
  nand GNAME2613(G2613,G4555,G4553,G4554);
  nand GNAME2614(G2614,G4552,G4550,G4551);
  nand GNAME2615(G2615,G4549,G4547,G4548);
  nand GNAME2616(G2616,G4546,G4544,G4545);
  nand GNAME2617(G2617,G4543,G4541,G4542);
  nand GNAME2618(G2618,G4540,G4538,G4539);
  nand GNAME2619(G2619,G4537,G4535,G4536);
  nand GNAME2620(G2620,G4534,G4532,G4533);
  nand GNAME2621(G2621,G4531,G4529,G4530);
  nand GNAME2622(G2622,G4528,G4526,G4527);
  nand GNAME2623(G2623,G4525,G4523,G4524);
  nand GNAME2624(G2624,G4522,G4520,G4521);
  nand GNAME2625(G2625,G4519,G4517,G4518);
  nand GNAME2626(G2626,G4516,G4514,G4515);
  nand GNAME2627(G2627,G4513,G4511,G4512);
  nand GNAME2628(G2628,G4510,G4508,G4509);
  nand GNAME2629(G2629,G4507,G4505,G4506);
  nand GNAME2630(G2630,G4504,G4502,G4503);
  nand GNAME2631(G2631,G4501,G4499,G4500);
  nand GNAME2632(G2632,G4498,G4496,G4497);
  nand GNAME2633(G2633,G4495,G4493,G4494);
  nand GNAME2634(G2634,G4492,G4490,G4491);
  nand GNAME2635(G2635,G4489,G4487,G4488);
  nand GNAME2636(G2636,G4486,G4484,G4485);
  nand GNAME2637(G2637,G4483,G4481,G4482);
  nand GNAME2638(G2638,G4480,G4478,G4479);
  and GNAME2639(G2639,G2876,G59244);
  nand GNAME2640(G2640,G4469,G4470,G4471,G4472);
  nand GNAME2641(G2641,G4465,G4466,G4467,G4468);
  nand GNAME2642(G2642,G4461,G4462,G4463,G4464);
  nand GNAME2643(G2643,G4457,G4458,G4459,G4460);
  nand GNAME2644(G2644,G4453,G4454,G4455,G4456);
  nand GNAME2645(G2645,G4449,G4450,G4451,G4452);
  nand GNAME2646(G2646,G4445,G4446,G4447,G4448);
  nand GNAME2647(G2647,G4441,G4442,G4443,G4444);
  nand GNAME2648(G2648,G4437,G4438,G4439,G4440);
  nand GNAME2649(G2649,G4433,G4434,G4435,G4436);
  nand GNAME2650(G2650,G4429,G4430,G4431,G4432);
  nand GNAME2651(G2651,G4425,G4426,G4427,G4428);
  nand GNAME2652(G2652,G4421,G4422,G4423,G4424);
  nand GNAME2653(G2653,G4417,G4418,G4419,G4420);
  nand GNAME2654(G2654,G4413,G4414,G4415,G4416);
  nand GNAME2655(G2655,G4409,G4410,G4411,G4412);
  nand GNAME2656(G2656,G4407,G4408,G4406,G4404,G4405);
  nand GNAME2657(G2657,G4402,G4403,G4401,G4399,G4400);
  nand GNAME2658(G2658,G4397,G4398,G4396,G4394,G4395);
  nand GNAME2659(G2659,G4392,G4393,G4391,G4389,G4390);
  nand GNAME2660(G2660,G4387,G4388,G4386,G4384,G4385);
  nand GNAME2661(G2661,G4382,G4383,G4381,G4379,G4380);
  nand GNAME2662(G2662,G4377,G4378,G4376,G4374,G4375);
  nand GNAME2663(G2663,G4372,G4373,G4371,G4369,G4370);
  nand GNAME2664(G2664,G4367,G4368,G4366,G4364,G4365);
  nand GNAME2665(G2665,G4362,G4363,G4361,G4359,G4360);
  nand GNAME2666(G2666,G4357,G4358,G4356,G4354,G4355);
  nand GNAME2667(G2667,G4352,G4353,G4351,G4349,G4350);
  nand GNAME2668(G2668,G4347,G4348,G4346,G4344,G4345);
  nand GNAME2669(G2669,G4342,G4343,G4341,G4339,G4340);
  nand GNAME2670(G2670,G4337,G4338,G4336,G4334,G4335);
  nand GNAME2671(G2671,G4333,G4331,G4332);
  nand GNAME2672(G2672,G4321,G4319,G4320);
  nand GNAME2673(G2673,G4318,G4316,G4317);
  nand GNAME2674(G2674,G4315,G4313,G4314);
  nand GNAME2675(G2675,G4312,G4310,G4311);
  nand GNAME2676(G2676,G4309,G4307,G4308);
  nand GNAME2677(G2677,G4306,G4304,G4305);
  nand GNAME2678(G2678,G4303,G4301,G4302);
  nand GNAME2679(G2679,G4300,G4298,G4299);
  nand GNAME2680(G2680,G4297,G4295,G4296);
  nand GNAME2681(G2681,G4294,G4292,G4293);
  nand GNAME2682(G2682,G4291,G4289,G4290);
  nand GNAME2683(G2683,G4288,G4286,G4287);
  nand GNAME2684(G2684,G4285,G4283,G4284);
  nand GNAME2685(G2685,G4282,G4280,G4281);
  nand GNAME2686(G2686,G4279,G4277,G4278);
  nand GNAME2687(G2687,G4276,G4274,G4275);
  nand GNAME2688(G2688,G4273,G4271,G4272);
  nand GNAME2689(G2689,G4270,G4268,G4269);
  nand GNAME2690(G2690,G4267,G4265,G4266);
  nand GNAME2691(G2691,G4264,G4262,G4263);
  nand GNAME2692(G2692,G4261,G4259,G4260);
  nand GNAME2693(G2693,G4258,G4256,G4257);
  nand GNAME2694(G2694,G4255,G4253,G4254);
  nand GNAME2695(G2695,G4252,G4250,G4251);
  nand GNAME2696(G2696,G4249,G4247,G4248);
  nand GNAME2697(G2697,G4246,G4244,G4245);
  nand GNAME2698(G2698,G4243,G4241,G4242);
  nand GNAME2699(G2699,G4240,G4238,G4239);
  nand GNAME2700(G2700,G4237,G4235,G4236);
  nand GNAME2701(G2701,G4234,G4232,G4233);
  nand GNAME2702(G2702,G4231,G4229,G4230);
  nand GNAME2703(G2703,G4227,G4228);
  nand GNAME2704(G2704,G3365,G4218,G4220,G4221);
  nand GNAME2705(G2705,G3364,G4212,G4214,G4215);
  nand GNAME2706(G2706,G4210,G3363,G4207,G4205,G4206);
  nand GNAME2707(G2707,G4204,G3362,G4201,G4199,G4200);
  nand GNAME2708(G2708,G3361,G4194,G4196,G4197);
  nand GNAME2709(G2709,G3360,G4188,G4190,G4191);
  nand GNAME2710(G2710,G3359,G4180,G4177,G4178,G4179);
  nand GNAME2711(G2711,G3358,G4174,G4171,G4172,G4173);
  nand GNAME2712(G2712,G3357,G4168,G4165,G4166,G4167);
  nand GNAME2713(G2713,G3356,G4162,G4159,G4160,G4163);
  nand GNAME2714(G2714,G3355,G4157,G4153,G4154,G4155);
  nand GNAME2715(G2715,G3354,G4151,G4147,G4148,G4149);
  nand GNAME2716(G2716,G3353,G4145,G4141,G4142,G4143);
  nand GNAME2717(G2717,G3352,G4139,G4135,G4136,G4137);
  nand GNAME2718(G2718,G3351,G4133,G4129,G4130,G4131);
  nand GNAME2719(G2719,G3350,G4127,G4123,G4124,G4125);
  nand GNAME2720(G2720,G3349,G4121,G4117,G4118,G4119);
  nand GNAME2721(G2721,G3348,G4115,G4111,G4112,G4113);
  nand GNAME2722(G2722,G3347,G4109,G4105,G4106,G4107);
  nand GNAME2723(G2723,G3346,G4103,G4099,G4100,G4101);
  nand GNAME2724(G2724,G3345,G4096,G4092,G4093);
  nand GNAME2725(G2725,G3344,G4090,G4086,G4087);
  nand GNAME2726(G2726,G3343,G4084,G4080,G4081);
  nand GNAME2727(G2727,G3342,G4078,G4074,G4075);
  nand GNAME2728(G2728,G3341,G4072,G4068,G4069);
  nand GNAME2729(G2729,G3340,G4066,G4062,G4063);
  nand GNAME2730(G2730,G3339,G4060,G4056,G4057);
  nand GNAME2731(G2731,G3338,G4054,G4050,G4051);
  nand GNAME2732(G2732,G3337,G4048,G4044,G4045);
  nand GNAME2733(G2733,G3336,G4042,G4038,G4039);
  nand GNAME2734(G2734,G3335,G4036,G4032,G4033);
  nand GNAME2735(G2735,G3334,G4030,G4026,G4027);
  nand GNAME2736(G2736,G4014,G3811,G2834);
  nand GNAME2737(G2737,G4013,G4011,G4012);
  nand GNAME2738(G2738,G4009,G3811,G2835);
  nand GNAME2739(G2739,G2835,G7853,G7854);
  nand GNAME2740(G2740,G4007,G4006);
  nand GNAME2741(G2741,G4004,G4005);
  nand GNAME2742(G2742,G3817,G7846,G7847);
  nand GNAME2743(G2743,G3817,G7842,G7843);
  nand GNAME2744(G2744,G3973,G3974);
  nand GNAME2745(G2745,G3965,G3964);
  and GNAME2746(G2746,G2783,G3852);
  nand GNAME2747(G2747,G7863,G7864,G5050,G5051);
  and GNAME2748(G2748,G2799,G3835);
  nand GNAME2749(G2749,G3302,G3303,G3304,G3305);
  and GNAME2750(G2750,G6187,G3107);
  not GNAME2751(G2751,G33);
  not GNAME2752(G2752,G1590);
  nand GNAME2753(G2753,G2894,G3835,G3852);
  not GNAME2754(G2754,G58977);
  not GNAME2755(G2755,G59112);
  and GNAME2756(G2756,G2771,G2764);
  and GNAME2757(G2757,G2759,G59112);
  and GNAME2758(G2758,G2756,G2757);
  not GNAME2759(G2759,G59111);
  and GNAME2760(G2760,G2755,G59111);
  and GNAME2761(G2761,G2756,G2760);
  and GNAME2762(G2762,G59112,G59111);
  and GNAME2763(G2763,G2756,G2762);
  not GNAME2764(G2764,G59110);
  nor GNAME2765(G2765,G59109,G2764);
  nor GNAME2766(G2766,G59112,G59111);
  and GNAME2767(G2767,G2765,G2766);
  and GNAME2768(G2768,G2757,G2765);
  and GNAME2769(G2769,G2760,G2765);
  and GNAME2770(G2770,G2762,G2765);
  not GNAME2771(G2771,G59109);
  and GNAME2772(G2772,G2764,G59109);
  and GNAME2773(G2773,G2766,G2772);
  and GNAME2774(G2774,G2757,G2772);
  and GNAME2775(G2775,G2760,G2772);
  nor GNAME2776(G2776,G3790,G3791);
  nor GNAME2777(G2777,G2764,G2771);
  and GNAME2778(G2778,G2766,G2777);
  and GNAME2779(G2779,G2757,G2777);
  and GNAME2780(G2780,G2760,G2777);
  and GNAME2781(G2781,G2762,G2777);
  and GNAME2782(G2782,G2756,G2766);
  nand GNAME2783(G2783,G3318,G3319,G3320,G3321);
  nand GNAME2784(G2784,G3322,G3323,G3324,G3325);
  nand GNAME2785(G2785,G3306,G3307,G3308,G3309);
  nand GNAME2786(G2786,G3310,G3311,G3312,G3313);
  and GNAME2787(G2787,G3920,G3903);
  and GNAME2788(G2788,G3886,G2748,G2795);
  and GNAME2789(G2789,G2855,G2749,G2787,G2788);
  not GNAME2790(G2790,G58979);
  and GNAME2791(G2791,G2789,G58979);
  not GNAME2792(G2792,G20773);
  and GNAME2793(G2793,G2817,G58977);
  nor GNAME2794(G2794,G3835,G2786);
  nand GNAME2795(G2795,G3294,G3295,G3296,G3297);
  and GNAME2796(G2796,G2794,G2785,G2855);
  nand GNAME2797(G2797,G2784,G3954,G3869,G2796);
  nor GNAME2798(G2798,G58978,G2790);
  nand GNAME2799(G2799,G3314,G3315,G3316,G3317);
  nor GNAME2800(G2800,G2785,G2799);
  nor GNAME2801(G2801,G2784,G3937,G3954);
  nand GNAME2802(G2802,G2800,G2801,G3903,G2795,G3835);
  and GNAME2803(G2803,G58979,G2793);
  not GNAME2804(G2804,G20108);
  and GNAME2805(G2805,G2817,G2754);
  nand GNAME2806(G2806,G2881,G3960);
  not GNAME2807(G2807,G58942);
  nand GNAME2808(G2808,G2820,G58942);
  not GNAME2809(G2809,G58943);
  or GNAME2810(G2810,G3963,G2815);
  and GNAME2811(G2811,G3967,G3808,G2855);
  and GNAME2812(G2812,G3806,G3970,G3971,G2811);
  and GNAME2813(G2813,G2837,G2805);
  and GNAME2814(G2814,G2809,G58942);
  and GNAME2815(G2815,G2807,G2809);
  and GNAME2816(G2816,G2790,G58977);
  not GNAME2817(G2817,G58978);
  nand GNAME2818(G2818,G2816,G58978);
  nor GNAME2819(G2819,G2910,G58976);
  not GNAME2820(G2820,G58941);
  nand GNAME2821(G2821,G3979,G2809);
  not GNAME2822(G2822,G59348);
  and GNAME2823(G2823,G58977,G3852);
  and GNAME2824(G2824,G3886,G2796);
  and GNAME2825(G2825,G2824,G2795,G2749);
  and GNAME2826(G2826,G2855,G3920);
  and GNAME2827(G2827,G2749,G3869);
  and GNAME2828(G2828,G2826,G2827,G3886,G2746,G2786);
  and GNAME2829(G2829,G2795,G2786);
  and GNAME2830(G2830,G2799,G3920);
  and GNAME2831(G2831,G2783,G2801,G2829,G2830);
  and GNAME2832(G2832,G3327,G3329,G3331,G3333);
  not GNAME2833(G2833,G59309);
  or GNAME2834(G2834,G7988,G59310,G58945);
  nand GNAME2835(G2835,G2832,G59310);
  and GNAME2836(G2836,G2822,G58978);
  not GNAME2837(G2837,G58976);
  and GNAME2838(G2838,G2752,G2822);
  nor GNAME2839(G2839,G4015,G2754);
  and GNAME2840(G2840,G4025,G2839);
  not GNAME2841(G2841,G3285);
  nor GNAME2842(G2842,G58977,G2790);
  and GNAME2843(G2843,G2845,G2842);
  and GNAME2844(G2844,G2800,G3980,G2838,G2839);
  nand GNAME2845(G2845,G3814,G3815,G4831,G7983);
  nand GNAME2846(G2846,G4017,G4018);
  not GNAME2847(G2847,G20180);
  not GNAME2848(G2848,G20507);
  not GNAME2849(G2849,G20141);
  not GNAME2850(G2850,G20446);
  not GNAME2851(G2851,G20233);
  not GNAME2852(G2852,G20552);
  not GNAME2853(G2853,G20209);
  not GNAME2854(G2854,G20505);
  nand GNAME2855(G2855,G3298,G3299,G3300,G3301);
  and GNAME2856(G2856,G3954,G3886);
  nor GNAME2857(G2857,G3808,G2786,G2855);
  nand GNAME2858(G2858,G2748,G2795,G2785,G2857);
  and GNAME2859(G2859,G58979,G2831);
  nand GNAME2860(G2860,G4226,G2793);
  nor GNAME2861(G2861,G2749,G2860);
  nor GNAME2862(G2862,G3954,G2860);
  and GNAME2863(G2863,G2785,G3835);
  nand GNAME2864(G2864,G3869,G3852,G2857,G2863);
  and GNAME2865(G2865,G7989,G3852);
  nand GNAME2866(G2866,G58979,G2865);
  and GNAME2867(G2867,G58979,G2828);
  nand GNAME2868(G2868,G4330,G2793);
  nor GNAME2869(G2869,G3808,G2868);
  nor GNAME2870(G2870,G3886,G2868);
  nor GNAME2871(G2871,G3869,G2868);
  nor GNAME2872(G2872,G3792,G2868);
  nor GNAME2873(G2873,G2890,G2868);
  and GNAME2874(G2874,G2799,G7989);
  nand GNAME2875(G2875,G3958,G3979,G58979);
  and GNAME2876(G2876,G2818,G4477);
  nor GNAME2877(G2877,G2876,G58979);
  nor GNAME2878(G2878,G2876,G2790);
  and GNAME2879(G2879,G2795,G2878);
  nand GNAME2880(G2880,G3958,G2803);
  nand GNAME2881(G2881,G2793,G2791,G20773);
  and GNAME2882(G2882,G4571,G4572);
  nor GNAME2883(G2883,G2882,G2799);
  nor GNAME2884(G2884,G2882,G3852);
  and GNAME2885(G2885,G4006,G4651);
  nor GNAME2886(G2886,G3246,G2885);
  nor GNAME2887(G2887,G2885,G3799);
  nor GNAME2888(G2888,G2885,G2790);
  nor GNAME2889(G2889,G2885,G3800);
  and GNAME2890(G2890,G3886,G3869);
  and GNAME2891(G2891,G3366,G2811,G4816,G4817);
  nor GNAME2892(G2892,G2909,G2754);
  and GNAME2893(G2893,G2828,G2892);
  nor GNAME2894(G2894,G3808,G3937,G2795);
  and GNAME2895(G2895,G4812,G7855,G7856);
  and GNAME2896(G2896,G4813,G4837);
  and GNAME2897(G2897,G2799,G3869);
  and GNAME2898(G2898,G3368,G2896,G4842,G2895);
  and GNAME2899(G2899,G3367,G3937,G3903,G2800);
  and GNAME2900(G2900,G2794,G2897,G3954,G2784,G2785);
  and GNAME2901(G2901,G4845,G4846);
  and GNAME2902(G2902,G2858,G2901);
  and GNAME2903(G2903,G3369,G2802,G2898);
  and GNAME2904(G2904,G4847,G2892);
  and GNAME2905(G2905,G5103,G4473);
  and GNAME2906(G2906,G4835,G2892);
  and GNAME2907(G2907,G4832,G2892);
  nor GNAME2908(G2908,G58977,G2909);
  and GNAME2909(G2909,G4830,G4831);
  and GNAME2910(G2910,G58977,G58978);
  and GNAME2911(G2911,G58979,G2910);
  nand GNAME2912(G2912,G2790,G58976);
  nand GNAME2913(G2913,G5040,G7861,G7862);
  not GNAME2914(G2914,G59117);
  nor GNAME2915(G2915,G2935,G5045,G2754,G2790);
  and GNAME2916(G2916,G7868,G7869,G3797,G5044);
  nand GNAME2917(G2917,G5046,G2922);
  nor GNAME2918(G2918,G3799,G58977,G5043);
  and GNAME2919(G2919,G2920,G5049);
  nand GNAME2920(G2920,G5041,G3816,G5042);
  not GNAME2921(G2921,G59116);
  or GNAME2922(G2922,G2916,G2915);
  nand GNAME2923(G2923,G5052,G5053);
  nand GNAME2924(G2924,G5057,G5055,G5056);
  not GNAME2925(G2925,G59115);
  and GNAME2926(G2926,G59117,G59116);
  and GNAME2927(G2927,G5064,G5062,G5063);
  nand GNAME2928(G2928,G5066,G5067);
  nand GNAME2929(G2929,G5068,G3775);
  nor GNAME2930(G2930,G59114,G2925);
  not GNAME2931(G2931,G59114);
  nor GNAME2932(G2932,G58977,G2804);
  nand GNAME2933(G2933,G5092,G59112);
  nand GNAME2934(G2934,G5098,G2936);
  and GNAME2935(G2935,G7867,G58978);
  nand GNAME2936(G2936,G5095,G5096);
  nand GNAME2937(G2937,G5120,G5121);
  nand GNAME2938(G2938,G5142,G5143);
  nand GNAME2939(G2939,G5139,G5140);
  nand GNAME2940(G2940,G5145,G3780);
  nand GNAME2941(G2941,G5174,G7904,G7905);
  nand GNAME2942(G2942,G5169,G5171);
  and GNAME2943(G2943,G58978,G59348);
  nand GNAME2944(G2944,G5167,G5162);
  nor GNAME2945(G2945,G7889,G2944);
  nor GNAME2946(G2946,G5099,G7895);
  nor GNAME2947(G2947,G5041,G3798);
  nor GNAME2948(G2948,G7882,G3253);
  nor GNAME2949(G2949,G5069,G5047);
  nand GNAME2950(G2950,G2948,G2949);
  nor GNAME2951(G2951,G2963,G7986);
  and GNAME2952(G2952,G5189,G2951);
  nor GNAME2953(G2953,G59115,G59114);
  nor GNAME2954(G2954,G59116,G59117);
  or GNAME2955(G2955,G2985,G2996);
  or GNAME2956(G2956,G5073,G3041,G3048);
  nor GNAME2957(G2957,G3254,G2956);
  nor GNAME2958(G2958,G2914,G2955);
  and GNAME2959(G2959,G2957,G2958);
  and GNAME2960(G2960,G2953,G2954);
  nor GNAME2961(G2961,G2959,G5194);
  and GNAME2962(G2962,G2913,G58871);
  and GNAME2963(G2963,G2945,G2946);
  and GNAME2964(G2964,G58895,G2947);
  nor GNAME2965(G2965,G5041,G3800);
  and GNAME2966(G2966,G2913,G58872);
  and GNAME2967(G2967,G58896,G2947);
  and GNAME2968(G2968,G2913,G58873);
  and GNAME2969(G2969,G58897,G2947);
  and GNAME2970(G2970,G2913,G58874);
  and GNAME2971(G2971,G58898,G2947);
  and GNAME2972(G2972,G2913,G58875);
  and GNAME2973(G2973,G58899,G2947);
  and GNAME2974(G2974,G2913,G58876);
  and GNAME2975(G2975,G58900,G2947);
  and GNAME2976(G2976,G2913,G58877);
  and GNAME2977(G2977,G58901,G2947);
  and GNAME2978(G2978,G2913,G58878);
  and GNAME2979(G2979,G58902,G2947);
  nor GNAME2980(G2980,G7895,G2934);
  nor GNAME2981(G2981,G5069,G2917);
  nand GNAME2982(G2982,G2948,G2981);
  nor GNAME2983(G2983,G2990,G7986);
  and GNAME2984(G2984,G5271,G2983);
  and GNAME2985(G2985,G2921,G59117);
  nor GNAME2986(G2986,G59117,G2955);
  and GNAME2987(G2987,G2957,G2986);
  and GNAME2988(G2988,G2953,G2985);
  nor GNAME2989(G2989,G2987,G5276);
  and GNAME2990(G2990,G2945,G2980);
  nor GNAME2991(G2991,G3256,G2944);
  nor GNAME2992(G2992,G7876,G7882);
  nand GNAME2993(G2993,G2949,G2992);
  nor GNAME2994(G2994,G3001,G7986);
  and GNAME2995(G2995,G5332,G2994);
  and GNAME2996(G2996,G2914,G59116);
  and GNAME2997(G2997,G2955,G59117);
  and GNAME2998(G2998,G2957,G2997);
  and GNAME2999(G2999,G2953,G2996);
  nor GNAME3000(G3000,G2998,G5337);
  and GNAME3001(G3001,G2946,G2991);
  nand GNAME3002(G3002,G2981,G2992);
  nor GNAME3003(G3003,G3009,G7986);
  and GNAME3004(G3004,G5393,G3003);
  and GNAME3005(G3005,G2955,G2914);
  and GNAME3006(G3006,G2957,G3005);
  and GNAME3007(G3007,G2926,G2953);
  nor GNAME3008(G3008,G3006,G5398);
  and GNAME3009(G3009,G2980,G2991);
  nor GNAME3010(G3010,G5099,G3267);
  nor GNAME3011(G3011,G5047,G2929);
  nand GNAME3012(G3012,G2948,G3011);
  nor GNAME3013(G3013,G3019,G7986);
  and GNAME3014(G3014,G5454,G3013);
  nor GNAME3015(G3015,G7879,G2956);
  and GNAME3016(G3016,G2958,G3015);
  and GNAME3017(G3017,G2930,G2954);
  nor GNAME3018(G3018,G3016,G5459);
  and GNAME3019(G3019,G2945,G3010);
  nor GNAME3020(G3020,G2934,G3267);
  nor GNAME3021(G3021,G2917,G2929);
  nand GNAME3022(G3022,G2948,G3021);
  nor GNAME3023(G3023,G3028,G7986);
  and GNAME3024(G3024,G5515,G3023);
  and GNAME3025(G3025,G2986,G3015);
  and GNAME3026(G3026,G2930,G2985);
  nor GNAME3027(G3027,G3025,G5520);
  and GNAME3028(G3028,G2945,G3020);
  nand GNAME3029(G3029,G2992,G3011);
  nor GNAME3030(G3030,G3035,G7986);
  and GNAME3031(G3031,G5576,G3030);
  and GNAME3032(G3032,G2997,G3015);
  and GNAME3033(G3033,G2930,G2996);
  nor GNAME3034(G3034,G3032,G5581);
  and GNAME3035(G3035,G2991,G3010);
  nand GNAME3036(G3036,G2992,G3021);
  nor GNAME3037(G3037,G3042,G7986);
  and GNAME3038(G3038,G5637,G3037);
  and GNAME3039(G3039,G3005,G3015);
  nor GNAME3040(G3040,G3039,G5642);
  and GNAME3041(G3041,G2926,G2930);
  and GNAME3042(G3042,G2991,G3020);
  nor GNAME3043(G3043,G5168,G7889);
  nor GNAME3044(G3044,G3255,G3253);
  nand GNAME3045(G3045,G2949,G3044);
  nor GNAME3046(G3046,G3053,G7986);
  and GNAME3047(G3047,G5698,G3046);
  and GNAME3048(G3048,G2925,G59114);
  and GNAME3049(G3049,G2956,G7879);
  and GNAME3050(G3050,G2958,G3049);
  and GNAME3051(G3051,G2954,G3048);
  nor GNAME3052(G3052,G3050,G5703);
  and GNAME3053(G3053,G2946,G3043);
  nand GNAME3054(G3054,G2981,G3044);
  nor GNAME3055(G3055,G3060,G7986);
  and GNAME3056(G3056,G5759,G3055);
  and GNAME3057(G3057,G2986,G3049);
  and GNAME3058(G3058,G2985,G3048);
  nor GNAME3059(G3059,G3057,G5764);
  and GNAME3060(G3060,G2980,G3043);
  nor GNAME3061(G3061,G5168,G3256);
  nor GNAME3062(G3062,G7876,G3255);
  nand GNAME3063(G3063,G2949,G3062);
  nor GNAME3064(G3064,G3069,G7986);
  and GNAME3065(G3065,G5820,G3064);
  and GNAME3066(G3066,G2997,G3049);
  and GNAME3067(G3067,G2996,G3048);
  nor GNAME3068(G3068,G3066,G5825);
  and GNAME3069(G3069,G2946,G3061);
  nand GNAME3070(G3070,G2981,G3062);
  nor GNAME3071(G3071,G3076,G7986);
  and GNAME3072(G3072,G5881,G3071);
  and GNAME3073(G3073,G3005,G3049);
  and GNAME3074(G3074,G2926,G3048);
  nor GNAME3075(G3075,G3073,G5886);
  and GNAME3076(G3076,G2980,G3061);
  nand GNAME3077(G3077,G3011,G3044);
  nor GNAME3078(G3078,G3085,G7986);
  and GNAME3079(G3079,G5942,G3078);
  nor GNAME3080(G3080,G2925,G2931);
  and GNAME3081(G3081,G2956,G3254);
  and GNAME3082(G3082,G2958,G3081);
  and GNAME3083(G3083,G2954,G3080);
  nor GNAME3084(G3084,G3082,G5947);
  and GNAME3085(G3085,G3010,G3043);
  nand GNAME3086(G3086,G3021,G3044);
  nor GNAME3087(G3087,G3092,G7986);
  and GNAME3088(G3088,G6003,G3087);
  and GNAME3089(G3089,G2986,G3081);
  and GNAME3090(G3090,G2985,G3080);
  nor GNAME3091(G3091,G3089,G6008);
  and GNAME3092(G3092,G3020,G3043);
  nand GNAME3093(G3093,G3011,G3062);
  nor GNAME3094(G3094,G3099,G7986);
  and GNAME3095(G3095,G6064,G3094);
  and GNAME3096(G3096,G2997,G3081);
  and GNAME3097(G3097,G2996,G3080);
  nor GNAME3098(G3098,G3096,G6069);
  and GNAME3099(G3099,G3010,G3061);
  nand GNAME3100(G3100,G3021,G3062);
  nor GNAME3101(G3101,G3106,G7986);
  and GNAME3102(G3102,G6125,G3101);
  and GNAME3103(G3103,G3005,G3081);
  nor GNAME3104(G3104,G3103,G6130);
  and GNAME3105(G3105,G2926,G3080);
  and GNAME3106(G3106,G3020,G3061);
  and GNAME3107(G3107,G3992,G2812);
  and GNAME3108(G3108,G3796,G3795);
  nor GNAME3109(G3109,G3535,G2750,G20784,G2825);
  nand GNAME3110(G3110,G7910,G7911,G6192,G58977);
  nor GNAME3111(G3111,G58978,G58976);
  not GNAME3112(G3112,G34);
  nand GNAME3113(G3113,G6208,G58941);
  and GNAME3114(G3114,G2820,G2814);
  and GNAME3115(G3115,G2814,G58941);
  nor GNAME3116(G3116,G20552,G20446);
  nor GNAME3117(G3117,G20507,G2854);
  and GNAME3118(G3118,G3116,G3117);
  nor GNAME3119(G3119,G20446,G2852);
  nor GNAME3120(G3120,G20505,G20507);
  and GNAME3121(G3121,G3119,G3120);
  and GNAME3122(G3122,G3117,G3119);
  nor GNAME3123(G3123,G20552,G2850);
  and GNAME3124(G3124,G3120,G3123);
  and GNAME3125(G3125,G3117,G3123);
  nor GNAME3126(G3126,G2850,G2852);
  and GNAME3127(G3127,G3120,G3126);
  and GNAME3128(G3128,G3117,G3126);
  nor GNAME3129(G3129,G20505,G2848);
  and GNAME3130(G3130,G3116,G3129);
  nor GNAME3131(G3131,G2848,G2854);
  and GNAME3132(G3132,G3116,G3131);
  and GNAME3133(G3133,G3119,G3129);
  and GNAME3134(G3134,G3119,G3131);
  and GNAME3135(G3135,G3123,G3129);
  and GNAME3136(G3136,G3123,G3131);
  and GNAME3137(G3137,G3126,G3129);
  and GNAME3138(G3138,G3126,G3131);
  and GNAME3139(G3139,G3116,G3120);
  nand GNAME3140(G3140,G3791,G7933,G7934);
  nor GNAME3141(G3141,G3259,G3140);
  and GNAME3142(G3142,G2762,G3141);
  and GNAME3143(G3143,G2766,G3141);
  and GNAME3144(G3144,G2757,G3141);
  nor GNAME3145(G3145,G7932,G3140);
  and GNAME3146(G3146,G2760,G3145);
  and GNAME3147(G3147,G2762,G3145);
  and GNAME3148(G3148,G2766,G3145);
  and GNAME3149(G3149,G2757,G3145);
  nor GNAME3150(G3150,G6437,G3259);
  and GNAME3151(G3151,G2760,G3150);
  and GNAME3152(G3152,G2762,G3150);
  and GNAME3153(G3153,G2766,G3150);
  and GNAME3154(G3154,G2757,G3150);
  nor GNAME3155(G3155,G6437,G7932);
  and GNAME3156(G3156,G2760,G3155);
  and GNAME3157(G3157,G2762,G3155);
  and GNAME3158(G3158,G2766,G3155);
  and GNAME3159(G3159,G2757,G3155);
  and GNAME3160(G3160,G2760,G3141);
  nor GNAME3161(G3161,G3809,G7901);
  nor GNAME3162(G3162,G5125,G2755);
  and GNAME3163(G3163,G3161,G3162);
  nand GNAME3164(G3164,G5124,G59111);
  nor GNAME3165(G3165,G59112,G3164);
  and GNAME3166(G3166,G3161,G3165);
  nor GNAME3167(G3167,G2755,G3164);
  and GNAME3168(G3168,G3161,G3167);
  nor GNAME3169(G3169,G3809,G3257);
  nor GNAME3170(G3170,G59112,G5125);
  and GNAME3171(G3171,G3169,G3170);
  and GNAME3172(G3172,G3162,G3169);
  and GNAME3173(G3173,G3165,G3169);
  and GNAME3174(G3174,G3167,G3169);
  nor GNAME3175(G3175,G7901,G2942);
  and GNAME3176(G3176,G3170,G3175);
  and GNAME3177(G3177,G3162,G3175);
  and GNAME3178(G3178,G3165,G3175);
  and GNAME3179(G3179,G3167,G3175);
  nor GNAME3180(G3180,G3257,G2942);
  and GNAME3181(G3181,G3170,G3180);
  and GNAME3182(G3182,G3162,G3180);
  and GNAME3183(G3183,G3165,G3180);
  and GNAME3184(G3184,G3167,G3180);
  and GNAME3185(G3185,G3161,G3170);
  nor GNAME3186(G3186,G20108,G3852);
  and GNAME3187(G3187,G2794,G3186);
  nand GNAME3188(G3188,G3835,G2795,G3979);
  nor GNAME3189(G3189,G2799,G3188);
  or GNAME3190(G3190,G2757,G2760);
  nor GNAME3191(G3191,G5175,G3190);
  nor GNAME3192(G3192,G59112,G5146);
  and GNAME3193(G3193,G3191,G3192);
  nor GNAME3194(G3194,G5123,G5175);
  nor GNAME3195(G3195,G5146,G2755);
  and GNAME3196(G3196,G3194,G3195);
  and GNAME3197(G3197,G3192,G3194);
  nor GNAME3198(G3198,G2755,G2940);
  and GNAME3199(G3199,G3191,G3198);
  nor GNAME3200(G3200,G59112,G2940);
  and GNAME3201(G3201,G3191,G3200);
  and GNAME3202(G3202,G3194,G3198);
  and GNAME3203(G3203,G3194,G3200);
  nor GNAME3204(G3204,G2941,G3190);
  and GNAME3205(G3205,G3195,G3204);
  and GNAME3206(G3206,G3192,G3204);
  nor GNAME3207(G3207,G5123,G2941);
  and GNAME3208(G3208,G3195,G3207);
  and GNAME3209(G3209,G3192,G3207);
  and GNAME3210(G3210,G3198,G3204);
  and GNAME3211(G3211,G3200,G3204);
  and GNAME3212(G3212,G3198,G3207);
  and GNAME3213(G3213,G3200,G3207);
  and GNAME3214(G3214,G3191,G3195);
  nor GNAME3215(G3215,G20141,G20180);
  nor GNAME3216(G3216,G20233,G2853);
  and GNAME3217(G3217,G3215,G3216);
  nor GNAME3218(G3218,G20209,G2851);
  and GNAME3219(G3219,G3215,G3218);
  nor GNAME3220(G3220,G2851,G2853);
  and GNAME3221(G3221,G3215,G3220);
  nor GNAME3222(G3222,G20180,G2849);
  nor GNAME3223(G3223,G20209,G20233);
  and GNAME3224(G3224,G3222,G3223);
  and GNAME3225(G3225,G3216,G3222);
  and GNAME3226(G3226,G3218,G3222);
  and GNAME3227(G3227,G3220,G3222);
  nor GNAME3228(G3228,G20141,G2847);
  and GNAME3229(G3229,G3223,G3228);
  and GNAME3230(G3230,G3216,G3228);
  and GNAME3231(G3231,G3218,G3228);
  and GNAME3232(G3232,G3220,G3228);
  nor GNAME3233(G3233,G2847,G2849);
  and GNAME3234(G3234,G3223,G3233);
  and GNAME3235(G3235,G3216,G3233);
  and GNAME3236(G3236,G3218,G3233);
  and GNAME3237(G3237,G3220,G3233);
  and GNAME3238(G3238,G3215,G3223);
  and GNAME3239(G3239,G20108,G2799,G2794);
  and GNAME3240(G3240,G2746,G2795);
  and GNAME3241(G3241,G58979,G2825);
  and GNAME3242(G3242,G7446,G2866);
  and GNAME3243(G3243,G7971,G7972,G7449,G2896);
  and GNAME3244(G3244,G7467,G2875);
  and GNAME3245(G3245,G2866,G7508);
  and GNAME3246(G3246,G3798,G3802);
  and GNAME3247(G3247,G58979,G4322);
  nand GNAME3248(G3248,G3111,G2785,G2749);
  nor GNAME3249(G3249,G3954,G3835,G3852);
  and GNAME3250(G3250,G7818,G3111);
  nor GNAME3251(G3251,G58976,G7805);
  nand GNAME3252(G3252,G7848,G7849);
  nand GNAME3253(G3253,G7874,G7875);
  nand GNAME3254(G3254,G7877,G7878);
  nand GNAME3255(G3255,G7880,G7881);
  nand GNAME3256(G3256,G7887,G7888);
  nand GNAME3257(G3257,G7899,G7900);
  nand GNAME3258(G3258,G7896,G7897);
  nand GNAME3259(G3259,G7930,G7931);
  nand GNAME3260(G3260,G7836,G7837);
  nand GNAME3261(G3261,G7838,G7839);
  nand GNAME3262(G3262,G7840,G7841);
  nand GNAME3263(G3263,G7844,G7845);
  nand GNAME3264(G3264,G7851,G7852);
  nand GNAME3265(G3265,G7883,G7884);
  nand GNAME3266(G3266,G7890,G7891);
  nand GNAME3267(G3267,G7893,G7894);
  nand GNAME3268(G3268,G7902,G7903);
  nand GNAME3269(G3269,G7906,G7907);
  nand GNAME3270(G3270,G7908,G7909);
  nand GNAME3271(G3271,G7914,G7915);
  nand GNAME3272(G3272,G7916,G7917);
  nand GNAME3273(G3273,G7922,G7923);
  nand GNAME3274(G3274,G7924,G7925);
  nand GNAME3275(G3275,G7926,G7927);
  nand GNAME3276(G3276,G7928,G7929);
  nand GNAME3277(G3277,G7935,G7936);
  nand GNAME3278(G3278,G7937,G7938);
  nand GNAME3279(G3279,G7939,G7940);
  nand GNAME3280(G3280,G7941,G7942);
  nand GNAME3281(G3281,G7943,G7944);
  nand GNAME3282(G3282,G7945,G7946);
  nand GNAME3283(G3283,G7947,G7948);
  nand GNAME3284(G3284,G7949,G7950);
  nand GNAME3285(G3285,G7951,G7952);
  nand GNAME3286(G3286,G7953,G7954);
  nand GNAME3287(G3287,G7955,G7956);
  nand GNAME3288(G3288,G7957,G7958);
  nand GNAME3289(G3289,G7959,G7960);
  nand GNAME3290(G3290,G7961,G7962);
  nand GNAME3291(G3291,G7963,G7964);
  nand GNAME3292(G3292,G7965,G7966);
  nand GNAME3293(G3293,G7967,G7968);
  and GNAME3294(G3294,G3853,G3854,G3855,G3856);
  and GNAME3295(G3295,G3857,G3858,G3859,G3860);
  and GNAME3296(G3296,G3861,G3862,G3863,G3864);
  and GNAME3297(G3297,G3865,G3866,G3867,G3868);
  and GNAME3298(G3298,G3921,G3922,G3923,G3924);
  and GNAME3299(G3299,G3925,G3926,G3927,G3928);
  and GNAME3300(G3300,G3929,G3930,G3931,G3932);
  and GNAME3301(G3301,G3933,G3934,G3935,G3936);
  and GNAME3302(G3302,G3938,G3939,G3940,G3941);
  and GNAME3303(G3303,G3942,G3943,G3944,G3945);
  and GNAME3304(G3304,G3946,G3947,G3948,G3949);
  and GNAME3305(G3305,G3950,G3951,G3952,G3953);
  and GNAME3306(G3306,G3904,G3905,G3906,G3907);
  and GNAME3307(G3307,G3908,G3909,G3910,G3911);
  and GNAME3308(G3308,G3912,G3913,G3914,G3915);
  and GNAME3309(G3309,G3916,G3917,G3918,G3919);
  and GNAME3310(G3310,G3887,G3888,G3889,G3890);
  and GNAME3311(G3311,G3891,G3892,G3893,G3894);
  and GNAME3312(G3312,G3895,G3896,G3897,G3898);
  and GNAME3313(G3313,G3899,G3900,G3901,G3902);
  and GNAME3314(G3314,G3836,G3837,G3838,G3839);
  and GNAME3315(G3315,G3840,G3841,G3842,G3843);
  and GNAME3316(G3316,G3844,G3845,G3846,G3847);
  and GNAME3317(G3317,G3848,G3849,G3850,G3851);
  and GNAME3318(G3318,G3819,G3820,G3821,G3822);
  and GNAME3319(G3319,G3823,G3824,G3825,G3826);
  and GNAME3320(G3320,G3827,G3828,G3829,G3830);
  and GNAME3321(G3321,G3831,G3832,G3833,G3834);
  and GNAME3322(G3322,G3870,G3871,G3872,G3873);
  and GNAME3323(G3323,G3874,G3875,G3876,G3877);
  and GNAME3324(G3324,G3878,G3879,G3880,G3881);
  and GNAME3325(G3325,G3882,G3883,G3884,G3885);
  or GNAME3326(G3326,G58949,G58948,G58947,G58946);
  nor GNAME3327(G3327,G3326,G58950,G58951,G58952,G58953);
  or GNAME3328(G3328,G58957,G58956,G58955,G58954);
  nor GNAME3329(G3329,G3328,G58958,G58959,G58960,G58961);
  or GNAME3330(G3330,G58965,G58964,G58963,G58962);
  nor GNAME3331(G3331,G3330,G58966,G58967,G58968,G58969);
  or GNAME3332(G3332,G58973,G58972,G58971,G58970);
  nor GNAME3333(G3333,G3332,G4008,G58974,G58975);
  and GNAME3334(G3334,G4031,G4029,G4028);
  and GNAME3335(G3335,G4037,G4035,G4034);
  and GNAME3336(G3336,G4043,G4041,G4040);
  and GNAME3337(G3337,G4049,G4047,G4046);
  and GNAME3338(G3338,G4055,G4053,G4052);
  and GNAME3339(G3339,G4061,G4059,G4058);
  and GNAME3340(G3340,G4067,G4065,G4064);
  and GNAME3341(G3341,G4073,G4071,G4070);
  and GNAME3342(G3342,G4079,G4077,G4076);
  and GNAME3343(G3343,G4085,G4083,G4082);
  and GNAME3344(G3344,G4091,G4089,G4088);
  and GNAME3345(G3345,G4097,G4095,G4094);
  and GNAME3346(G3346,G4104,G4102,G4098);
  and GNAME3347(G3347,G4110,G4108,G4098);
  and GNAME3348(G3348,G4116,G4114,G4098);
  and GNAME3349(G3349,G4122,G4120,G4098);
  and GNAME3350(G3350,G4128,G4126,G4098);
  and GNAME3351(G3351,G4134,G4132,G4098);
  and GNAME3352(G3352,G4140,G4138,G4098);
  and GNAME3353(G3353,G4146,G4144,G4098);
  and GNAME3354(G3354,G4152,G4150,G4098);
  and GNAME3355(G3355,G4158,G4156,G4098);
  and GNAME3356(G3356,G4164,G4098,G4161);
  and GNAME3357(G3357,G4170,G4098,G4169);
  and GNAME3358(G3358,G4176,G4098,G4175);
  and GNAME3359(G3359,G4182,G4098,G4181);
  and GNAME3360(G3360,G4098,G4187,G4192,G4189);
  and GNAME3361(G3361,G4098,G4193,G4198,G4195);
  and GNAME3362(G3362,G4202,G4203);
  and GNAME3363(G3363,G4208,G4209);
  and GNAME3364(G3364,G4213,G4211,G4216);
  and GNAME3365(G3365,G4219,G4217,G4222);
  and GNAME3366(G3366,G4815,G4812,G4813);
  and GNAME3367(G3367,G3835,G2784,G3954);
  and GNAME3368(G3368,G4841,G4839,G4840);
  and GNAME3369(G3369,G7857,G7858,G7859,G7860);
  and GNAME3370(G3370,G4850,G4848,G4849);
  and GNAME3371(G3371,G4856,G4854,G4855);
  and GNAME3372(G3372,G4862,G4860,G4861);
  and GNAME3373(G3373,G4868,G4866,G4867);
  and GNAME3374(G3374,G4874,G4872,G4873);
  and GNAME3375(G3375,G4880,G4878,G4879);
  and GNAME3376(G3376,G4886,G4884,G4885);
  and GNAME3377(G3377,G4892,G4890,G4891);
  and GNAME3378(G3378,G4898,G4896,G4897);
  and GNAME3379(G3379,G4904,G4902,G4903);
  and GNAME3380(G3380,G4910,G4908,G4909);
  and GNAME3381(G3381,G4916,G4914,G4915);
  and GNAME3382(G3382,G4922,G4920,G4921);
  and GNAME3383(G3383,G4928,G4926,G4927);
  and GNAME3384(G3384,G4934,G4932,G4933);
  and GNAME3385(G3385,G4940,G4938,G4939);
  and GNAME3386(G3386,G4946,G4944,G4945);
  and GNAME3387(G3387,G4952,G4950,G4951);
  and GNAME3388(G3388,G4958,G4956,G4957);
  and GNAME3389(G3389,G4964,G4962,G4963);
  and GNAME3390(G3390,G4970,G4968,G4969);
  and GNAME3391(G3391,G4976,G4974,G4975);
  and GNAME3392(G3392,G4982,G4980,G4981);
  and GNAME3393(G3393,G4988,G4986,G4987);
  and GNAME3394(G3394,G4994,G4992,G4993);
  and GNAME3395(G3395,G5000,G4998,G4999);
  and GNAME3396(G3396,G5006,G5004,G5005);
  and GNAME3397(G3397,G5012,G5010,G5011);
  and GNAME3398(G3398,G5018,G5016,G5021);
  and GNAME3399(G3399,G5024,G5022,G5027);
  and GNAME3400(G3400,G5030,G5028,G5033);
  and GNAME3401(G3401,G5036,G5034,G5039);
  and GNAME3402(G3402,G7872,G7873);
  and GNAME3403(G3403,G7885,G7886);
  and GNAME3404(G3404,G5132,G5130,G5127);
  and GNAME3405(G3405,G5153,G5149,G5152);
  and GNAME3406(G3406,G5181,G5177,G5180);
  and GNAME3407(G3407,G5207,G5205,G5206);
  and GNAME3408(G3408,G5216,G5214,G5215);
  and GNAME3409(G3409,G5225,G5223,G5224);
  and GNAME3410(G3410,G5234,G5232,G5233);
  and GNAME3411(G3411,G5243,G5241,G5242);
  and GNAME3412(G3412,G5252,G5250,G5251);
  and GNAME3413(G3413,G5261,G5259,G5260);
  and GNAME3414(G3414,G5270,G5268,G5269);
  and GNAME3415(G3415,G5289,G5287,G5288);
  and GNAME3416(G3416,G5295,G5293,G5294);
  and GNAME3417(G3417,G5301,G5299,G5300);
  and GNAME3418(G3418,G5307,G5305,G5306);
  and GNAME3419(G3419,G5313,G5311,G5312);
  and GNAME3420(G3420,G5319,G5317,G5318);
  and GNAME3421(G3421,G5325,G5323,G5324);
  and GNAME3422(G3422,G5331,G5329,G5330);
  and GNAME3423(G3423,G5350,G5348,G5349);
  and GNAME3424(G3424,G5356,G5354,G5355);
  and GNAME3425(G3425,G5362,G5360,G5361);
  and GNAME3426(G3426,G5368,G5366,G5367);
  and GNAME3427(G3427,G5374,G5372,G5373);
  and GNAME3428(G3428,G5380,G5378,G5379);
  and GNAME3429(G3429,G5386,G5384,G5385);
  and GNAME3430(G3430,G5392,G5390,G5391);
  and GNAME3431(G3431,G5411,G5409,G5410);
  and GNAME3432(G3432,G5417,G5415,G5416);
  and GNAME3433(G3433,G5423,G5421,G5422);
  and GNAME3434(G3434,G5429,G5427,G5428);
  and GNAME3435(G3435,G5435,G5433,G5434);
  and GNAME3436(G3436,G5441,G5439,G5440);
  and GNAME3437(G3437,G5447,G5445,G5446);
  and GNAME3438(G3438,G5453,G5451,G5452);
  and GNAME3439(G3439,G5472,G5470,G5471);
  and GNAME3440(G3440,G5478,G5476,G5477);
  and GNAME3441(G3441,G5484,G5482,G5483);
  and GNAME3442(G3442,G5490,G5488,G5489);
  and GNAME3443(G3443,G5496,G5494,G5495);
  and GNAME3444(G3444,G5502,G5500,G5501);
  and GNAME3445(G3445,G5508,G5506,G5507);
  and GNAME3446(G3446,G5514,G5512,G5513);
  and GNAME3447(G3447,G5533,G5531,G5532);
  and GNAME3448(G3448,G5539,G5537,G5538);
  and GNAME3449(G3449,G5545,G5543,G5544);
  and GNAME3450(G3450,G5551,G5549,G5550);
  and GNAME3451(G3451,G5557,G5555,G5556);
  and GNAME3452(G3452,G5563,G5561,G5562);
  and GNAME3453(G3453,G5569,G5567,G5568);
  and GNAME3454(G3454,G5575,G5573,G5574);
  and GNAME3455(G3455,G5594,G5592,G5593);
  and GNAME3456(G3456,G5600,G5598,G5599);
  and GNAME3457(G3457,G5606,G5604,G5605);
  and GNAME3458(G3458,G5612,G5610,G5611);
  and GNAME3459(G3459,G5618,G5616,G5617);
  and GNAME3460(G3460,G5624,G5622,G5623);
  and GNAME3461(G3461,G5630,G5628,G5629);
  and GNAME3462(G3462,G5636,G5634,G5635);
  and GNAME3463(G3463,G5655,G5653,G5654);
  and GNAME3464(G3464,G5661,G5659,G5660);
  and GNAME3465(G3465,G5667,G5665,G5666);
  and GNAME3466(G3466,G5673,G5671,G5672);
  and GNAME3467(G3467,G5679,G5677,G5678);
  and GNAME3468(G3468,G5685,G5683,G5684);
  and GNAME3469(G3469,G5691,G5689,G5690);
  and GNAME3470(G3470,G5697,G5695,G5696);
  and GNAME3471(G3471,G5716,G5714,G5715);
  and GNAME3472(G3472,G5722,G5720,G5721);
  and GNAME3473(G3473,G5728,G5726,G5727);
  and GNAME3474(G3474,G5734,G5732,G5733);
  and GNAME3475(G3475,G5740,G5738,G5739);
  and GNAME3476(G3476,G5746,G5744,G5745);
  and GNAME3477(G3477,G5752,G5750,G5751);
  and GNAME3478(G3478,G5758,G5756,G5757);
  and GNAME3479(G3479,G5777,G5775,G5776);
  and GNAME3480(G3480,G5783,G5781,G5782);
  and GNAME3481(G3481,G5789,G5787,G5788);
  and GNAME3482(G3482,G5795,G5793,G5794);
  and GNAME3483(G3483,G5801,G5799,G5800);
  and GNAME3484(G3484,G5807,G5805,G5806);
  and GNAME3485(G3485,G5813,G5811,G5812);
  and GNAME3486(G3486,G5819,G5817,G5818);
  and GNAME3487(G3487,G5838,G5836,G5837);
  and GNAME3488(G3488,G5844,G5842,G5843);
  and GNAME3489(G3489,G5850,G5848,G5849);
  and GNAME3490(G3490,G5856,G5854,G5855);
  and GNAME3491(G3491,G5862,G5860,G5861);
  and GNAME3492(G3492,G5868,G5866,G5867);
  and GNAME3493(G3493,G5874,G5872,G5873);
  and GNAME3494(G3494,G5880,G5878,G5879);
  and GNAME3495(G3495,G5899,G5897,G5898);
  and GNAME3496(G3496,G5905,G5903,G5904);
  and GNAME3497(G3497,G5911,G5909,G5910);
  and GNAME3498(G3498,G5917,G5915,G5916);
  and GNAME3499(G3499,G5923,G5921,G5922);
  and GNAME3500(G3500,G5929,G5927,G5928);
  and GNAME3501(G3501,G5935,G5933,G5934);
  and GNAME3502(G3502,G5941,G5939,G5940);
  and GNAME3503(G3503,G5960,G5958,G5959);
  and GNAME3504(G3504,G5966,G5964,G5965);
  and GNAME3505(G3505,G5972,G5970,G5971);
  and GNAME3506(G3506,G5978,G5976,G5977);
  and GNAME3507(G3507,G5984,G5982,G5983);
  and GNAME3508(G3508,G5990,G5988,G5989);
  and GNAME3509(G3509,G5996,G5994,G5995);
  and GNAME3510(G3510,G6002,G6000,G6001);
  and GNAME3511(G3511,G6021,G6019,G6020);
  and GNAME3512(G3512,G6027,G6025,G6026);
  and GNAME3513(G3513,G6033,G6031,G6032);
  and GNAME3514(G3514,G6039,G6037,G6038);
  and GNAME3515(G3515,G6045,G6043,G6044);
  and GNAME3516(G3516,G6051,G6049,G6050);
  and GNAME3517(G3517,G6057,G6055,G6056);
  and GNAME3518(G3518,G6063,G6061,G6062);
  and GNAME3519(G3519,G6082,G6080,G6081);
  and GNAME3520(G3520,G6088,G6086,G6087);
  and GNAME3521(G3521,G6094,G6092,G6093);
  and GNAME3522(G3522,G6100,G6098,G6099);
  and GNAME3523(G3523,G6106,G6104,G6105);
  and GNAME3524(G3524,G6112,G6110,G6111);
  and GNAME3525(G3525,G6118,G6116,G6117);
  and GNAME3526(G3526,G6124,G6122,G6123);
  and GNAME3527(G3527,G6143,G6141,G6142);
  and GNAME3528(G3528,G6149,G6147,G6148);
  and GNAME3529(G3529,G6155,G6153,G6154);
  and GNAME3530(G3530,G6161,G6159,G6160);
  and GNAME3531(G3531,G6167,G6165,G6166);
  and GNAME3532(G3532,G6173,G6171,G6172);
  and GNAME3533(G3533,G6179,G6177,G6178);
  and GNAME3534(G3534,G6185,G6183,G6184);
  nand GNAME3535(G3535,G20786,G6188,G6189);
  and GNAME3536(G3536,G6309,G6310,G6311,G6312);
  and GNAME3537(G3537,G6313,G6314,G6315,G6316);
  and GNAME3538(G3538,G6317,G6318,G6319,G6320);
  and GNAME3539(G3539,G6321,G6322,G6323,G6324);
  and GNAME3540(G3540,G6325,G6326,G6327,G6328);
  and GNAME3541(G3541,G6329,G6330,G6331,G6332);
  and GNAME3542(G3542,G6333,G6334,G6335,G6336);
  and GNAME3543(G3543,G6337,G6338,G6339,G6340);
  and GNAME3544(G3544,G6341,G6342,G6343,G6344);
  and GNAME3545(G3545,G6345,G6346,G6347,G6348);
  and GNAME3546(G3546,G6349,G6350,G6351,G6352);
  and GNAME3547(G3547,G6353,G6354,G6355,G6356);
  and GNAME3548(G3548,G6357,G6358,G6359,G6360);
  and GNAME3549(G3549,G6361,G6362,G6363,G6364);
  and GNAME3550(G3550,G6365,G6366,G6367,G6368);
  and GNAME3551(G3551,G6369,G6370,G6371,G6372);
  and GNAME3552(G3552,G6373,G6374,G6375,G6376);
  and GNAME3553(G3553,G6377,G6378,G6379,G6380);
  and GNAME3554(G3554,G6381,G6382,G6383,G6384);
  and GNAME3555(G3555,G6385,G6386,G6387,G6388);
  and GNAME3556(G3556,G6389,G6390,G6391,G6392);
  and GNAME3557(G3557,G6393,G6394,G6395,G6396);
  and GNAME3558(G3558,G6397,G6398,G6399,G6400);
  and GNAME3559(G3559,G6401,G6402,G6403,G6404);
  and GNAME3560(G3560,G6405,G6406,G6407,G6408);
  and GNAME3561(G3561,G6409,G6410,G6411,G6412);
  and GNAME3562(G3562,G6413,G6414,G6415,G6416);
  and GNAME3563(G3563,G6417,G6418,G6419,G6420);
  and GNAME3564(G3564,G6421,G6422,G6423,G6424);
  and GNAME3565(G3565,G6425,G6426,G6427,G6428);
  and GNAME3566(G3566,G6429,G6430,G6431,G6432);
  and GNAME3567(G3567,G6433,G6434,G6435,G6436);
  and GNAME3568(G3568,G6438,G6439,G6440,G6441);
  and GNAME3569(G3569,G6442,G6443,G6444,G6445);
  and GNAME3570(G3570,G6446,G6447,G6448,G6449);
  and GNAME3571(G3571,G6450,G6451,G6452,G6453);
  and GNAME3572(G3572,G6454,G6455,G6456,G6457);
  and GNAME3573(G3573,G6458,G6459,G6460,G6461);
  and GNAME3574(G3574,G6462,G6463,G6464,G6465);
  and GNAME3575(G3575,G6466,G6467,G6468,G6469);
  and GNAME3576(G3576,G6470,G6471,G6472,G6473);
  and GNAME3577(G3577,G6474,G6475,G6476,G6477);
  and GNAME3578(G3578,G6478,G6479,G6480,G6481);
  and GNAME3579(G3579,G6482,G6483,G6484,G6485);
  and GNAME3580(G3580,G6486,G6487,G6488,G6489);
  and GNAME3581(G3581,G6490,G6491,G6492,G6493);
  and GNAME3582(G3582,G6494,G6495,G6496,G6497);
  and GNAME3583(G3583,G6498,G6499,G6500,G6501);
  and GNAME3584(G3584,G6502,G6503,G6504,G6505);
  and GNAME3585(G3585,G6506,G6507,G6508,G6509);
  and GNAME3586(G3586,G6510,G6511,G6512,G6513);
  and GNAME3587(G3587,G6514,G6515,G6516,G6517);
  and GNAME3588(G3588,G6518,G6519,G6520,G6521);
  and GNAME3589(G3589,G6522,G6523,G6524,G6525);
  and GNAME3590(G3590,G6526,G6527,G6528,G6529);
  and GNAME3591(G3591,G6530,G6531,G6532,G6533);
  and GNAME3592(G3592,G6534,G6535,G6536,G6537);
  and GNAME3593(G3593,G6538,G6539,G6540,G6541);
  and GNAME3594(G3594,G6542,G6543,G6544,G6545);
  and GNAME3595(G3595,G6546,G6547,G6548,G6549);
  and GNAME3596(G3596,G6550,G6551,G6552,G6553);
  and GNAME3597(G3597,G6554,G6555,G6556,G6557);
  and GNAME3598(G3598,G6558,G6559,G6560,G6561);
  and GNAME3599(G3599,G6562,G6563,G6564,G6565);
  and GNAME3600(G3600,G6566,G6567,G6568,G6569);
  and GNAME3601(G3601,G6570,G6571,G6572,G6573);
  and GNAME3602(G3602,G6574,G6575,G6576,G6577);
  and GNAME3603(G3603,G6578,G6579,G6580,G6581);
  and GNAME3604(G3604,G6583,G6584,G6585,G6586);
  and GNAME3605(G3605,G6587,G6588,G6589,G6590);
  and GNAME3606(G3606,G6591,G6592,G6593,G6594);
  and GNAME3607(G3607,G6595,G6596,G6597,G6598);
  and GNAME3608(G3608,G6600,G6601,G6602,G6603);
  and GNAME3609(G3609,G6604,G6605,G6606,G6607);
  and GNAME3610(G3610,G6608,G6609,G6610,G6611);
  and GNAME3611(G3611,G6612,G6613,G6614,G6615);
  and GNAME3612(G3612,G6617,G6618,G6619,G6620);
  and GNAME3613(G3613,G6621,G6622,G6623,G6624);
  and GNAME3614(G3614,G6625,G6626,G6627,G6628);
  and GNAME3615(G3615,G6629,G6630,G6631,G6632);
  and GNAME3616(G3616,G6634,G6635,G6636,G6637);
  and GNAME3617(G3617,G6638,G6639,G6640,G6641);
  and GNAME3618(G3618,G6642,G6643,G6644,G6645);
  and GNAME3619(G3619,G6646,G6647,G6648,G6649);
  and GNAME3620(G3620,G6651,G6652,G6653,G6654);
  and GNAME3621(G3621,G6655,G6656,G6657,G6658);
  and GNAME3622(G3622,G6659,G6660,G6661,G6662);
  and GNAME3623(G3623,G6663,G6664,G6665,G6666);
  and GNAME3624(G3624,G6668,G6669,G6670,G6671);
  and GNAME3625(G3625,G6672,G6673,G6674,G6675);
  and GNAME3626(G3626,G6676,G6677,G6678,G6679);
  and GNAME3627(G3627,G6680,G6681,G6682,G6683);
  and GNAME3628(G3628,G6685,G6686,G6687,G6688);
  and GNAME3629(G3629,G6689,G6690,G6691,G6692);
  and GNAME3630(G3630,G6693,G6694,G6695,G6696);
  and GNAME3631(G3631,G6697,G6698,G6699,G6700);
  and GNAME3632(G3632,G6702,G6703,G6704,G6705);
  and GNAME3633(G3633,G6706,G6707,G6708,G6709);
  and GNAME3634(G3634,G6710,G6711,G6712,G6713);
  and GNAME3635(G3635,G6714,G6715,G6716,G6717);
  and GNAME3636(G3636,G6719,G6720,G6721,G6722);
  and GNAME3637(G3637,G6723,G6724,G6725,G6726);
  and GNAME3638(G3638,G6727,G6728,G6729,G6730);
  and GNAME3639(G3639,G6731,G6732,G6733,G6734);
  and GNAME3640(G3640,G6736,G6737,G6738,G6739);
  and GNAME3641(G3641,G6740,G6741,G6742,G6743);
  and GNAME3642(G3642,G6744,G6745,G6746,G6747);
  and GNAME3643(G3643,G6748,G6749,G6750,G6751);
  and GNAME3644(G3644,G6753,G6754,G6755,G6756);
  and GNAME3645(G3645,G6757,G6758,G6759,G6760);
  and GNAME3646(G3646,G6761,G6762,G6763,G6764);
  and GNAME3647(G3647,G6765,G6766,G6767,G6768);
  and GNAME3648(G3648,G6770,G6771,G6772,G6773);
  and GNAME3649(G3649,G6774,G6775,G6776,G6777);
  and GNAME3650(G3650,G6778,G6779,G6780,G6781);
  and GNAME3651(G3651,G6782,G6783,G6784,G6785);
  and GNAME3652(G3652,G6787,G6788,G6789,G6790);
  and GNAME3653(G3653,G6791,G6792,G6793,G6794);
  and GNAME3654(G3654,G6795,G6796,G6797,G6798);
  and GNAME3655(G3655,G6799,G6800,G6801,G6802);
  and GNAME3656(G3656,G6804,G6805,G6806,G6807);
  and GNAME3657(G3657,G6808,G6809,G6810,G6811);
  and GNAME3658(G3658,G6812,G6813,G6814,G6815);
  and GNAME3659(G3659,G6816,G6817,G6818,G6819);
  and GNAME3660(G3660,G6821,G6822,G6823,G6824);
  and GNAME3661(G3661,G6825,G6826,G6827,G6828);
  and GNAME3662(G3662,G6829,G6830,G6831,G6832);
  and GNAME3663(G3663,G6833,G6834,G6835,G6836);
  and GNAME3664(G3664,G3886,G6997,G6998);
  and GNAME3665(G3665,G7033,G7034,G7035,G7036);
  and GNAME3666(G3666,G7037,G7038,G7039,G7040);
  and GNAME3667(G3667,G7041,G7042,G7043,G7044);
  and GNAME3668(G3668,G7045,G7046,G7047,G7048);
  and GNAME3669(G3669,G7016,G7017,G7018,G7019);
  and GNAME3670(G3670,G7020,G7021,G7022,G7023);
  and GNAME3671(G3671,G7024,G7025,G7026,G7027);
  and GNAME3672(G3672,G7028,G7029,G7030,G7031);
  and GNAME3673(G3673,G6999,G7000,G7001,G7002);
  and GNAME3674(G3674,G7003,G7004,G7005,G7006);
  and GNAME3675(G3675,G7007,G7008,G7009,G7010);
  and GNAME3676(G3676,G7011,G7012,G7013,G7014);
  and GNAME3677(G3677,G7088,G7089,G7090,G7091);
  and GNAME3678(G3678,G7092,G7093,G7094,G7095);
  and GNAME3679(G3679,G7096,G7097,G7098,G7099);
  and GNAME3680(G3680,G7100,G7101,G7102,G7103);
  and GNAME3681(G3681,G7071,G7072,G7073,G7074);
  and GNAME3682(G3682,G7075,G7076,G7077,G7078);
  and GNAME3683(G3683,G7079,G7080,G7081,G7082);
  and GNAME3684(G3684,G7083,G7084,G7085,G7086);
  and GNAME3685(G3685,G7054,G7055,G7056,G7057);
  and GNAME3686(G3686,G7058,G7059,G7060,G7061);
  and GNAME3687(G3687,G7062,G7063,G7064,G7065);
  and GNAME3688(G3688,G7066,G7067,G7068,G7069);
  and GNAME3689(G3689,G7143,G7144,G7145,G7146);
  and GNAME3690(G3690,G7147,G7148,G7149,G7150);
  and GNAME3691(G3691,G7151,G7152,G7153,G7154);
  and GNAME3692(G3692,G7155,G7156,G7157,G7158);
  and GNAME3693(G3693,G7126,G7127,G7128,G7129);
  and GNAME3694(G3694,G7130,G7131,G7132,G7133);
  and GNAME3695(G3695,G7134,G7135,G7136,G7137);
  and GNAME3696(G3696,G7138,G7139,G7140,G7141);
  and GNAME3697(G3697,G7109,G7110,G7111,G7112);
  and GNAME3698(G3698,G7113,G7114,G7115,G7116);
  and GNAME3699(G3699,G7117,G7118,G7119,G7120);
  and GNAME3700(G3700,G7121,G7122,G7123,G7124);
  and GNAME3701(G3701,G7198,G7199,G7200,G7201);
  and GNAME3702(G3702,G7202,G7203,G7204,G7205);
  and GNAME3703(G3703,G7206,G7207,G7208,G7209);
  and GNAME3704(G3704,G7210,G7211,G7212,G7213);
  and GNAME3705(G3705,G7181,G7182,G7183,G7184);
  and GNAME3706(G3706,G7185,G7186,G7187,G7188);
  and GNAME3707(G3707,G7189,G7190,G7191,G7192);
  and GNAME3708(G3708,G7193,G7194,G7195,G7196);
  and GNAME3709(G3709,G7164,G7165,G7166,G7167);
  and GNAME3710(G3710,G7168,G7169,G7170,G7171);
  and GNAME3711(G3711,G7172,G7173,G7174,G7175);
  and GNAME3712(G3712,G7176,G7177,G7178,G7179);
  and GNAME3713(G3713,G7254,G7255,G7256,G7257);
  and GNAME3714(G3714,G7258,G7259,G7260,G7261);
  and GNAME3715(G3715,G7262,G7263,G7264,G7265);
  and GNAME3716(G3716,G7266,G7267,G7268,G7269);
  and GNAME3717(G3717,G7237,G7238,G7239,G7240);
  and GNAME3718(G3718,G7241,G7242,G7243,G7244);
  and GNAME3719(G3719,G7245,G7246,G7247,G7248);
  and GNAME3720(G3720,G7249,G7250,G7251,G7252);
  and GNAME3721(G3721,G7220,G7221,G7222,G7223);
  and GNAME3722(G3722,G7224,G7225,G7226,G7227);
  and GNAME3723(G3723,G7228,G7229,G7230,G7231);
  and GNAME3724(G3724,G7232,G7233,G7234,G7235);
  and GNAME3725(G3725,G7310,G7311,G7312,G7313);
  and GNAME3726(G3726,G7314,G7315,G7316,G7317);
  and GNAME3727(G3727,G7318,G7319,G7320,G7321);
  and GNAME3728(G3728,G7322,G7323,G7324,G7325);
  and GNAME3729(G3729,G7293,G7294,G7295,G7296);
  and GNAME3730(G3730,G7297,G7298,G7299,G7300);
  and GNAME3731(G3731,G7301,G7302,G7303,G7304);
  and GNAME3732(G3732,G7305,G7306,G7307,G7308);
  and GNAME3733(G3733,G7276,G7277,G7278,G7279);
  and GNAME3734(G3734,G7280,G7281,G7282,G7283);
  and GNAME3735(G3735,G7284,G7285,G7286,G7287);
  and GNAME3736(G3736,G7288,G7289,G7290,G7291);
  and GNAME3737(G3737,G7331,G7329,G7330);
  and GNAME3738(G3738,G7366,G7367,G7368,G7369);
  and GNAME3739(G3739,G7370,G7371,G7372,G7373);
  and GNAME3740(G3740,G7374,G7375,G7376,G7377);
  and GNAME3741(G3741,G7378,G7379,G7380,G7381);
  and GNAME3742(G3742,G7349,G7350,G7351,G7352);
  and GNAME3743(G3743,G7353,G7354,G7355,G7356);
  and GNAME3744(G3744,G7357,G7358,G7359,G7360);
  and GNAME3745(G3745,G7361,G7362,G7363,G7364);
  and GNAME3746(G3746,G7332,G7333,G7334,G7335);
  and GNAME3747(G3747,G7336,G7337,G7338,G7339);
  and GNAME3748(G3748,G7340,G7341,G7342,G7343);
  and GNAME3749(G3749,G7344,G7345,G7346,G7347);
  and GNAME3750(G3750,G7387,G7385,G7386);
  and GNAME3751(G3751,G7422,G7423,G7424,G7425);
  and GNAME3752(G3752,G7426,G7427,G7428,G7429);
  and GNAME3753(G3753,G7430,G7431,G7432,G7433);
  and GNAME3754(G3754,G7434,G7435,G7436,G7437);
  and GNAME3755(G3755,G7405,G7406,G7407,G7408);
  and GNAME3756(G3756,G7409,G7410,G7411,G7412);
  and GNAME3757(G3757,G7413,G7414,G7415,G7416);
  and GNAME3758(G3758,G7417,G7418,G7419,G7420);
  and GNAME3759(G3759,G7388,G7389,G7390,G7391);
  and GNAME3760(G3760,G7392,G7393,G7394,G7395);
  and GNAME3761(G3761,G7396,G7397,G7398,G7399);
  and GNAME3762(G3762,G7400,G7401,G7402,G7403);
  and GNAME3763(G3763,G7443,G7441,G7442);
  and GNAME3764(G3764,G7447,G7448);
  and GNAME3765(G3765,G3818,G2855,G7450,G7969);
  and GNAME3766(G3766,G7463,G7461,G7462);
  and GNAME3767(G3767,G7621,G7619,G7620);
  and GNAME3768(G3768,G7672,G7673,G7677,G7674,G7670);
  and GNAME3769(G3769,G7731,G7732,G7736,G7733,G7729);
  and GNAME3770(G3770,G7790,G7791,G7795,G7792,G7788);
  and GNAME3771(G3771,G7799,G7800,G7804,G7801,G7797);
  or GNAME3772(G3772,G2813,G2806);
  and GNAME3773(G3773,G7983,G3975,G3977);
  not GNAME3774(G3774,G35);
  or GNAME3775(G3775,G2927,G2928);
  and GNAME3776(G3776,G5076,G5074,G5075);
  nand GNAME3777(G3777,G5088,G3816,G2912);
  nand GNAME3778(G3778,G5090,G58977);
  and GNAME3779(G3779,G2762,G3869);
  nand GNAME3780(G3780,G2762,G7898);
  nand GNAME3781(G3781,G2891,G5086,G5087);
  not GNAME3782(G3782,G2859);
  not GNAME3783(G3783,G3246);
  not GNAME3784(G3784,G2746);
  not GNAME3785(G3785,G2748);
  not GNAME3786(G3786,G2787);
  not GNAME3787(G3787,G2814);
  not GNAME3788(G3788,G3114);
  not GNAME3789(G3789,G3115);
  not GNAME3790(G3790,G2762);
  not GNAME3791(G3791,G2772);
  not GNAME3792(G3792,G2827);
  not GNAME3793(G3793,G2830);
  not GNAME3794(G3794,G2829);
  not GNAME3795(G3795,G2831);
  not GNAME3796(G3796,G2828);
  not GNAME3797(G3797,G2910);
  not GNAME3798(G3798,G2943);
  not GNAME3799(G3799,G2836);
  not GNAME3800(G3800,G2805);
  not GNAME3801(G3801,G2793);
  not GNAME3802(G3802,G2816);
  nand GNAME3803(G3803,G2913,G2836);
  not GNAME3804(G3804,G2922);
  not GNAME3805(G3805,G2823);
  not GNAME3806(G3806,G2890);
  not GNAME3807(G3807,G2803);
  not GNAME3808(G3808,G2856);
  not GNAME3809(G3809,G2942);
  nand GNAME3810(G3810,G3241,G2799,G20108);
  or GNAME3811(G3811,G58944,G58945,G59309,G7988);
  nand GNAME3812(G3812,G2900,G3979,G58979);
  nand GNAME3813(G3813,G1590,G2842);
  nand GNAME3814(G3814,G2836,G2754,G2790);
  nand GNAME3815(G3815,G58976,G58979,G2805);
  nand GNAME3816(G3816,G59346,G2911);
  nand GNAME3817(G3817,G2820,G2815);
  not GNAME3818(G3818,G2897);
  nand GNAME3819(G3819,G59094,G2758);
  nand GNAME3820(G3820,G59086,G2761);
  nand GNAME3821(G3821,G59078,G2763);
  nand GNAME3822(G3822,G59070,G2767);
  nand GNAME3823(G3823,G59062,G2768);
  nand GNAME3824(G3824,G59054,G2769);
  nand GNAME3825(G3825,G59046,G2770);
  nand GNAME3826(G3826,G59038,G2773);
  nand GNAME3827(G3827,G59030,G2774);
  nand GNAME3828(G3828,G59022,G2775);
  nand GNAME3829(G3829,G59014,G2776);
  nand GNAME3830(G3830,G59006,G2778);
  nand GNAME3831(G3831,G58998,G2779);
  nand GNAME3832(G3832,G58990,G2780);
  nand GNAME3833(G3833,G58982,G2781);
  nand GNAME3834(G3834,G2782,G59102);
  not GNAME3835(G3835,G2783);
  nand GNAME3836(G3836,G2782,G59106);
  nand GNAME3837(G3837,G2758,G59098);
  nand GNAME3838(G3838,G2761,G59090);
  nand GNAME3839(G3839,G2763,G59082);
  nand GNAME3840(G3840,G2767,G59074);
  nand GNAME3841(G3841,G2768,G59066);
  nand GNAME3842(G3842,G2769,G59058);
  nand GNAME3843(G3843,G2770,G59050);
  nand GNAME3844(G3844,G2773,G59042);
  nand GNAME3845(G3845,G2774,G59034);
  nand GNAME3846(G3846,G2775,G59026);
  nand GNAME3847(G3847,G2776,G59018);
  nand GNAME3848(G3848,G2778,G59010);
  nand GNAME3849(G3849,G2779,G59002);
  nand GNAME3850(G3850,G2780,G58994);
  nand GNAME3851(G3851,G2781,G58986);
  not GNAME3852(G3852,G2799);
  nand GNAME3853(G3853,G2782,G59107);
  nand GNAME3854(G3854,G2758,G59099);
  nand GNAME3855(G3855,G2761,G59091);
  nand GNAME3856(G3856,G2763,G59083);
  nand GNAME3857(G3857,G2767,G59075);
  nand GNAME3858(G3858,G2768,G59067);
  nand GNAME3859(G3859,G2769,G59059);
  nand GNAME3860(G3860,G2770,G59051);
  nand GNAME3861(G3861,G2773,G59043);
  nand GNAME3862(G3862,G2774,G59035);
  nand GNAME3863(G3863,G2775,G59027);
  nand GNAME3864(G3864,G2776,G59019);
  nand GNAME3865(G3865,G2778,G59011);
  nand GNAME3866(G3866,G2779,G59003);
  nand GNAME3867(G3867,G2780,G58995);
  nand GNAME3868(G3868,G2781,G58987);
  not GNAME3869(G3869,G2795);
  nand GNAME3870(G3870,G2782,G59105);
  nand GNAME3871(G3871,G2758,G59097);
  nand GNAME3872(G3872,G2761,G59089);
  nand GNAME3873(G3873,G2763,G59081);
  nand GNAME3874(G3874,G2767,G59073);
  nand GNAME3875(G3875,G2768,G59065);
  nand GNAME3876(G3876,G2769,G59057);
  nand GNAME3877(G3877,G2770,G59049);
  nand GNAME3878(G3878,G2773,G59041);
  nand GNAME3879(G3879,G2774,G59033);
  nand GNAME3880(G3880,G2775,G59025);
  nand GNAME3881(G3881,G2776,G59017);
  nand GNAME3882(G3882,G2778,G59009);
  nand GNAME3883(G3883,G2779,G59001);
  nand GNAME3884(G3884,G2780,G58993);
  nand GNAME3885(G3885,G2781,G58985);
  not GNAME3886(G3886,G2784);
  nand GNAME3887(G3887,G2758,G59095);
  nand GNAME3888(G3888,G2761,G59087);
  nand GNAME3889(G3889,G2763,G59079);
  nand GNAME3890(G3890,G2767,G59071);
  nand GNAME3891(G3891,G2768,G59063);
  nand GNAME3892(G3892,G2769,G59055);
  nand GNAME3893(G3893,G2770,G59047);
  nand GNAME3894(G3894,G2773,G59039);
  nand GNAME3895(G3895,G2774,G59031);
  nand GNAME3896(G3896,G2775,G59023);
  nand GNAME3897(G3897,G2776,G59015);
  nand GNAME3898(G3898,G2778,G59007);
  nand GNAME3899(G3899,G2779,G58999);
  nand GNAME3900(G3900,G2780,G58991);
  nand GNAME3901(G3901,G2781,G58983);
  nand GNAME3902(G3902,G2782,G59103);
  not GNAME3903(G3903,G2786);
  nand GNAME3904(G3904,G2758,G59093);
  nand GNAME3905(G3905,G2761,G59085);
  nand GNAME3906(G3906,G2763,G59077);
  nand GNAME3907(G3907,G2767,G59069);
  nand GNAME3908(G3908,G2768,G59061);
  nand GNAME3909(G3909,G2769,G59053);
  nand GNAME3910(G3910,G2770,G59045);
  nand GNAME3911(G3911,G2773,G59037);
  nand GNAME3912(G3912,G2774,G59029);
  nand GNAME3913(G3913,G2775,G59021);
  nand GNAME3914(G3914,G2776,G59013);
  nand GNAME3915(G3915,G2778,G59005);
  nand GNAME3916(G3916,G2779,G58997);
  nand GNAME3917(G3917,G2780,G58989);
  nand GNAME3918(G3918,G2781,G58981);
  nand GNAME3919(G3919,G2782,G59101);
  not GNAME3920(G3920,G2785);
  nand GNAME3921(G3921,G2758,G59092);
  nand GNAME3922(G3922,G2761,G59084);
  nand GNAME3923(G3923,G2763,G59076);
  nand GNAME3924(G3924,G2767,G59068);
  nand GNAME3925(G3925,G2768,G59060);
  nand GNAME3926(G3926,G2769,G59052);
  nand GNAME3927(G3927,G2770,G59044);
  nand GNAME3928(G3928,G2773,G59036);
  nand GNAME3929(G3929,G2774,G59028);
  nand GNAME3930(G3930,G2775,G59020);
  nand GNAME3931(G3931,G2776,G59012);
  nand GNAME3932(G3932,G2778,G59004);
  nand GNAME3933(G3933,G2779,G58996);
  nand GNAME3934(G3934,G2780,G58988);
  nand GNAME3935(G3935,G2781,G58980);
  nand GNAME3936(G3936,G2782,G59100);
  not GNAME3937(G3937,G2855);
  nand GNAME3938(G3938,G2758,G59096);
  nand GNAME3939(G3939,G2761,G59088);
  nand GNAME3940(G3940,G2763,G59080);
  nand GNAME3941(G3941,G2767,G59072);
  nand GNAME3942(G3942,G2768,G59064);
  nand GNAME3943(G3943,G2769,G59056);
  nand GNAME3944(G3944,G2770,G59048);
  nand GNAME3945(G3945,G2773,G59040);
  nand GNAME3946(G3946,G2774,G59032);
  nand GNAME3947(G3947,G2775,G59024);
  nand GNAME3948(G3948,G2776,G59016);
  nand GNAME3949(G3949,G2778,G59008);
  nand GNAME3950(G3950,G2779,G59000);
  nand GNAME3951(G3951,G2780,G58992);
  nand GNAME3952(G3952,G2781,G58984);
  nand GNAME3953(G3953,G2782,G59104);
  not GNAME3954(G3954,G2749);
  not GNAME3955(G3955,G2789);
  not GNAME3956(G3956,G2791);
  nand GNAME3957(G3957,G2798,G58977,G7989);
  not GNAME3958(G3958,G2802);
  nand GNAME3959(G3959,G3957,G2880);
  nand GNAME3960(G3960,G3959,G20108);
  nand GNAME3961(G3961,G58977,G3869);
  or GNAME3962(G3962,G2754,G2746,G2788);
  nor GNAME3963(G3963,G2808,G2809);
  not GNAME3964(G3964,G2810);
  nand GNAME3965(G3965,G58943,G59353);
  nand GNAME3966(G3966,G2796,G3954,G3869);
  nand GNAME3967(G3967,G3966,G2784);
  nand GNAME3968(G3968,G2792,G2799);
  nand GNAME3969(G3969,G2787,G3968,G3835);
  nand GNAME3970(G3970,G2804,G7849);
  nand GNAME3971(G3971,G3969,G3886);
  nand GNAME3972(G3972,G2803,G2812);
  nand GNAME3973(G3973,G3972,G59352);
  nand GNAME3974(G3974,G58979,G2813);
  or GNAME3975(G3975,G1590,G2818);
  nand GNAME3976(G3976,G58977,G58979);
  nand GNAME3977(G3977,G3976,G2819);
  nand GNAME3978(G3978,G2807,G58941);
  nand GNAME3979(G3979,G3978,G2808);
  not GNAME3980(G3980,G2821);
  nand GNAME3981(G3981,G2821,G3869);
  nand GNAME3982(G3982,G2799,G3981);
  nand GNAME3983(G3983,G3980,G59348);
  nand GNAME3984(G3984,G3982,G3983);
  nand GNAME3985(G3985,G3984,G58977);
  nand GNAME3986(G3986,G3869,G2823);
  nand GNAME3987(G3987,G3985,G3986);
  nand GNAME3988(G3988,G2752,G3987);
  nand GNAME3989(G3989,G3988,G58979);
  and GNAME3990(G3990,G3800,G3989);
  nand GNAME3991(G3991,G2821,G7850);
  nand GNAME3992(G3992,G2752,G3991);
  or GNAME3993(G3993,G3107,G3807);
  not GNAME3994(G3994,G2867);
  nand GNAME3995(G3995,G3994,G3782);
  nand GNAME3996(G3996,G3995,G2793);
  nand GNAME3997(G3997,G3996,G3957,G2880);
  nand GNAME3998(G3998,G2825,G58977,G2798);
  nand GNAME3999(G3999,G2791,G2793);
  nand GNAME4000(G4000,G3998,G3999);
  nand GNAME4001(G4001,G2792,G4000);
  nand GNAME4002(G4002,G2804,G3997);
  and GNAME4003(G4003,G4001,G4002);
  or GNAME4004(G4004,G3107,G4003);
  nand GNAME4005(G4005,G3993,G59347);
  nand GNAME4006(G4006,G58977,G20773,G2798,G2825);
  nand GNAME4007(G4007,G3993,G59346);
  and GNAME4008(G4008,G58945,G58944);
  nand GNAME4009(G4009,G7988,G59343);
  and GNAME4010(G4010,G58944,G59309);
  or GNAME4011(G4011,G4010,G2834);
  or GNAME4012(G4012,G2833,G2835);
  nand GNAME4013(G4013,G7988,G59342);
  nand GNAME4014(G4014,G7988,G59341);
  not GNAME4015(G4015,G2845);
  not GNAME4016(G4016,G2838);
  nand GNAME4017(G4017,G2839,G2830,G2838);
  nand GNAME4018(G4018,G20210,G2845,G58978);
  nand GNAME4019(G4019,G4016,G2830,G2839,G3285);
  or GNAME4020(G4020,G2817,G20210,G4015);
  nand GNAME4021(G4021,G4019,G4020);
  nand GNAME4022(G4022,G3980,G2838);
  nand GNAME4023(G4023,G2830,G2841,G4016);
  nand GNAME4024(G4024,G4022,G2800);
  nand GNAME4025(G4025,G4023,G4024);
  nand GNAME4026(G4026,G2840,G59308);
  nand GNAME4027(G4027,G4021,G20210);
  nand GNAME4028(G4028,G59181,G2843);
  nand GNAME4029(G4029,G2846,G20508);
  nand GNAME4030(G4030,G20921,G2844);
  nand GNAME4031(G4031,G4015,G59340);
  nand GNAME4032(G4032,G2840,G59307);
  nand GNAME4033(G4033,G4021,G20142);
  nand GNAME4034(G4034,G2843,G59180);
  nand GNAME4035(G4035,G2846,G20447);
  nand GNAME4036(G4036,G2844,G20922);
  nand GNAME4037(G4037,G4015,G59339);
  nand GNAME4038(G4038,G2840,G59306);
  nand GNAME4039(G4039,G4021,G20196);
  nand GNAME4040(G4040,G2843,G59179);
  nand GNAME4041(G4041,G2846,G20495);
  nand GNAME4042(G4042,G2844,G20960);
  nand GNAME4043(G4043,G4015,G59338);
  nand GNAME4044(G4044,G2840,G59305);
  nand GNAME4045(G4045,G4021,G20197);
  nand GNAME4046(G4046,G2843,G59178);
  nand GNAME4047(G4047,G2846,G20496);
  nand GNAME4048(G4048,G2844,G20961);
  nand GNAME4049(G4049,G4015,G59337);
  nand GNAME4050(G4050,G2840,G59304);
  nand GNAME4051(G4051,G4021,G20198);
  nand GNAME4052(G4052,G2843,G59177);
  nand GNAME4053(G4053,G2846,G20497);
  nand GNAME4054(G4054,G2844,G20962);
  nand GNAME4055(G4055,G4015,G59336);
  nand GNAME4056(G4056,G2840,G59303);
  nand GNAME4057(G4057,G4021,G20199);
  nand GNAME4058(G4058,G2843,G59176);
  nand GNAME4059(G4059,G2846,G20498);
  nand GNAME4060(G4060,G2844,G20963);
  nand GNAME4061(G4061,G4015,G59335);
  nand GNAME4062(G4062,G2840,G59302);
  nand GNAME4063(G4063,G4021,G20200);
  nand GNAME4064(G4064,G2843,G59175);
  nand GNAME4065(G4065,G2846,G20499);
  nand GNAME4066(G4066,G2844,G20964);
  nand GNAME4067(G4067,G4015,G59334);
  nand GNAME4068(G4068,G2840,G59301);
  nand GNAME4069(G4069,G4021,G20201);
  nand GNAME4070(G4070,G2843,G59174);
  nand GNAME4071(G4071,G2846,G20537);
  nand GNAME4072(G4072,G2844,G20965);
  nand GNAME4073(G4073,G4015,G59333);
  nand GNAME4074(G4074,G2840,G59300);
  nand GNAME4075(G4075,G4021,G20202);
  nand GNAME4076(G4076,G2843,G59173);
  nand GNAME4077(G4077,G2846,G20540);
  nand GNAME4078(G4078,G2844,G20966);
  nand GNAME4079(G4079,G4015,G59332);
  nand GNAME4080(G4080,G2840,G59299);
  nand GNAME4081(G4081,G4021,G20203);
  nand GNAME4082(G4082,G2843,G59172);
  nand GNAME4083(G4083,G2846,G20543);
  nand GNAME4084(G4084,G2844,G20967);
  nand GNAME4085(G4085,G4015,G59331);
  nand GNAME4086(G4086,G2840,G59298);
  nand GNAME4087(G4087,G4021,G20204);
  nand GNAME4088(G4088,G2843,G59171);
  nand GNAME4089(G4089,G2846,G20546);
  nand GNAME4090(G4090,G2844,G20968);
  nand GNAME4091(G4091,G4015,G59330);
  nand GNAME4092(G4092,G2840,G59297);
  nand GNAME4093(G4093,G4021,G20205);
  nand GNAME4094(G4094,G2843,G59170);
  nand GNAME4095(G4095,G2846,G20549);
  nand GNAME4096(G4096,G2844,G20969);
  nand GNAME4097(G4097,G4015,G59329);
  nand GNAME4098(G4098,G2845,G2790,G2817);
  nand GNAME4099(G4099,G2840,G59296);
  nand GNAME4100(G4100,G4021,G20206);
  nand GNAME4101(G4101,G2843,G59169);
  nand GNAME4102(G4102,G2846,G20555);
  nand GNAME4103(G4103,G2844,G20973);
  nand GNAME4104(G4104,G4015,G59328);
  nand GNAME4105(G4105,G2840,G59295);
  nand GNAME4106(G4106,G4021,G20207);
  nand GNAME4107(G4107,G2843,G59168);
  nand GNAME4108(G4108,G2846,G20558);
  nand GNAME4109(G4109,G2844,G20974);
  nand GNAME4110(G4110,G4015,G59327);
  nand GNAME4111(G4111,G2840,G59294);
  nand GNAME4112(G4112,G4021,G20208);
  nand GNAME4113(G4113,G2843,G59167);
  nand GNAME4114(G4114,G2846,G20561);
  nand GNAME4115(G4115,G2844,G20975);
  nand GNAME4116(G4116,G4015,G59326);
  nand GNAME4117(G4117,G2840,G59293);
  nand GNAME4118(G4118,G4021,G20236);
  nand GNAME4119(G4119,G2843,G59166);
  nand GNAME4120(G4120,G2846,G20500);
  nand GNAME4121(G4121,G2844,G20976);
  nand GNAME4122(G4122,G4015,G59325);
  nand GNAME4123(G4123,G2840,G59292);
  nand GNAME4124(G4124,G4021,G20239);
  nand GNAME4125(G4125,G2843,G59165);
  nand GNAME4126(G4126,G2846,G20501);
  nand GNAME4127(G4127,G2844,G20977);
  nand GNAME4128(G4128,G4015,G59324);
  nand GNAME4129(G4129,G2840,G59291);
  nand GNAME4130(G4130,G4021,G20211);
  nand GNAME4131(G4131,G2843,G59164);
  nand GNAME4132(G4132,G2846,G20445);
  nand GNAME4133(G4133,G2844,G20923);
  nand GNAME4134(G4134,G4015,G59323);
  nand GNAME4135(G4135,G2840,G59290);
  nand GNAME4136(G4136,G4021,G20243);
  nand GNAME4137(G4137,G2843,G59163);
  nand GNAME4138(G4138,G2846,G20502);
  nand GNAME4139(G4139,G2844,G20978);
  nand GNAME4140(G4140,G4015,G59322);
  nand GNAME4141(G4141,G2840,G59289);
  nand GNAME4142(G4142,G4021,G20246);
  nand GNAME4143(G4143,G2843,G59162);
  nand GNAME4144(G4144,G2846,G20503);
  nand GNAME4145(G4145,G2844,G20979);
  nand GNAME4146(G4146,G4015,G59321);
  nand GNAME4147(G4147,G2840,G59288);
  nand GNAME4148(G4148,G4021,G20212);
  nand GNAME4149(G4149,G2843,G59161);
  nand GNAME4150(G4150,G2846,G20504);
  nand GNAME4151(G4151,G2844,G20859);
  nand GNAME4152(G4152,G4015,G59320);
  nand GNAME4153(G4153,G2840,G59287);
  nand GNAME4154(G4154,G4021,G20140);
  nand GNAME4155(G4155,G2843,G59160);
  nand GNAME4156(G4156,G2846,G20444);
  nand GNAME4157(G4157,G2844,G20858);
  nand GNAME4158(G4158,G4015,G59319);
  nand GNAME4159(G4159,G2840,G59286);
  nand GNAME4160(G4160,G4021,G20219);
  nand GNAME4161(G4161,G2843,G59159);
  nand GNAME4162(G4162,G2846,G20481);
  nand GNAME4163(G4163,G2844,G20950);
  nand GNAME4164(G4164,G4015,G59318);
  nand GNAME4165(G4165,G2840,G59285);
  nand GNAME4166(G4166,G4021,G20176);
  nand GNAME4167(G4167,G2843,G59158);
  nand GNAME4168(G4168,G2846,G20516);
  nand GNAME4169(G4169,G2844,G20951);
  nand GNAME4170(G4170,G4015,G59317);
  nand GNAME4171(G4171,G2840,G59284);
  nand GNAME4172(G4172,G4021,G20177);
  nand GNAME4173(G4173,G2843,G59157);
  nand GNAME4174(G4174,G2846,G20506);
  nand GNAME4175(G4175,G2844,G20919);
  nand GNAME4176(G4176,G4015,G59316);
  nand GNAME4177(G4177,G2840,G59283);
  nand GNAME4178(G4178,G4021,G20143);
  nand GNAME4179(G4179,G2843,G59156);
  nand GNAME4180(G4180,G2846,G20448);
  nand GNAME4181(G4181,G2844,G20861);
  nand GNAME4182(G4182,G4015,G59315);
  and GNAME4183(G4183,G2839,G2799,G2785);
  or GNAME4184(G4184,G4183,G2846);
  and GNAME4185(G4185,G2823,G2785,G2845);
  or GNAME4186(G4186,G4185,G2844);
  nand GNAME4187(G4187,G2840,G59282);
  nand GNAME4188(G4188,G4021,G20178);
  nand GNAME4189(G4189,G4186,G20955);
  nand GNAME4190(G4190,G2843,G59155);
  nand GNAME4191(G4191,G4184,G20520);
  nand GNAME4192(G4192,G4015,G59314);
  nand GNAME4193(G4193,G2840,G59281);
  nand GNAME4194(G4194,G4021,G20179);
  nand GNAME4195(G4195,G4186,G20958);
  nand GNAME4196(G4196,G2843,G59154);
  nand GNAME4197(G4197,G4184,G20523);
  nand GNAME4198(G4198,G4015,G59313);
  nand GNAME4199(G4199,G2840,G59280);
  nand GNAME4200(G4200,G4021,G20180);
  nand GNAME4201(G4201,G4186,G20920);
  nand GNAME4202(G4202,G2843,G59153);
  nand GNAME4203(G4203,G4015,G59312);
  nand GNAME4204(G4204,G4184,G20507);
  nand GNAME4205(G4205,G2840,G59279);
  nand GNAME4206(G4206,G4021,G20141);
  nand GNAME4207(G4207,G4186,G20860);
  nand GNAME4208(G4208,G2843,G59152);
  nand GNAME4209(G4209,G4015,G59311);
  nand GNAME4210(G4210,G4184,G20446);
  nand GNAME4211(G4211,G2840,G59278);
  nand GNAME4212(G4212,G4021,G20233);
  nand GNAME4213(G4213,G4186,G20972);
  nand GNAME4214(G4214,G2843,G59151);
  nand GNAME4215(G4215,G4184,G20552);
  nand GNAME4216(G4216,G59310,G4015);
  nand GNAME4217(G4217,G2840,G59277);
  nand GNAME4218(G4218,G4021,G20209);
  nand GNAME4219(G4219,G4186,G20918);
  nand GNAME4220(G4220,G2843,G59150);
  nand GNAME4221(G4221,G4184,G20505);
  nand GNAME4222(G4222,G59309,G4015);
  not GNAME4223(G4223,G2858);
  nand GNAME4224(G4224,G58979,G4223);
  nand GNAME4225(G4225,G20108,G2859);
  nand GNAME4226(G4226,G4224,G4225);
  nand GNAME4227(G4227,G2860,G59308);
  nand GNAME4228(G4228,G20210,G2861);
  nand GNAME4229(G4229,G2860,G59307);
  nand GNAME4230(G4230,G20447,G2862);
  nand GNAME4231(G4231,G20142,G2861);
  nand GNAME4232(G4232,G2860,G59306);
  nand GNAME4233(G4233,G20495,G2862);
  nand GNAME4234(G4234,G20196,G2861);
  nand GNAME4235(G4235,G2860,G59305);
  nand GNAME4236(G4236,G20496,G2862);
  nand GNAME4237(G4237,G20197,G2861);
  nand GNAME4238(G4238,G2860,G59304);
  nand GNAME4239(G4239,G20497,G2862);
  nand GNAME4240(G4240,G20198,G2861);
  nand GNAME4241(G4241,G2860,G59303);
  nand GNAME4242(G4242,G20498,G2862);
  nand GNAME4243(G4243,G20199,G2861);
  nand GNAME4244(G4244,G2860,G59302);
  nand GNAME4245(G4245,G20499,G2862);
  nand GNAME4246(G4246,G20200,G2861);
  nand GNAME4247(G4247,G2860,G59301);
  nand GNAME4248(G4248,G20537,G2862);
  nand GNAME4249(G4249,G20201,G2861);
  nand GNAME4250(G4250,G2860,G59300);
  nand GNAME4251(G4251,G20540,G2862);
  nand GNAME4252(G4252,G20202,G2861);
  nand GNAME4253(G4253,G2860,G59299);
  nand GNAME4254(G4254,G20543,G2862);
  nand GNAME4255(G4255,G20203,G2861);
  nand GNAME4256(G4256,G2860,G59298);
  nand GNAME4257(G4257,G20546,G2862);
  nand GNAME4258(G4258,G20204,G2861);
  nand GNAME4259(G4259,G2860,G59297);
  nand GNAME4260(G4260,G20549,G2862);
  nand GNAME4261(G4261,G20205,G2861);
  nand GNAME4262(G4262,G2860,G59296);
  nand GNAME4263(G4263,G20555,G2862);
  nand GNAME4264(G4264,G20206,G2861);
  nand GNAME4265(G4265,G2860,G59295);
  nand GNAME4266(G4266,G20558,G2862);
  nand GNAME4267(G4267,G20207,G2861);
  nand GNAME4268(G4268,G2860,G59294);
  nand GNAME4269(G4269,G20561,G2862);
  nand GNAME4270(G4270,G20208,G2861);
  nand GNAME4271(G4271,G2860,G59293);
  nand GNAME4272(G4272,G20500,G2862);
  nand GNAME4273(G4273,G20236,G2861);
  nand GNAME4274(G4274,G2860,G59292);
  nand GNAME4275(G4275,G20501,G2862);
  nand GNAME4276(G4276,G20239,G2861);
  nand GNAME4277(G4277,G2860,G59291);
  nand GNAME4278(G4278,G20445,G2862);
  nand GNAME4279(G4279,G20211,G2861);
  nand GNAME4280(G4280,G2860,G59290);
  nand GNAME4281(G4281,G20502,G2862);
  nand GNAME4282(G4282,G20243,G2861);
  nand GNAME4283(G4283,G2860,G59289);
  nand GNAME4284(G4284,G20503,G2862);
  nand GNAME4285(G4285,G20246,G2861);
  nand GNAME4286(G4286,G2860,G59288);
  nand GNAME4287(G4287,G20504,G2862);
  nand GNAME4288(G4288,G20212,G2861);
  nand GNAME4289(G4289,G2860,G59287);
  nand GNAME4290(G4290,G20444,G2862);
  nand GNAME4291(G4291,G20140,G2861);
  nand GNAME4292(G4292,G2860,G59286);
  nand GNAME4293(G4293,G20481,G2862);
  nand GNAME4294(G4294,G20219,G2861);
  nand GNAME4295(G4295,G2860,G59285);
  nand GNAME4296(G4296,G20516,G2862);
  nand GNAME4297(G4297,G20176,G2861);
  nand GNAME4298(G4298,G2860,G59284);
  nand GNAME4299(G4299,G20506,G2862);
  nand GNAME4300(G4300,G20177,G2861);
  nand GNAME4301(G4301,G2860,G59283);
  nand GNAME4302(G4302,G20448,G2862);
  nand GNAME4303(G4303,G20143,G2861);
  nand GNAME4304(G4304,G2860,G59282);
  nand GNAME4305(G4305,G20520,G2862);
  nand GNAME4306(G4306,G20178,G2861);
  nand GNAME4307(G4307,G2860,G59281);
  nand GNAME4308(G4308,G20523,G2862);
  nand GNAME4309(G4309,G20179,G2861);
  nand GNAME4310(G4310,G2860,G59280);
  nand GNAME4311(G4311,G20180,G2861);
  nand GNAME4312(G4312,G20507,G2862);
  nand GNAME4313(G4313,G2860,G59279);
  nand GNAME4314(G4314,G20141,G2861);
  nand GNAME4315(G4315,G20446,G2862);
  nand GNAME4316(G4316,G2860,G59278);
  nand GNAME4317(G4317,G20552,G2862);
  nand GNAME4318(G4318,G20233,G2861);
  nand GNAME4319(G4319,G2860,G59277);
  nand GNAME4320(G4320,G20209,G2861);
  nand GNAME4321(G4321,G20505,G2862);
  not GNAME4322(G4322,G2864);
  not GNAME4323(G4323,G3247);
  not GNAME4324(G4324,G2865);
  or GNAME4325(G4325,G2804,G2866);
  nand GNAME4326(G4326,G2791,G20773);
  nand GNAME4327(G4327,G4325,G4326);
  nand GNAME4328(G4328,G2752,G4327);
  nand GNAME4329(G4329,G20108,G2867);
  nand GNAME4330(G4330,G4329,G4323,G4328);
  nand GNAME4331(G4331,G2868,G59276);
  nand GNAME4332(G4332,G20210,G2869);
  nand GNAME4333(G4333,G2870,G58902);
  nand GNAME4334(G4334,G58885,G2871);
  nand GNAME4335(G4335,G2868,G59275);
  nand GNAME4336(G4336,G20142,G2869);
  nand GNAME4337(G4337,G20922,G2872);
  nand GNAME4338(G4338,G2870,G58901);
  nand GNAME4339(G4339,G2871,G58884);
  nand GNAME4340(G4340,G2868,G59274);
  nand GNAME4341(G4341,G20196,G2869);
  nand GNAME4342(G4342,G20960,G2872);
  nand GNAME4343(G4343,G2870,G58900);
  nand GNAME4344(G4344,G2871,G58883);
  nand GNAME4345(G4345,G2868,G59273);
  nand GNAME4346(G4346,G20197,G2869);
  nand GNAME4347(G4347,G20961,G2872);
  nand GNAME4348(G4348,G2870,G58899);
  nand GNAME4349(G4349,G2871,G58882);
  nand GNAME4350(G4350,G2868,G59272);
  nand GNAME4351(G4351,G20198,G2869);
  nand GNAME4352(G4352,G20962,G2872);
  nand GNAME4353(G4353,G2870,G58898);
  nand GNAME4354(G4354,G2871,G58881);
  nand GNAME4355(G4355,G2868,G59271);
  nand GNAME4356(G4356,G20199,G2869);
  nand GNAME4357(G4357,G20963,G2872);
  nand GNAME4358(G4358,G2870,G58897);
  nand GNAME4359(G4359,G2871,G58880);
  nand GNAME4360(G4360,G2868,G59270);
  nand GNAME4361(G4361,G20200,G2869);
  nand GNAME4362(G4362,G20964,G2872);
  nand GNAME4363(G4363,G2870,G58896);
  nand GNAME4364(G4364,G2871,G58879);
  nand GNAME4365(G4365,G2868,G59269);
  nand GNAME4366(G4366,G20201,G2869);
  nand GNAME4367(G4367,G20965,G2872);
  nand GNAME4368(G4368,G2870,G58895);
  nand GNAME4369(G4369,G2868,G59268);
  nand GNAME4370(G4370,G20202,G2869);
  nand GNAME4371(G4371,G20966,G2872);
  nand GNAME4372(G4372,G2870,G58894);
  nand GNAME4373(G4373,G2871,G58878);
  nand GNAME4374(G4374,G2868,G59267);
  nand GNAME4375(G4375,G20203,G2869);
  nand GNAME4376(G4376,G20967,G2872);
  nand GNAME4377(G4377,G2870,G58893);
  nand GNAME4378(G4378,G2871,G58877);
  nand GNAME4379(G4379,G2868,G59266);
  nand GNAME4380(G4380,G20204,G2869);
  nand GNAME4381(G4381,G20968,G2872);
  nand GNAME4382(G4382,G2870,G58892);
  nand GNAME4383(G4383,G2871,G58876);
  nand GNAME4384(G4384,G2868,G59265);
  nand GNAME4385(G4385,G20205,G2869);
  nand GNAME4386(G4386,G20969,G2872);
  nand GNAME4387(G4387,G2870,G58891);
  nand GNAME4388(G4388,G2871,G58875);
  nand GNAME4389(G4389,G2868,G59264);
  nand GNAME4390(G4390,G20206,G2869);
  nand GNAME4391(G4391,G20973,G2872);
  nand GNAME4392(G4392,G2870,G58890);
  nand GNAME4393(G4393,G2871,G58874);
  nand GNAME4394(G4394,G2868,G59263);
  nand GNAME4395(G4395,G20207,G2869);
  nand GNAME4396(G4396,G20974,G2872);
  nand GNAME4397(G4397,G2870,G58889);
  nand GNAME4398(G4398,G2871,G58873);
  nand GNAME4399(G4399,G2868,G59262);
  nand GNAME4400(G4400,G20208,G2869);
  nand GNAME4401(G4401,G20975,G2872);
  nand GNAME4402(G4402,G2870,G58888);
  nand GNAME4403(G4403,G2871,G58872);
  nand GNAME4404(G4404,G2868,G59261);
  nand GNAME4405(G4405,G20236,G2869);
  nand GNAME4406(G4406,G20976,G2872);
  nand GNAME4407(G4407,G2870,G58887);
  nand GNAME4408(G4408,G2871,G58871);
  nand GNAME4409(G4409,G58886,G2873);
  nand GNAME4410(G4410,G2868,G59260);
  nand GNAME4411(G4411,G20239,G2869);
  nand GNAME4412(G4412,G20977,G2872);
  nand GNAME4413(G4413,G58885,G2873);
  nand GNAME4414(G4414,G2868,G59259);
  nand GNAME4415(G4415,G20211,G2869);
  nand GNAME4416(G4416,G20923,G2872);
  nand GNAME4417(G4417,G58884,G2873);
  nand GNAME4418(G4418,G2868,G59258);
  nand GNAME4419(G4419,G20243,G2869);
  nand GNAME4420(G4420,G20978,G2872);
  nand GNAME4421(G4421,G58883,G2873);
  nand GNAME4422(G4422,G2868,G59257);
  nand GNAME4423(G4423,G20246,G2869);
  nand GNAME4424(G4424,G20979,G2872);
  nand GNAME4425(G4425,G58882,G2873);
  nand GNAME4426(G4426,G2868,G59256);
  nand GNAME4427(G4427,G20212,G2869);
  nand GNAME4428(G4428,G20859,G2872);
  nand GNAME4429(G4429,G58881,G2873);
  nand GNAME4430(G4430,G2868,G59255);
  nand GNAME4431(G4431,G20140,G2869);
  nand GNAME4432(G4432,G20858,G2872);
  nand GNAME4433(G4433,G58880,G2873);
  nand GNAME4434(G4434,G2868,G59254);
  nand GNAME4435(G4435,G20219,G2869);
  nand GNAME4436(G4436,G20950,G2872);
  nand GNAME4437(G4437,G58879,G2873);
  nand GNAME4438(G4438,G2868,G59253);
  nand GNAME4439(G4439,G20176,G2869);
  nand GNAME4440(G4440,G20951,G2872);
  nand GNAME4441(G4441,G2868,G59252);
  nand GNAME4442(G4442,G20177,G2869);
  nand GNAME4443(G4443,G20919,G2872);
  nand GNAME4444(G4444,G58878,G2873);
  nand GNAME4445(G4445,G2868,G59251);
  nand GNAME4446(G4446,G20143,G2869);
  nand GNAME4447(G4447,G20861,G2872);
  nand GNAME4448(G4448,G58877,G2873);
  nand GNAME4449(G4449,G2868,G59250);
  nand GNAME4450(G4450,G20178,G2869);
  nand GNAME4451(G4451,G20955,G2872);
  nand GNAME4452(G4452,G58876,G2873);
  nand GNAME4453(G4453,G2868,G59249);
  nand GNAME4454(G4454,G20179,G2869);
  nand GNAME4455(G4455,G20958,G2872);
  nand GNAME4456(G4456,G58875,G2873);
  nand GNAME4457(G4457,G2868,G59248);
  nand GNAME4458(G4458,G20920,G2872);
  nand GNAME4459(G4459,G20180,G2869);
  nand GNAME4460(G4460,G58874,G2873);
  nand GNAME4461(G4461,G2868,G59247);
  nand GNAME4462(G4462,G20860,G2872);
  nand GNAME4463(G4463,G20141,G2869);
  nand GNAME4464(G4464,G58873,G2873);
  nand GNAME4465(G4465,G2868,G59246);
  nand GNAME4466(G4466,G20972,G2872);
  nand GNAME4467(G4467,G20233,G2869);
  nand GNAME4468(G4468,G58872,G2873);
  nand GNAME4469(G4469,G2868,G59245);
  nand GNAME4470(G4470,G20918,G2872);
  nand GNAME4471(G4471,G20209,G2869);
  nand GNAME4472(G4472,G58871,G2873);
  not GNAME4473(G4473,G2874);
  nand GNAME4474(G4474,G2874,G58979,G3980);
  or GNAME4475(G4475,G58943,G2875);
  nand GNAME4476(G4476,G4474,G4475);
  nand GNAME4477(G4477,G20108,G4476,G2793);
  nand GNAME4478(G4478,G2876,G59243);
  nand GNAME4479(G4479,G59198,G2877);
  nand GNAME4480(G4480,G59275,G2879);
  nand GNAME4481(G4481,G2876,G59242);
  nand GNAME4482(G4482,G2877,G59199);
  nand GNAME4483(G4483,G59274,G2879);
  nand GNAME4484(G4484,G2876,G59241);
  nand GNAME4485(G4485,G2877,G59200);
  nand GNAME4486(G4486,G59273,G2879);
  nand GNAME4487(G4487,G2876,G59240);
  nand GNAME4488(G4488,G2877,G59201);
  nand GNAME4489(G4489,G59272,G2879);
  nand GNAME4490(G4490,G2876,G59239);
  nand GNAME4491(G4491,G2877,G59202);
  nand GNAME4492(G4492,G59271,G2879);
  nand GNAME4493(G4493,G2876,G59238);
  nand GNAME4494(G4494,G2877,G59203);
  nand GNAME4495(G4495,G59270,G2879);
  nand GNAME4496(G4496,G2876,G59237);
  nand GNAME4497(G4497,G2877,G59204);
  nand GNAME4498(G4498,G59269,G2879);
  nand GNAME4499(G4499,G2876,G59236);
  nand GNAME4500(G4500,G2877,G59205);
  nand GNAME4501(G4501,G59268,G2879);
  nand GNAME4502(G4502,G2876,G59235);
  nand GNAME4503(G4503,G2877,G59206);
  nand GNAME4504(G4504,G59267,G2879);
  nand GNAME4505(G4505,G2876,G59234);
  nand GNAME4506(G4506,G2877,G59207);
  nand GNAME4507(G4507,G59266,G2879);
  nand GNAME4508(G4508,G2876,G59233);
  nand GNAME4509(G4509,G2877,G59208);
  nand GNAME4510(G4510,G59265,G2879);
  nand GNAME4511(G4511,G2876,G59232);
  nand GNAME4512(G4512,G2877,G59209);
  nand GNAME4513(G4513,G59264,G2879);
  nand GNAME4514(G4514,G2876,G59231);
  nand GNAME4515(G4515,G2877,G59210);
  nand GNAME4516(G4516,G59263,G2879);
  nand GNAME4517(G4517,G2876,G59230);
  nand GNAME4518(G4518,G2877,G59211);
  nand GNAME4519(G4519,G59262,G2879);
  nand GNAME4520(G4520,G2876,G59229);
  nand GNAME4521(G4521,G2877,G59212);
  nand GNAME4522(G4522,G59261,G2879);
  nand GNAME4523(G4523,G2876,G59228);
  nand GNAME4524(G4524,G2877,G59182);
  nand GNAME4525(G4525,G59260,G2878);
  nand GNAME4526(G4526,G2876,G59227);
  nand GNAME4527(G4527,G2877,G59183);
  nand GNAME4528(G4528,G59259,G2878);
  nand GNAME4529(G4529,G2876,G59226);
  nand GNAME4530(G4530,G2877,G59184);
  nand GNAME4531(G4531,G59258,G2878);
  nand GNAME4532(G4532,G2876,G59225);
  nand GNAME4533(G4533,G2877,G59185);
  nand GNAME4534(G4534,G59257,G2878);
  nand GNAME4535(G4535,G2876,G59224);
  nand GNAME4536(G4536,G2877,G59186);
  nand GNAME4537(G4537,G59256,G2878);
  nand GNAME4538(G4538,G2876,G59223);
  nand GNAME4539(G4539,G2877,G59187);
  nand GNAME4540(G4540,G59255,G2878);
  nand GNAME4541(G4541,G2876,G59222);
  nand GNAME4542(G4542,G2877,G59188);
  nand GNAME4543(G4543,G59254,G2878);
  nand GNAME4544(G4544,G2876,G59221);
  nand GNAME4545(G4545,G2877,G59189);
  nand GNAME4546(G4546,G59253,G2878);
  nand GNAME4547(G4547,G2876,G59220);
  nand GNAME4548(G4548,G2877,G59190);
  nand GNAME4549(G4549,G59252,G2878);
  nand GNAME4550(G4550,G2876,G59219);
  nand GNAME4551(G4551,G2877,G59191);
  nand GNAME4552(G4552,G59251,G2878);
  nand GNAME4553(G4553,G2876,G59218);
  nand GNAME4554(G4554,G2877,G59192);
  nand GNAME4555(G4555,G59250,G2878);
  nand GNAME4556(G4556,G2876,G59217);
  nand GNAME4557(G4557,G2877,G59193);
  nand GNAME4558(G4558,G59249,G2878);
  nand GNAME4559(G4559,G2876,G59216);
  nand GNAME4560(G4560,G2877,G59194);
  nand GNAME4561(G4561,G59248,G2878);
  nand GNAME4562(G4562,G2876,G59215);
  nand GNAME4563(G4563,G2877,G59195);
  nand GNAME4564(G4564,G59247,G2878);
  nand GNAME4565(G4565,G2876,G59214);
  nand GNAME4566(G4566,G2877,G59196);
  nand GNAME4567(G4567,G59246,G2878);
  nand GNAME4568(G4568,G2876,G59213);
  nand GNAME4569(G4569,G2877,G59197);
  nand GNAME4570(G4570,G59245,G2878);
  or GNAME4571(G4571,G2804,G2880);
  or GNAME4572(G4572,G1590,G2881);
  nand GNAME4573(G4573,G59212,G2882);
  nand GNAME4574(G4574,G59261,G2883);
  nand GNAME4575(G4575,G59211,G2882);
  nand GNAME4576(G4576,G59262,G2883);
  nand GNAME4577(G4577,G59210,G2882);
  nand GNAME4578(G4578,G59263,G2883);
  nand GNAME4579(G4579,G59209,G2882);
  nand GNAME4580(G4580,G59264,G2883);
  nand GNAME4581(G4581,G59208,G2882);
  nand GNAME4582(G4582,G59265,G2883);
  nand GNAME4583(G4583,G59207,G2882);
  nand GNAME4584(G4584,G59266,G2883);
  nand GNAME4585(G4585,G59206,G2882);
  nand GNAME4586(G4586,G59267,G2883);
  nand GNAME4587(G4587,G59205,G2882);
  nand GNAME4588(G4588,G59268,G2883);
  nand GNAME4589(G4589,G59204,G2882);
  nand GNAME4590(G4590,G59269,G2883);
  nand GNAME4591(G4591,G59203,G2882);
  nand GNAME4592(G4592,G59270,G2883);
  nand GNAME4593(G4593,G59202,G2882);
  nand GNAME4594(G4594,G59271,G2883);
  nand GNAME4595(G4595,G59201,G2882);
  nand GNAME4596(G4596,G59272,G2883);
  nand GNAME4597(G4597,G59200,G2882);
  nand GNAME4598(G4598,G59273,G2883);
  nand GNAME4599(G4599,G59199,G2882);
  nand GNAME4600(G4600,G59274,G2883);
  nand GNAME4601(G4601,G59198,G2882);
  nand GNAME4602(G4602,G59275,G2883);
  nand GNAME4603(G4603,G59197,G2882);
  nand GNAME4604(G4604,G59245,G2883);
  nand GNAME4605(G4605,G58871,G2884);
  nand GNAME4606(G4606,G59196,G2882);
  nand GNAME4607(G4607,G59246,G2883);
  nand GNAME4608(G4608,G58872,G2884);
  nand GNAME4609(G4609,G59195,G2882);
  nand GNAME4610(G4610,G59247,G2883);
  nand GNAME4611(G4611,G58873,G2884);
  nand GNAME4612(G4612,G59194,G2882);
  nand GNAME4613(G4613,G59248,G2883);
  nand GNAME4614(G4614,G58874,G2884);
  nand GNAME4615(G4615,G59193,G2882);
  nand GNAME4616(G4616,G59249,G2883);
  nand GNAME4617(G4617,G58875,G2884);
  nand GNAME4618(G4618,G59192,G2882);
  nand GNAME4619(G4619,G59250,G2883);
  nand GNAME4620(G4620,G58876,G2884);
  nand GNAME4621(G4621,G59191,G2882);
  nand GNAME4622(G4622,G59251,G2883);
  nand GNAME4623(G4623,G58877,G2884);
  nand GNAME4624(G4624,G59190,G2882);
  nand GNAME4625(G4625,G59252,G2883);
  nand GNAME4626(G4626,G58878,G2884);
  nand GNAME4627(G4627,G58879,G2884);
  nand GNAME4628(G4628,G59189,G2882);
  nand GNAME4629(G4629,G59253,G2883);
  nand GNAME4630(G4630,G58880,G2884);
  nand GNAME4631(G4631,G59188,G2882);
  nand GNAME4632(G4632,G59254,G2883);
  nand GNAME4633(G4633,G58881,G2884);
  nand GNAME4634(G4634,G59187,G2882);
  nand GNAME4635(G4635,G59255,G2883);
  nand GNAME4636(G4636,G58882,G2884);
  nand GNAME4637(G4637,G59186,G2882);
  nand GNAME4638(G4638,G59256,G2883);
  nand GNAME4639(G4639,G58883,G2884);
  nand GNAME4640(G4640,G59185,G2882);
  nand GNAME4641(G4641,G59257,G2883);
  nand GNAME4642(G4642,G58884,G2884);
  nand GNAME4643(G4643,G59184,G2882);
  nand GNAME4644(G4644,G59258,G2883);
  nand GNAME4645(G4645,G58885,G2884);
  nand GNAME4646(G4646,G59183,G2882);
  nand GNAME4647(G4647,G59259,G2883);
  nand GNAME4648(G4648,G59182,G2882);
  nand GNAME4649(G4649,G58886,G2884);
  nand GNAME4650(G4650,G59260,G2883);
  nand GNAME4651(G4651,G2790,G2819);
  nand GNAME4652(G4652,G59181,G2885);
  nand GNAME4653(G4653,G20508,G2886);
  nand GNAME4654(G4654,G20210,G2887);
  nand GNAME4655(G4655,G20921,G2888);
  nand GNAME4656(G4656,G59340,G2889);
  nand GNAME4657(G4657,G59180,G2885);
  nand GNAME4658(G4658,G20447,G2886);
  nand GNAME4659(G4659,G20142,G2887);
  nand GNAME4660(G4660,G20922,G2888);
  nand GNAME4661(G4661,G59339,G2889);
  nand GNAME4662(G4662,G59179,G2885);
  nand GNAME4663(G4663,G20495,G2886);
  nand GNAME4664(G4664,G20196,G2887);
  nand GNAME4665(G4665,G20960,G2888);
  nand GNAME4666(G4666,G59338,G2889);
  nand GNAME4667(G4667,G59178,G2885);
  nand GNAME4668(G4668,G20496,G2886);
  nand GNAME4669(G4669,G20197,G2887);
  nand GNAME4670(G4670,G20961,G2888);
  nand GNAME4671(G4671,G59337,G2889);
  nand GNAME4672(G4672,G59177,G2885);
  nand GNAME4673(G4673,G20497,G2886);
  nand GNAME4674(G4674,G20198,G2887);
  nand GNAME4675(G4675,G20962,G2888);
  nand GNAME4676(G4676,G59336,G2889);
  nand GNAME4677(G4677,G59176,G2885);
  nand GNAME4678(G4678,G20498,G2886);
  nand GNAME4679(G4679,G20199,G2887);
  nand GNAME4680(G4680,G20963,G2888);
  nand GNAME4681(G4681,G59335,G2889);
  nand GNAME4682(G4682,G59175,G2885);
  nand GNAME4683(G4683,G20499,G2886);
  nand GNAME4684(G4684,G20200,G2887);
  nand GNAME4685(G4685,G20964,G2888);
  nand GNAME4686(G4686,G59334,G2889);
  nand GNAME4687(G4687,G59174,G2885);
  nand GNAME4688(G4688,G20537,G2886);
  nand GNAME4689(G4689,G20201,G2887);
  nand GNAME4690(G4690,G20965,G2888);
  nand GNAME4691(G4691,G59333,G2889);
  nand GNAME4692(G4692,G59173,G2885);
  nand GNAME4693(G4693,G20540,G2886);
  nand GNAME4694(G4694,G20202,G2887);
  nand GNAME4695(G4695,G20966,G2888);
  nand GNAME4696(G4696,G59332,G2889);
  nand GNAME4697(G4697,G59172,G2885);
  nand GNAME4698(G4698,G20543,G2886);
  nand GNAME4699(G4699,G20203,G2887);
  nand GNAME4700(G4700,G20967,G2888);
  nand GNAME4701(G4701,G59331,G2889);
  nand GNAME4702(G4702,G59171,G2885);
  nand GNAME4703(G4703,G20546,G2886);
  nand GNAME4704(G4704,G20204,G2887);
  nand GNAME4705(G4705,G20968,G2888);
  nand GNAME4706(G4706,G59330,G2889);
  nand GNAME4707(G4707,G59170,G2885);
  nand GNAME4708(G4708,G20549,G2886);
  nand GNAME4709(G4709,G20205,G2887);
  nand GNAME4710(G4710,G20969,G2888);
  nand GNAME4711(G4711,G59329,G2889);
  nand GNAME4712(G4712,G59169,G2885);
  nand GNAME4713(G4713,G20555,G2886);
  nand GNAME4714(G4714,G20206,G2887);
  nand GNAME4715(G4715,G20973,G2888);
  nand GNAME4716(G4716,G59328,G2889);
  nand GNAME4717(G4717,G59168,G2885);
  nand GNAME4718(G4718,G20558,G2886);
  nand GNAME4719(G4719,G20207,G2887);
  nand GNAME4720(G4720,G20974,G2888);
  nand GNAME4721(G4721,G59327,G2889);
  nand GNAME4722(G4722,G59167,G2885);
  nand GNAME4723(G4723,G20561,G2886);
  nand GNAME4724(G4724,G20208,G2887);
  nand GNAME4725(G4725,G20975,G2888);
  nand GNAME4726(G4726,G59326,G2889);
  nand GNAME4727(G4727,G59166,G2885);
  nand GNAME4728(G4728,G20500,G2886);
  nand GNAME4729(G4729,G20236,G2887);
  nand GNAME4730(G4730,G20976,G2888);
  nand GNAME4731(G4731,G59325,G2889);
  nand GNAME4732(G4732,G59165,G2885);
  nand GNAME4733(G4733,G20501,G2886);
  nand GNAME4734(G4734,G20239,G2887);
  nand GNAME4735(G4735,G20977,G2888);
  nand GNAME4736(G4736,G59324,G2889);
  nand GNAME4737(G4737,G59164,G2885);
  nand GNAME4738(G4738,G20445,G2886);
  nand GNAME4739(G4739,G20211,G2887);
  nand GNAME4740(G4740,G20923,G2888);
  nand GNAME4741(G4741,G59323,G2889);
  nand GNAME4742(G4742,G59163,G2885);
  nand GNAME4743(G4743,G20502,G2886);
  nand GNAME4744(G4744,G20243,G2887);
  nand GNAME4745(G4745,G20978,G2888);
  nand GNAME4746(G4746,G59322,G2889);
  nand GNAME4747(G4747,G59162,G2885);
  nand GNAME4748(G4748,G20503,G2886);
  nand GNAME4749(G4749,G20246,G2887);
  nand GNAME4750(G4750,G20979,G2888);
  nand GNAME4751(G4751,G59321,G2889);
  nand GNAME4752(G4752,G59161,G2885);
  nand GNAME4753(G4753,G20504,G2886);
  nand GNAME4754(G4754,G20212,G2887);
  nand GNAME4755(G4755,G20859,G2888);
  nand GNAME4756(G4756,G59320,G2889);
  nand GNAME4757(G4757,G59160,G2885);
  nand GNAME4758(G4758,G20444,G2886);
  nand GNAME4759(G4759,G20140,G2887);
  nand GNAME4760(G4760,G20858,G2888);
  nand GNAME4761(G4761,G59319,G2889);
  nand GNAME4762(G4762,G59159,G2885);
  nand GNAME4763(G4763,G20481,G2886);
  nand GNAME4764(G4764,G20219,G2887);
  nand GNAME4765(G4765,G20950,G2888);
  nand GNAME4766(G4766,G59318,G2889);
  nand GNAME4767(G4767,G59158,G2885);
  nand GNAME4768(G4768,G20516,G2886);
  nand GNAME4769(G4769,G20176,G2887);
  nand GNAME4770(G4770,G20951,G2888);
  nand GNAME4771(G4771,G59317,G2889);
  nand GNAME4772(G4772,G59157,G2885);
  nand GNAME4773(G4773,G20506,G2886);
  nand GNAME4774(G4774,G20177,G2887);
  nand GNAME4775(G4775,G20919,G2888);
  nand GNAME4776(G4776,G59316,G2889);
  nand GNAME4777(G4777,G59156,G2885);
  nand GNAME4778(G4778,G20448,G2886);
  nand GNAME4779(G4779,G20143,G2887);
  nand GNAME4780(G4780,G20861,G2888);
  nand GNAME4781(G4781,G59315,G2889);
  nand GNAME4782(G4782,G59155,G2885);
  nand GNAME4783(G4783,G20520,G2886);
  nand GNAME4784(G4784,G20178,G2887);
  nand GNAME4785(G4785,G20955,G2888);
  nand GNAME4786(G4786,G59314,G2889);
  nand GNAME4787(G4787,G59154,G2885);
  nand GNAME4788(G4788,G20523,G2886);
  nand GNAME4789(G4789,G20179,G2887);
  nand GNAME4790(G4790,G20958,G2888);
  nand GNAME4791(G4791,G59313,G2889);
  nand GNAME4792(G4792,G59153,G2885);
  nand GNAME4793(G4793,G20920,G2888);
  nand GNAME4794(G4794,G59312,G2889);
  nand GNAME4795(G4795,G20180,G2887);
  nand GNAME4796(G4796,G20507,G2886);
  nand GNAME4797(G4797,G59152,G2885);
  nand GNAME4798(G4798,G20860,G2888);
  nand GNAME4799(G4799,G59311,G2889);
  nand GNAME4800(G4800,G20141,G2887);
  nand GNAME4801(G4801,G20446,G2886);
  nand GNAME4802(G4802,G59151,G2885);
  nand GNAME4803(G4803,G20972,G2888);
  nand GNAME4804(G4804,G20552,G2886);
  nand GNAME4805(G4805,G20233,G2887);
  nand GNAME4806(G4806,G59310,G2889);
  nand GNAME4807(G4807,G59150,G2885);
  nand GNAME4808(G4808,G20918,G2888);
  nand GNAME4809(G4809,G20209,G2887);
  nand GNAME4810(G4810,G59309,G2889);
  nand GNAME4811(G4811,G20505,G2886);
  nand GNAME4812(G4812,G2783,G2787);
  nand GNAME4813(G4813,G3852,G2829);
  nand GNAME4814(G4814,G2786,G3852);
  nand GNAME4815(G4815,G4814,G2890);
  nand GNAME4816(G4816,G2786,G2785);
  nand GNAME4817(G4817,G3786,G3835);
  nand GNAME4818(G4818,G3903,G2752,G2799);
  nand GNAME4819(G4819,G4818,G3920);
  nand GNAME4820(G4820,G3835,G3980);
  nand GNAME4821(G4821,G4820,G3886);
  nand GNAME4822(G4822,G4821,G3852);
  nand GNAME4823(G4823,G2784,G3980);
  nand GNAME4824(G4824,G4822,G4823);
  nand GNAME4825(G4825,G2752,G4824);
  nand GNAME4826(G4826,G4825,G3903);
  nand GNAME4827(G4827,G20773,G4819,G3886);
  nand GNAME4828(G4828,G4826,G20108);
  nand GNAME4829(G4829,G2891,G4827,G4828);
  nand GNAME4830(G4830,G4829,G2803);
  nand GNAME4831(G4831,G2790,G2813);
  or GNAME4832(G4832,G2831,G2825,G2789,G4322);
  nand GNAME4833(G4833,G2894,G2786,G2800);
  or GNAME4834(G4834,G3903,G2753);
  nand GNAME4835(G4835,G4324,G4833,G4834,G2905);
  nand GNAME4836(G4836,G3252,G3937);
  nand GNAME4837(G4837,G2784,G2749);
  nand GNAME4838(G4838,G3903,G3784,G3954);
  nand GNAME4839(G4839,G4838,G3937);
  nand GNAME4840(G4840,G2784,G2826);
  nand GNAME4841(G4841,G3808,G2863);
  or GNAME4842(G4842,G2753,G2786);
  nand GNAME4843(G4843,G7973,G2856);
  nand GNAME4844(G4844,G4843,G3792);
  nand GNAME4845(G4845,G2795,G2899);
  nand GNAME4846(G4846,G3937,G2900);
  nand GNAME4847(G4847,G2902,G2903);
  nand GNAME4848(G4848,G21441,G2893);
  nand GNAME4849(G4849,G20508,G2904);
  nand GNAME4850(G4850,G20210,G2906);
  nand GNAME4851(G4851,G20921,G2907);
  nand GNAME4852(G4852,G59340,G2908);
  nand GNAME4853(G4853,G2909,G59149);
  nand GNAME4854(G4854,G2909,G59148);
  nand GNAME4855(G4855,G2893,G21442);
  nand GNAME4856(G4856,G20447,G2904);
  nand GNAME4857(G4857,G20142,G2906);
  nand GNAME4858(G4858,G20922,G2907);
  nand GNAME4859(G4859,G59339,G2908);
  nand GNAME4860(G4860,G2909,G59147);
  nand GNAME4861(G4861,G2893,G21393);
  nand GNAME4862(G4862,G20495,G2904);
  nand GNAME4863(G4863,G20196,G2906);
  nand GNAME4864(G4864,G20960,G2907);
  nand GNAME4865(G4865,G59338,G2908);
  nand GNAME4866(G4866,G2909,G59146);
  nand GNAME4867(G4867,G2893,G21392);
  nand GNAME4868(G4868,G20496,G2904);
  nand GNAME4869(G4869,G20197,G2906);
  nand GNAME4870(G4870,G20961,G2907);
  nand GNAME4871(G4871,G59337,G2908);
  nand GNAME4872(G4872,G2909,G59145);
  nand GNAME4873(G4873,G2893,G21444);
  nand GNAME4874(G4874,G20497,G2904);
  nand GNAME4875(G4875,G20198,G2906);
  nand GNAME4876(G4876,G20962,G2907);
  nand GNAME4877(G4877,G59336,G2908);
  nand GNAME4878(G4878,G2909,G59144);
  nand GNAME4879(G4879,G2893,G21391);
  nand GNAME4880(G4880,G20498,G2904);
  nand GNAME4881(G4881,G20199,G2906);
  nand GNAME4882(G4882,G20963,G2907);
  nand GNAME4883(G4883,G59335,G2908);
  nand GNAME4884(G4884,G2909,G59143);
  nand GNAME4885(G4885,G2893,G21390);
  nand GNAME4886(G4886,G20499,G2904);
  nand GNAME4887(G4887,G20200,G2906);
  nand GNAME4888(G4888,G20964,G2907);
  nand GNAME4889(G4889,G59334,G2908);
  nand GNAME4890(G4890,G2909,G59142);
  nand GNAME4891(G4891,G2893,G21468);
  nand GNAME4892(G4892,G20537,G2904);
  nand GNAME4893(G4893,G20201,G2906);
  nand GNAME4894(G4894,G20965,G2907);
  nand GNAME4895(G4895,G59333,G2908);
  nand GNAME4896(G4896,G2909,G59141);
  nand GNAME4897(G4897,G2893,G21469);
  nand GNAME4898(G4898,G20540,G2904);
  nand GNAME4899(G4899,G20202,G2906);
  nand GNAME4900(G4900,G20966,G2907);
  nand GNAME4901(G4901,G59332,G2908);
  nand GNAME4902(G4902,G2893,G21470);
  nand GNAME4903(G4903,G20543,G2904);
  nand GNAME4904(G4904,G20203,G2906);
  nand GNAME4905(G4905,G20967,G2907);
  nand GNAME4906(G4906,G59331,G2908);
  nand GNAME4907(G4907,G2909,G59140);
  nand GNAME4908(G4908,G2893,G21471);
  nand GNAME4909(G4909,G20546,G2904);
  nand GNAME4910(G4910,G20204,G2906);
  nand GNAME4911(G4911,G20968,G2907);
  nand GNAME4912(G4912,G59330,G2908);
  nand GNAME4913(G4913,G2909,G59139);
  nand GNAME4914(G4914,G2893,G21472);
  nand GNAME4915(G4915,G20549,G2904);
  nand GNAME4916(G4916,G20205,G2906);
  nand GNAME4917(G4917,G20969,G2907);
  nand GNAME4918(G4918,G59329,G2908);
  nand GNAME4919(G4919,G2909,G59138);
  nand GNAME4920(G4920,G2893,G21474);
  nand GNAME4921(G4921,G20555,G2904);
  nand GNAME4922(G4922,G20206,G2906);
  nand GNAME4923(G4923,G20973,G2907);
  nand GNAME4924(G4924,G59328,G2908);
  nand GNAME4925(G4925,G2909,G59137);
  nand GNAME4926(G4926,G2893,G21475);
  nand GNAME4927(G4927,G20558,G2904);
  nand GNAME4928(G4928,G20207,G2906);
  nand GNAME4929(G4929,G20974,G2907);
  nand GNAME4930(G4930,G59327,G2908);
  nand GNAME4931(G4931,G2909,G59136);
  nand GNAME4932(G4932,G2893,G21476);
  nand GNAME4933(G4933,G20561,G2904);
  nand GNAME4934(G4934,G20208,G2906);
  nand GNAME4935(G4935,G20975,G2907);
  nand GNAME4936(G4936,G59326,G2908);
  nand GNAME4937(G4937,G2909,G59135);
  nand GNAME4938(G4938,G2893,G21446);
  nand GNAME4939(G4939,G20500,G2904);
  nand GNAME4940(G4940,G20236,G2906);
  nand GNAME4941(G4941,G20976,G2907);
  nand GNAME4942(G4942,G59325,G2908);
  nand GNAME4943(G4943,G2909,G59134);
  nand GNAME4944(G4944,G2893,G21447);
  nand GNAME4945(G4945,G20501,G2904);
  nand GNAME4946(G4946,G20239,G2906);
  nand GNAME4947(G4947,G20977,G2907);
  nand GNAME4948(G4948,G59324,G2908);
  nand GNAME4949(G4949,G2909,G59133);
  nand GNAME4950(G4950,G2893,G21448);
  nand GNAME4951(G4951,G20445,G2904);
  nand GNAME4952(G4952,G20211,G2906);
  nand GNAME4953(G4953,G20923,G2907);
  nand GNAME4954(G4954,G59323,G2908);
  nand GNAME4955(G4955,G2909,G59132);
  nand GNAME4956(G4956,G2893,G21449);
  nand GNAME4957(G4957,G20502,G2904);
  nand GNAME4958(G4958,G20243,G2906);
  nand GNAME4959(G4959,G20978,G2907);
  nand GNAME4960(G4960,G59322,G2908);
  nand GNAME4961(G4961,G2909,G59131);
  nand GNAME4962(G4962,G2893,G21450);
  nand GNAME4963(G4963,G20503,G2904);
  nand GNAME4964(G4964,G20246,G2906);
  nand GNAME4965(G4965,G20979,G2907);
  nand GNAME4966(G4966,G59321,G2908);
  nand GNAME4967(G4967,G2909,G59130);
  nand GNAME4968(G4968,G2893,G21451);
  nand GNAME4969(G4969,G20504,G2904);
  nand GNAME4970(G4970,G20212,G2906);
  nand GNAME4971(G4971,G20859,G2907);
  nand GNAME4972(G4972,G59320,G2908);
  nand GNAME4973(G4973,G2909,G59129);
  nand GNAME4974(G4974,G2893,G21452);
  nand GNAME4975(G4975,G20444,G2904);
  nand GNAME4976(G4976,G20140,G2906);
  nand GNAME4977(G4977,G20858,G2907);
  nand GNAME4978(G4978,G59319,G2908);
  nand GNAME4979(G4979,G2909,G59128);
  nand GNAME4980(G4980,G2893,G21434);
  nand GNAME4981(G4981,G20481,G2904);
  nand GNAME4982(G4982,G20219,G2906);
  nand GNAME4983(G4983,G20950,G2907);
  nand GNAME4984(G4984,G59318,G2908);
  nand GNAME4985(G4985,G2909,G59127);
  nand GNAME4986(G4986,G2893,G21435);
  nand GNAME4987(G4987,G20516,G2904);
  nand GNAME4988(G4988,G20176,G2906);
  nand GNAME4989(G4989,G20951,G2907);
  nand GNAME4990(G4990,G59317,G2908);
  nand GNAME4991(G4991,G2909,G59126);
  nand GNAME4992(G4992,G2893,G21436);
  nand GNAME4993(G4993,G20506,G2904);
  nand GNAME4994(G4994,G20177,G2906);
  nand GNAME4995(G4995,G20919,G2907);
  nand GNAME4996(G4996,G59316,G2908);
  nand GNAME4997(G4997,G2909,G59125);
  nand GNAME4998(G4998,G2893,G21437);
  nand GNAME4999(G4999,G20448,G2904);
  nand GNAME5000(G5000,G20143,G2906);
  nand GNAME5001(G5001,G20861,G2907);
  nand GNAME5002(G5002,G59315,G2908);
  nand GNAME5003(G5003,G2909,G59124);
  nand GNAME5004(G5004,G2893,G21438);
  nand GNAME5005(G5005,G20520,G2904);
  nand GNAME5006(G5006,G20178,G2906);
  nand GNAME5007(G5007,G20955,G2907);
  nand GNAME5008(G5008,G59314,G2908);
  nand GNAME5009(G5009,G2909,G59123);
  nand GNAME5010(G5010,G2893,G21439);
  nand GNAME5011(G5011,G20523,G2904);
  nand GNAME5012(G5012,G20179,G2906);
  nand GNAME5013(G5013,G20958,G2907);
  nand GNAME5014(G5014,G59313,G2908);
  nand GNAME5015(G5015,G2909,G59122);
  nand GNAME5016(G5016,G2893,G21440);
  nand GNAME5017(G5017,G20920,G2907);
  nand GNAME5018(G5018,G59312,G2908);
  nand GNAME5019(G5019,G20180,G2906);
  nand GNAME5020(G5020,G20507,G2904);
  nand GNAME5021(G5021,G2909,G59121);
  nand GNAME5022(G5022,G2893,G21443);
  nand GNAME5023(G5023,G20860,G2907);
  nand GNAME5024(G5024,G59311,G2908);
  nand GNAME5025(G5025,G20141,G2906);
  nand GNAME5026(G5026,G20446,G2904);
  nand GNAME5027(G5027,G2909,G59120);
  nand GNAME5028(G5028,G2893,G21445);
  nand GNAME5029(G5029,G20972,G2907);
  nand GNAME5030(G5030,G20552,G2904);
  nand GNAME5031(G5031,G59310,G2908);
  nand GNAME5032(G5032,G20233,G2906);
  nand GNAME5033(G5033,G2909,G59119);
  nand GNAME5034(G5034,G2893,G21453);
  nand GNAME5035(G5035,G20918,G2907);
  nand GNAME5036(G5036,G59309,G2908);
  nand GNAME5037(G5037,G20505,G2904);
  nand GNAME5038(G5038,G20209,G2906);
  nand GNAME5039(G5039,G2909,G59118);
  or GNAME5040(G5040,G2804,G2912);
  not GNAME5041(G5041,G2913);
  or GNAME5042(G5042,G20108,G7987);
  not GNAME5043(G5043,G2920);
  nand GNAME5044(G5044,G59112,G2798);
  nor GNAME5045(G5045,G2788,G58978);
  nand GNAME5046(G5046,G2915,G2916);
  not GNAME5047(G5047,G2917);
  nand GNAME5048(G5048,G2754,G3799);
  nand GNAME5049(G5049,G5048,G3802);
  nand GNAME5050(G5050,G5047,G2918);
  nand GNAME5051(G5051,G20209,G2919);
  nand GNAME5052(G5052,G2910,G7870,G7871);
  nand GNAME5053(G5053,G2748,G2798);
  not GNAME5054(G5054,G2923);
  nand GNAME5055(G5055,G2754,G2955);
  nand GNAME5056(G5056,G59111,G2798);
  nand GNAME5057(G5057,G2816,G59116);
  not GNAME5058(G5058,G2924);
  nand GNAME5059(G5059,G3253,G2918);
  nand GNAME5060(G5060,G20233,G2919);
  nand GNAME5061(G5061,G5043,G59116);
  nand GNAME5062(G5062,G2754,G3254);
  nand GNAME5063(G5063,G59110,G2798);
  nand GNAME5064(G5064,G2816,G59115);
  nand GNAME5065(G5065,G2924,G3804);
  nand GNAME5066(G5066,G5065,G5054);
  nand GNAME5067(G5067,G2922,G5058);
  nand GNAME5068(G5068,G2928,G2927);
  not GNAME5069(G5069,G2929);
  nand GNAME5070(G5070,G2918,G5069);
  nand GNAME5071(G5071,G20141,G2919);
  nand GNAME5072(G5072,G5043,G59115);
  nor GNAME5073(G5073,G2926,G2931);
  nand GNAME5074(G5074,G2754,G2956);
  nand GNAME5075(G5075,G59109,G2798);
  nand GNAME5076(G5076,G2816,G59114);
  nand GNAME5077(G5077,G2918,G7882);
  nand GNAME5078(G5078,G20180,G2919);
  nand GNAME5079(G5079,G5043,G59114);
  nand GNAME5080(G5080,G4473,G2802);
  nand GNAME5081(G5081,G5080,G3980);
  nand GNAME5082(G5082,G5081,G4324);
  nand GNAME5083(G5083,G5082,G20108);
  nand GNAME5084(G5084,G2789,G20773);
  nand GNAME5085(G5085,G5083,G5084);
  nand GNAME5086(G5086,G2752,G5085);
  or GNAME5087(G5087,G3108,G2804);
  nand GNAME5088(G5088,G3781,G2803);
  nand GNAME5089(G5089,G3979,G2897);
  nand GNAME5090(G5090,G5089,G7458);
  nand GNAME5091(G5091,G2795,G58977);
  nand GNAME5092(G5092,G5091,G3778,G3805);
  not GNAME5093(G5093,G2933);
  nand GNAME5094(G5094,G2795,G5093);
  nand GNAME5095(G5095,G5094,G58977);
  nand GNAME5096(G5096,G2917,G2933);
  not GNAME5097(G5097,G2936);
  nand GNAME5098(G5098,G3869,G2933,G58977);
  not GNAME5099(G5099,G2934);
  nand GNAME5100(G5100,G2800,G2894);
  nand GNAME5101(G5101,G5100,G2753);
  nand GNAME5102(G5102,G2786,G5101);
  nand GNAME5103(G5103,G3869,G2899);
  nand GNAME5104(G5104,G2864,G4324,G5102,G5103);
  nand GNAME5105(G5105,G2799,G2824);
  nand GNAME5106(G5106,G5105,G2903);
  nand GNAME5107(G5107,G3955,G2901);
  nand GNAME5108(G5108,G2858,G4473);
  or GNAME5109(G5109,G59112,G3108);
  nand GNAME5110(G5110,G5108,G5099);
  nand GNAME5111(G5111,G5107,G5047);
  nand GNAME5112(G5112,G5106,G20209);
  nand GNAME5113(G5113,G5104,G20505);
  nand GNAME5114(G5114,G5112,G5113,G5111,G5109,G5110);
  nand GNAME5115(G5115,G2917,G7867);
  nand GNAME5116(G5116,G20505,G2932);
  nand GNAME5117(G5117,G5115,G58978);
  nand GNAME5118(G5118,G5114,G2793);
  nand GNAME5119(G5119,G5118,G5116,G5117);
  nand GNAME5120(G5120,G5092,G59111);
  nand GNAME5121(G5121,G2754,G3253);
  not GNAME5122(G5122,G2937);
  not GNAME5123(G5123,G3190);
  nand GNAME5124(G5124,G59112,G3869);
  not GNAME5125(G5125,G3164);
  or GNAME5126(G5126,G2757,G5125);
  nand GNAME5127(G5127,G5126,G2828);
  nand GNAME5128(G5128,G5108,G7889);
  nand GNAME5129(G5129,G5107,G3253);
  nand GNAME5130(G5130,G5106,G20233);
  nand GNAME5131(G5131,G5104,G20552);
  nand GNAME5132(G5132,G3190,G2831);
  nand GNAME5133(G5133,G3404,G5129,G5131,G5128);
  nand GNAME5134(G5134,G3253,G2935);
  nand GNAME5135(G5135,G20552,G2932);
  nand GNAME5136(G5136,G5133,G2793);
  nand GNAME5137(G5137,G5136,G5134,G5135);
  nand GNAME5138(G5138,G2937,G5097);
  nand GNAME5139(G5139,G3778,G5138);
  nand GNAME5140(G5140,G2936,G5122);
  not GNAME5141(G5141,G2939);
  nand GNAME5142(G5142,G5092,G59110);
  nand GNAME5143(G5143,G2754,G5069);
  not GNAME5144(G5144,G2938);
  nand GNAME5145(G5145,G3790,G3258);
  not GNAME5146(G5146,G2940);
  not GNAME5147(G5147,G3779);
  nand GNAME5148(G5148,G5108,G7895);
  nand GNAME5149(G5149,G5107,G5069);
  nand GNAME5150(G5150,G5106,G20141);
  nand GNAME5151(G5151,G5104,G20446);
  nand GNAME5152(G5152,G2828,G7901);
  nand GNAME5153(G5153,G2831,G5146);
  nand GNAME5154(G5154,G3405,G5150,G5148,G5151);
  nand GNAME5155(G5155,G5069,G2935);
  nand GNAME5156(G5156,G20446,G2932);
  nand GNAME5157(G5157,G5154,G2793);
  nand GNAME5158(G5158,G5157,G5155,G5156);
  nand GNAME5159(G5159,G5092,G59109);
  nand GNAME5160(G5160,G5159,G5165);
  nand GNAME5161(G5161,G5166,G5141);
  nand GNAME5162(G5162,G5163,G5160,G5161);
  nand GNAME5163(G5163,G2938,G2823);
  nand GNAME5164(G5164,G2939,G5163);
  nand GNAME5165(G5165,G2754,G7882);
  nand GNAME5166(G5166,G3805,G5144);
  nand GNAME5167(G5167,G5159,G5164,G5165,G5166);
  not GNAME5168(G5168,G2944);
  nand GNAME5169(G5169,G5147,G2756);
  nand GNAME5170(G5170,G2764,G5147);
  nand GNAME5171(G5171,G5170,G59109);
  and GNAME5172(G5172,G2771,G3869);
  or GNAME5173(G5173,G5172,G2756);
  nand GNAME5174(G5174,G2795,G2777);
  not GNAME5175(G5175,G2941);
  nand GNAME5176(G5176,G5108,G2944);
  nand GNAME5177(G5177,G5107,G7882);
  nand GNAME5178(G5178,G5106,G20180);
  nand GNAME5179(G5179,G5104,G20507);
  nand GNAME5180(G5180,G2831,G5175);
  nand GNAME5181(G5181,G2828,G3809);
  nand GNAME5182(G5182,G3406,G5178,G5176,G5179);
  nand GNAME5183(G5183,G20507,G2932);
  nand GNAME5184(G5184,G5182,G2793);
  nand GNAME5185(G5185,G5183,G5184);
  nand GNAME5186(G5186,G2795,G2965);
  nand GNAME5187(G5187,G58977,G2962);
  nand GNAME5188(G5188,G5186,G5187);
  not GNAME5189(G5189,G2950);
  nand GNAME5190(G5190,G2836,G2959);
  nand GNAME5191(G5191,G58977,G5189);
  nand GNAME5192(G5192,G5190,G5191);
  nand GNAME5193(G5193,G2950,G2951);
  and GNAME5194(G5194,G5193,G3803);
  nand GNAME5195(G5195,G2959,G2950,G2951);
  nand GNAME5196(G5196,G2960,G2961);
  nand GNAME5197(G5197,G5195,G5196);
  and GNAME5198(G5198,G2950,G58977);
  nor GNAME5199(G5199,G5198,G2805,G2961);
  or GNAME5200(G5200,G2960,G5199);
  nand GNAME5201(G5201,G5200,G2913);
  nand GNAME5202(G5202,G58887,G2952);
  nand GNAME5203(G5203,G5201,G59107);
  nand GNAME5204(G5204,G5197,G58871);
  nand GNAME5205(G5205,G5192,G2962);
  nand GNAME5206(G5206,G2963,G2964);
  nand GNAME5207(G5207,G5188,G2960);
  nand GNAME5208(G5208,G2799,G2965);
  nand GNAME5209(G5209,G58977,G2966);
  nand GNAME5210(G5210,G5208,G5209);
  nand GNAME5211(G5211,G58888,G2952);
  nand GNAME5212(G5212,G5201,G59106);
  nand GNAME5213(G5213,G5197,G58872);
  nand GNAME5214(G5214,G5192,G2966);
  nand GNAME5215(G5215,G2963,G2967);
  nand GNAME5216(G5216,G5210,G2960);
  nand GNAME5217(G5217,G2784,G2965);
  nand GNAME5218(G5218,G58977,G2968);
  nand GNAME5219(G5219,G5217,G5218);
  nand GNAME5220(G5220,G58889,G2952);
  nand GNAME5221(G5221,G5201,G59105);
  nand GNAME5222(G5222,G5197,G58873);
  nand GNAME5223(G5223,G5192,G2968);
  nand GNAME5224(G5224,G2963,G2969);
  nand GNAME5225(G5225,G5219,G2960);
  nand GNAME5226(G5226,G2749,G2965);
  nand GNAME5227(G5227,G58977,G2970);
  nand GNAME5228(G5228,G5226,G5227);
  nand GNAME5229(G5229,G58890,G2952);
  nand GNAME5230(G5230,G5201,G59104);
  nand GNAME5231(G5231,G5197,G58874);
  nand GNAME5232(G5232,G5192,G2970);
  nand GNAME5233(G5233,G2963,G2971);
  nand GNAME5234(G5234,G5228,G2960);
  nand GNAME5235(G5235,G2786,G2965);
  nand GNAME5236(G5236,G58977,G2972);
  nand GNAME5237(G5237,G5235,G5236);
  nand GNAME5238(G5238,G58891,G2952);
  nand GNAME5239(G5239,G5201,G59103);
  nand GNAME5240(G5240,G5197,G58875);
  nand GNAME5241(G5241,G5192,G2972);
  nand GNAME5242(G5242,G2963,G2973);
  nand GNAME5243(G5243,G5237,G2960);
  nand GNAME5244(G5244,G2783,G2965);
  nand GNAME5245(G5245,G58977,G2974);
  nand GNAME5246(G5246,G5244,G5245);
  nand GNAME5247(G5247,G58892,G2952);
  nand GNAME5248(G5248,G5201,G59102);
  nand GNAME5249(G5249,G5197,G58876);
  nand GNAME5250(G5250,G5192,G2974);
  nand GNAME5251(G5251,G2963,G2975);
  nand GNAME5252(G5252,G5246,G2960);
  nand GNAME5253(G5253,G2785,G2965);
  nand GNAME5254(G5254,G58977,G2976);
  nand GNAME5255(G5255,G5253,G5254);
  nand GNAME5256(G5256,G58893,G2952);
  nand GNAME5257(G5257,G5201,G59101);
  nand GNAME5258(G5258,G5197,G58877);
  nand GNAME5259(G5259,G5192,G2976);
  nand GNAME5260(G5260,G2963,G2977);
  nand GNAME5261(G5261,G5255,G2960);
  nand GNAME5262(G5262,G2855,G2965);
  nand GNAME5263(G5263,G58977,G2978);
  nand GNAME5264(G5264,G5262,G5263);
  nand GNAME5265(G5265,G58894,G2952);
  nand GNAME5266(G5266,G5201,G59100);
  nand GNAME5267(G5267,G5197,G58878);
  nand GNAME5268(G5268,G5192,G2978);
  nand GNAME5269(G5269,G2963,G2979);
  nand GNAME5270(G5270,G5264,G2960);
  not GNAME5271(G5271,G2982);
  nand GNAME5272(G5272,G2836,G2987);
  nand GNAME5273(G5273,G58977,G5271);
  nand GNAME5274(G5274,G5272,G5273);
  nand GNAME5275(G5275,G2982,G2983);
  and GNAME5276(G5276,G5275,G3803);
  nand GNAME5277(G5277,G2987,G2982,G2983);
  nand GNAME5278(G5278,G2988,G2989);
  nand GNAME5279(G5279,G5277,G5278);
  and GNAME5280(G5280,G2982,G58977);
  nor GNAME5281(G5281,G5280,G2805,G2989);
  or GNAME5282(G5282,G2988,G5281);
  nand GNAME5283(G5283,G5282,G2913);
  nand GNAME5284(G5284,G58887,G2984);
  nand GNAME5285(G5285,G5283,G59099);
  nand GNAME5286(G5286,G5279,G58871);
  nand GNAME5287(G5287,G5274,G2962);
  nand GNAME5288(G5288,G2964,G2990);
  nand GNAME5289(G5289,G5188,G2988);
  nand GNAME5290(G5290,G58888,G2984);
  nand GNAME5291(G5291,G5283,G59098);
  nand GNAME5292(G5292,G5279,G58872);
  nand GNAME5293(G5293,G5274,G2966);
  nand GNAME5294(G5294,G2967,G2990);
  nand GNAME5295(G5295,G5210,G2988);
  nand GNAME5296(G5296,G58889,G2984);
  nand GNAME5297(G5297,G5283,G59097);
  nand GNAME5298(G5298,G5279,G58873);
  nand GNAME5299(G5299,G5274,G2968);
  nand GNAME5300(G5300,G2969,G2990);
  nand GNAME5301(G5301,G5219,G2988);
  nand GNAME5302(G5302,G58890,G2984);
  nand GNAME5303(G5303,G5283,G59096);
  nand GNAME5304(G5304,G5279,G58874);
  nand GNAME5305(G5305,G5274,G2970);
  nand GNAME5306(G5306,G2971,G2990);
  nand GNAME5307(G5307,G5228,G2988);
  nand GNAME5308(G5308,G58891,G2984);
  nand GNAME5309(G5309,G5283,G59095);
  nand GNAME5310(G5310,G5279,G58875);
  nand GNAME5311(G5311,G5274,G2972);
  nand GNAME5312(G5312,G2973,G2990);
  nand GNAME5313(G5313,G5237,G2988);
  nand GNAME5314(G5314,G58892,G2984);
  nand GNAME5315(G5315,G5283,G59094);
  nand GNAME5316(G5316,G5279,G58876);
  nand GNAME5317(G5317,G5274,G2974);
  nand GNAME5318(G5318,G2975,G2990);
  nand GNAME5319(G5319,G5246,G2988);
  nand GNAME5320(G5320,G58893,G2984);
  nand GNAME5321(G5321,G5283,G59093);
  nand GNAME5322(G5322,G5279,G58877);
  nand GNAME5323(G5323,G5274,G2976);
  nand GNAME5324(G5324,G2977,G2990);
  nand GNAME5325(G5325,G5255,G2988);
  nand GNAME5326(G5326,G58894,G2984);
  nand GNAME5327(G5327,G5283,G59092);
  nand GNAME5328(G5328,G5279,G58878);
  nand GNAME5329(G5329,G5274,G2978);
  nand GNAME5330(G5330,G2979,G2990);
  nand GNAME5331(G5331,G5264,G2988);
  not GNAME5332(G5332,G2993);
  nand GNAME5333(G5333,G2836,G2998);
  nand GNAME5334(G5334,G58977,G5332);
  nand GNAME5335(G5335,G5333,G5334);
  nand GNAME5336(G5336,G2993,G2994);
  and GNAME5337(G5337,G5336,G3803);
  nand GNAME5338(G5338,G2998,G2993,G2994);
  nand GNAME5339(G5339,G2999,G3000);
  nand GNAME5340(G5340,G5338,G5339);
  and GNAME5341(G5341,G2993,G58977);
  nor GNAME5342(G5342,G5341,G2805,G3000);
  or GNAME5343(G5343,G2999,G5342);
  nand GNAME5344(G5344,G5343,G2913);
  nand GNAME5345(G5345,G58887,G2995);
  nand GNAME5346(G5346,G5344,G59091);
  nand GNAME5347(G5347,G5340,G58871);
  nand GNAME5348(G5348,G5335,G2962);
  nand GNAME5349(G5349,G2964,G3001);
  nand GNAME5350(G5350,G5188,G2999);
  nand GNAME5351(G5351,G58888,G2995);
  nand GNAME5352(G5352,G5344,G59090);
  nand GNAME5353(G5353,G5340,G58872);
  nand GNAME5354(G5354,G5335,G2966);
  nand GNAME5355(G5355,G2967,G3001);
  nand GNAME5356(G5356,G5210,G2999);
  nand GNAME5357(G5357,G58889,G2995);
  nand GNAME5358(G5358,G5344,G59089);
  nand GNAME5359(G5359,G5340,G58873);
  nand GNAME5360(G5360,G5335,G2968);
  nand GNAME5361(G5361,G2969,G3001);
  nand GNAME5362(G5362,G5219,G2999);
  nand GNAME5363(G5363,G58890,G2995);
  nand GNAME5364(G5364,G5344,G59088);
  nand GNAME5365(G5365,G5340,G58874);
  nand GNAME5366(G5366,G5335,G2970);
  nand GNAME5367(G5367,G2971,G3001);
  nand GNAME5368(G5368,G5228,G2999);
  nand GNAME5369(G5369,G58891,G2995);
  nand GNAME5370(G5370,G5344,G59087);
  nand GNAME5371(G5371,G5340,G58875);
  nand GNAME5372(G5372,G5335,G2972);
  nand GNAME5373(G5373,G2973,G3001);
  nand GNAME5374(G5374,G5237,G2999);
  nand GNAME5375(G5375,G58892,G2995);
  nand GNAME5376(G5376,G5344,G59086);
  nand GNAME5377(G5377,G5340,G58876);
  nand GNAME5378(G5378,G5335,G2974);
  nand GNAME5379(G5379,G2975,G3001);
  nand GNAME5380(G5380,G5246,G2999);
  nand GNAME5381(G5381,G58893,G2995);
  nand GNAME5382(G5382,G5344,G59085);
  nand GNAME5383(G5383,G5340,G58877);
  nand GNAME5384(G5384,G5335,G2976);
  nand GNAME5385(G5385,G2977,G3001);
  nand GNAME5386(G5386,G5255,G2999);
  nand GNAME5387(G5387,G58894,G2995);
  nand GNAME5388(G5388,G5344,G59084);
  nand GNAME5389(G5389,G5340,G58878);
  nand GNAME5390(G5390,G5335,G2978);
  nand GNAME5391(G5391,G2979,G3001);
  nand GNAME5392(G5392,G5264,G2999);
  not GNAME5393(G5393,G3002);
  nand GNAME5394(G5394,G2836,G3006);
  nand GNAME5395(G5395,G58977,G5393);
  nand GNAME5396(G5396,G5394,G5395);
  nand GNAME5397(G5397,G3002,G3003);
  and GNAME5398(G5398,G5397,G3803);
  nand GNAME5399(G5399,G3003,G3006);
  nand GNAME5400(G5400,G3007,G3008);
  nand GNAME5401(G5401,G5399,G5400);
  and GNAME5402(G5402,G3002,G58977);
  nor GNAME5403(G5403,G5402,G2805,G3008);
  or GNAME5404(G5404,G3007,G5403);
  nand GNAME5405(G5405,G5404,G2913);
  nand GNAME5406(G5406,G58887,G3004);
  nand GNAME5407(G5407,G5405,G59083);
  nand GNAME5408(G5408,G5401,G58871);
  nand GNAME5409(G5409,G5396,G2962);
  nand GNAME5410(G5410,G2964,G3009);
  nand GNAME5411(G5411,G5188,G3007);
  nand GNAME5412(G5412,G58888,G3004);
  nand GNAME5413(G5413,G5405,G59082);
  nand GNAME5414(G5414,G5401,G58872);
  nand GNAME5415(G5415,G5396,G2966);
  nand GNAME5416(G5416,G2967,G3009);
  nand GNAME5417(G5417,G5210,G3007);
  nand GNAME5418(G5418,G58889,G3004);
  nand GNAME5419(G5419,G5405,G59081);
  nand GNAME5420(G5420,G5401,G58873);
  nand GNAME5421(G5421,G5396,G2968);
  nand GNAME5422(G5422,G2969,G3009);
  nand GNAME5423(G5423,G5219,G3007);
  nand GNAME5424(G5424,G58890,G3004);
  nand GNAME5425(G5425,G5405,G59080);
  nand GNAME5426(G5426,G5401,G58874);
  nand GNAME5427(G5427,G5396,G2970);
  nand GNAME5428(G5428,G2971,G3009);
  nand GNAME5429(G5429,G5228,G3007);
  nand GNAME5430(G5430,G58891,G3004);
  nand GNAME5431(G5431,G5405,G59079);
  nand GNAME5432(G5432,G5401,G58875);
  nand GNAME5433(G5433,G5396,G2972);
  nand GNAME5434(G5434,G2973,G3009);
  nand GNAME5435(G5435,G5237,G3007);
  nand GNAME5436(G5436,G58892,G3004);
  nand GNAME5437(G5437,G5405,G59078);
  nand GNAME5438(G5438,G5401,G58876);
  nand GNAME5439(G5439,G5396,G2974);
  nand GNAME5440(G5440,G2975,G3009);
  nand GNAME5441(G5441,G5246,G3007);
  nand GNAME5442(G5442,G58893,G3004);
  nand GNAME5443(G5443,G5405,G59077);
  nand GNAME5444(G5444,G5401,G58877);
  nand GNAME5445(G5445,G5396,G2976);
  nand GNAME5446(G5446,G2977,G3009);
  nand GNAME5447(G5447,G5255,G3007);
  nand GNAME5448(G5448,G58894,G3004);
  nand GNAME5449(G5449,G5405,G59076);
  nand GNAME5450(G5450,G5401,G58878);
  nand GNAME5451(G5451,G5396,G2978);
  nand GNAME5452(G5452,G2979,G3009);
  nand GNAME5453(G5453,G5264,G3007);
  not GNAME5454(G5454,G3012);
  nand GNAME5455(G5455,G2836,G3016);
  nand GNAME5456(G5456,G58977,G5454);
  nand GNAME5457(G5457,G5455,G5456);
  nand GNAME5458(G5458,G3012,G3013);
  and GNAME5459(G5459,G5458,G3803);
  nand GNAME5460(G5460,G3016,G3012,G3013);
  nand GNAME5461(G5461,G3017,G3018);
  nand GNAME5462(G5462,G5460,G5461);
  and GNAME5463(G5463,G3012,G58977);
  nor GNAME5464(G5464,G5463,G2805,G3018);
  or GNAME5465(G5465,G3017,G5464);
  nand GNAME5466(G5466,G5465,G2913);
  nand GNAME5467(G5467,G58887,G3014);
  nand GNAME5468(G5468,G5466,G59075);
  nand GNAME5469(G5469,G5462,G58871);
  nand GNAME5470(G5470,G5457,G2962);
  nand GNAME5471(G5471,G2964,G3019);
  nand GNAME5472(G5472,G5188,G3017);
  nand GNAME5473(G5473,G58888,G3014);
  nand GNAME5474(G5474,G5466,G59074);
  nand GNAME5475(G5475,G5462,G58872);
  nand GNAME5476(G5476,G5457,G2966);
  nand GNAME5477(G5477,G2967,G3019);
  nand GNAME5478(G5478,G5210,G3017);
  nand GNAME5479(G5479,G58889,G3014);
  nand GNAME5480(G5480,G5466,G59073);
  nand GNAME5481(G5481,G5462,G58873);
  nand GNAME5482(G5482,G5457,G2968);
  nand GNAME5483(G5483,G2969,G3019);
  nand GNAME5484(G5484,G5219,G3017);
  nand GNAME5485(G5485,G58890,G3014);
  nand GNAME5486(G5486,G5466,G59072);
  nand GNAME5487(G5487,G5462,G58874);
  nand GNAME5488(G5488,G5457,G2970);
  nand GNAME5489(G5489,G2971,G3019);
  nand GNAME5490(G5490,G5228,G3017);
  nand GNAME5491(G5491,G58891,G3014);
  nand GNAME5492(G5492,G5466,G59071);
  nand GNAME5493(G5493,G5462,G58875);
  nand GNAME5494(G5494,G5457,G2972);
  nand GNAME5495(G5495,G2973,G3019);
  nand GNAME5496(G5496,G5237,G3017);
  nand GNAME5497(G5497,G58892,G3014);
  nand GNAME5498(G5498,G5466,G59070);
  nand GNAME5499(G5499,G5462,G58876);
  nand GNAME5500(G5500,G5457,G2974);
  nand GNAME5501(G5501,G2975,G3019);
  nand GNAME5502(G5502,G5246,G3017);
  nand GNAME5503(G5503,G58893,G3014);
  nand GNAME5504(G5504,G5466,G59069);
  nand GNAME5505(G5505,G5462,G58877);
  nand GNAME5506(G5506,G5457,G2976);
  nand GNAME5507(G5507,G2977,G3019);
  nand GNAME5508(G5508,G5255,G3017);
  nand GNAME5509(G5509,G58894,G3014);
  nand GNAME5510(G5510,G5466,G59068);
  nand GNAME5511(G5511,G5462,G58878);
  nand GNAME5512(G5512,G5457,G2978);
  nand GNAME5513(G5513,G2979,G3019);
  nand GNAME5514(G5514,G5264,G3017);
  not GNAME5515(G5515,G3022);
  nand GNAME5516(G5516,G2836,G3025);
  nand GNAME5517(G5517,G58977,G5515);
  nand GNAME5518(G5518,G5516,G5517);
  nand GNAME5519(G5519,G3022,G3023);
  and GNAME5520(G5520,G5519,G3803);
  nand GNAME5521(G5521,G3023,G3025);
  nand GNAME5522(G5522,G3026,G3027);
  nand GNAME5523(G5523,G5521,G5522);
  and GNAME5524(G5524,G3022,G58977);
  nor GNAME5525(G5525,G5524,G2805,G3027);
  or GNAME5526(G5526,G3026,G5525);
  nand GNAME5527(G5527,G5526,G2913);
  nand GNAME5528(G5528,G58887,G3024);
  nand GNAME5529(G5529,G5527,G59067);
  nand GNAME5530(G5530,G5523,G58871);
  nand GNAME5531(G5531,G5518,G2962);
  nand GNAME5532(G5532,G2964,G3028);
  nand GNAME5533(G5533,G5188,G3026);
  nand GNAME5534(G5534,G58888,G3024);
  nand GNAME5535(G5535,G5527,G59066);
  nand GNAME5536(G5536,G5523,G58872);
  nand GNAME5537(G5537,G5518,G2966);
  nand GNAME5538(G5538,G2967,G3028);
  nand GNAME5539(G5539,G5210,G3026);
  nand GNAME5540(G5540,G58889,G3024);
  nand GNAME5541(G5541,G5527,G59065);
  nand GNAME5542(G5542,G5523,G58873);
  nand GNAME5543(G5543,G5518,G2968);
  nand GNAME5544(G5544,G2969,G3028);
  nand GNAME5545(G5545,G5219,G3026);
  nand GNAME5546(G5546,G58890,G3024);
  nand GNAME5547(G5547,G5527,G59064);
  nand GNAME5548(G5548,G5523,G58874);
  nand GNAME5549(G5549,G5518,G2970);
  nand GNAME5550(G5550,G2971,G3028);
  nand GNAME5551(G5551,G5228,G3026);
  nand GNAME5552(G5552,G58891,G3024);
  nand GNAME5553(G5553,G5527,G59063);
  nand GNAME5554(G5554,G5523,G58875);
  nand GNAME5555(G5555,G5518,G2972);
  nand GNAME5556(G5556,G2973,G3028);
  nand GNAME5557(G5557,G5237,G3026);
  nand GNAME5558(G5558,G58892,G3024);
  nand GNAME5559(G5559,G5527,G59062);
  nand GNAME5560(G5560,G5523,G58876);
  nand GNAME5561(G5561,G5518,G2974);
  nand GNAME5562(G5562,G2975,G3028);
  nand GNAME5563(G5563,G5246,G3026);
  nand GNAME5564(G5564,G58893,G3024);
  nand GNAME5565(G5565,G5527,G59061);
  nand GNAME5566(G5566,G5523,G58877);
  nand GNAME5567(G5567,G5518,G2976);
  nand GNAME5568(G5568,G2977,G3028);
  nand GNAME5569(G5569,G5255,G3026);
  nand GNAME5570(G5570,G58894,G3024);
  nand GNAME5571(G5571,G5527,G59060);
  nand GNAME5572(G5572,G5523,G58878);
  nand GNAME5573(G5573,G5518,G2978);
  nand GNAME5574(G5574,G2979,G3028);
  nand GNAME5575(G5575,G5264,G3026);
  not GNAME5576(G5576,G3029);
  nand GNAME5577(G5577,G2836,G3032);
  nand GNAME5578(G5578,G58977,G5576);
  nand GNAME5579(G5579,G5577,G5578);
  nand GNAME5580(G5580,G3029,G3030);
  and GNAME5581(G5581,G5580,G3803);
  nand GNAME5582(G5582,G3032,G3029,G3030);
  nand GNAME5583(G5583,G3033,G3034);
  nand GNAME5584(G5584,G5582,G5583);
  and GNAME5585(G5585,G3029,G58977);
  nor GNAME5586(G5586,G5585,G2805,G3034);
  or GNAME5587(G5587,G3033,G5586);
  nand GNAME5588(G5588,G5587,G2913);
  nand GNAME5589(G5589,G58887,G3031);
  nand GNAME5590(G5590,G5588,G59059);
  nand GNAME5591(G5591,G5584,G58871);
  nand GNAME5592(G5592,G5579,G2962);
  nand GNAME5593(G5593,G2964,G3035);
  nand GNAME5594(G5594,G5188,G3033);
  nand GNAME5595(G5595,G58888,G3031);
  nand GNAME5596(G5596,G5588,G59058);
  nand GNAME5597(G5597,G5584,G58872);
  nand GNAME5598(G5598,G5579,G2966);
  nand GNAME5599(G5599,G2967,G3035);
  nand GNAME5600(G5600,G5210,G3033);
  nand GNAME5601(G5601,G58889,G3031);
  nand GNAME5602(G5602,G5588,G59057);
  nand GNAME5603(G5603,G5584,G58873);
  nand GNAME5604(G5604,G5579,G2968);
  nand GNAME5605(G5605,G2969,G3035);
  nand GNAME5606(G5606,G5219,G3033);
  nand GNAME5607(G5607,G58890,G3031);
  nand GNAME5608(G5608,G5588,G59056);
  nand GNAME5609(G5609,G5584,G58874);
  nand GNAME5610(G5610,G5579,G2970);
  nand GNAME5611(G5611,G2971,G3035);
  nand GNAME5612(G5612,G5228,G3033);
  nand GNAME5613(G5613,G58891,G3031);
  nand GNAME5614(G5614,G5588,G59055);
  nand GNAME5615(G5615,G5584,G58875);
  nand GNAME5616(G5616,G5579,G2972);
  nand GNAME5617(G5617,G2973,G3035);
  nand GNAME5618(G5618,G5237,G3033);
  nand GNAME5619(G5619,G58892,G3031);
  nand GNAME5620(G5620,G5588,G59054);
  nand GNAME5621(G5621,G5584,G58876);
  nand GNAME5622(G5622,G5579,G2974);
  nand GNAME5623(G5623,G2975,G3035);
  nand GNAME5624(G5624,G5246,G3033);
  nand GNAME5625(G5625,G58893,G3031);
  nand GNAME5626(G5626,G5588,G59053);
  nand GNAME5627(G5627,G5584,G58877);
  nand GNAME5628(G5628,G5579,G2976);
  nand GNAME5629(G5629,G2977,G3035);
  nand GNAME5630(G5630,G5255,G3033);
  nand GNAME5631(G5631,G58894,G3031);
  nand GNAME5632(G5632,G5588,G59052);
  nand GNAME5633(G5633,G5584,G58878);
  nand GNAME5634(G5634,G5579,G2978);
  nand GNAME5635(G5635,G2979,G3035);
  nand GNAME5636(G5636,G5264,G3033);
  not GNAME5637(G5637,G3036);
  nand GNAME5638(G5638,G2836,G3039);
  nand GNAME5639(G5639,G58977,G5637);
  nand GNAME5640(G5640,G5638,G5639);
  nand GNAME5641(G5641,G3036,G3037);
  and GNAME5642(G5642,G5641,G3803);
  nand GNAME5643(G5643,G3037,G3039);
  nand GNAME5644(G5644,G3040,G3041);
  nand GNAME5645(G5645,G5643,G5644);
  and GNAME5646(G5646,G3036,G58977);
  nor GNAME5647(G5647,G5646,G2805,G3040);
  or GNAME5648(G5648,G3041,G5647);
  nand GNAME5649(G5649,G5648,G2913);
  nand GNAME5650(G5650,G58887,G3038);
  nand GNAME5651(G5651,G5649,G59051);
  nand GNAME5652(G5652,G5645,G58871);
  nand GNAME5653(G5653,G5640,G2962);
  nand GNAME5654(G5654,G2964,G3042);
  nand GNAME5655(G5655,G5188,G3041);
  nand GNAME5656(G5656,G58888,G3038);
  nand GNAME5657(G5657,G5649,G59050);
  nand GNAME5658(G5658,G5645,G58872);
  nand GNAME5659(G5659,G5640,G2966);
  nand GNAME5660(G5660,G2967,G3042);
  nand GNAME5661(G5661,G5210,G3041);
  nand GNAME5662(G5662,G58889,G3038);
  nand GNAME5663(G5663,G5649,G59049);
  nand GNAME5664(G5664,G5645,G58873);
  nand GNAME5665(G5665,G5640,G2968);
  nand GNAME5666(G5666,G2969,G3042);
  nand GNAME5667(G5667,G5219,G3041);
  nand GNAME5668(G5668,G58890,G3038);
  nand GNAME5669(G5669,G5649,G59048);
  nand GNAME5670(G5670,G5645,G58874);
  nand GNAME5671(G5671,G5640,G2970);
  nand GNAME5672(G5672,G2971,G3042);
  nand GNAME5673(G5673,G5228,G3041);
  nand GNAME5674(G5674,G58891,G3038);
  nand GNAME5675(G5675,G5649,G59047);
  nand GNAME5676(G5676,G5645,G58875);
  nand GNAME5677(G5677,G5640,G2972);
  nand GNAME5678(G5678,G2973,G3042);
  nand GNAME5679(G5679,G5237,G3041);
  nand GNAME5680(G5680,G58892,G3038);
  nand GNAME5681(G5681,G5649,G59046);
  nand GNAME5682(G5682,G5645,G58876);
  nand GNAME5683(G5683,G5640,G2974);
  nand GNAME5684(G5684,G2975,G3042);
  nand GNAME5685(G5685,G5246,G3041);
  nand GNAME5686(G5686,G58893,G3038);
  nand GNAME5687(G5687,G5649,G59045);
  nand GNAME5688(G5688,G5645,G58877);
  nand GNAME5689(G5689,G5640,G2976);
  nand GNAME5690(G5690,G2977,G3042);
  nand GNAME5691(G5691,G5255,G3041);
  nand GNAME5692(G5692,G58894,G3038);
  nand GNAME5693(G5693,G5649,G59044);
  nand GNAME5694(G5694,G5645,G58878);
  nand GNAME5695(G5695,G5640,G2978);
  nand GNAME5696(G5696,G2979,G3042);
  nand GNAME5697(G5697,G5264,G3041);
  not GNAME5698(G5698,G3045);
  nand GNAME5699(G5699,G58977,G5698);
  nand GNAME5700(G5700,G2836,G3050);
  nand GNAME5701(G5701,G5699,G5700);
  nand GNAME5702(G5702,G3045,G3046);
  and GNAME5703(G5703,G5702,G3803);
  nand GNAME5704(G5704,G3050,G3045,G3046);
  nand GNAME5705(G5705,G3051,G3052);
  nand GNAME5706(G5706,G5704,G5705);
  and GNAME5707(G5707,G3045,G58977);
  nor GNAME5708(G5708,G5707,G2805,G3052);
  or GNAME5709(G5709,G3051,G5708);
  nand GNAME5710(G5710,G5709,G2913);
  nand GNAME5711(G5711,G58887,G3047);
  nand GNAME5712(G5712,G5710,G59043);
  nand GNAME5713(G5713,G5706,G58871);
  nand GNAME5714(G5714,G5701,G2962);
  nand GNAME5715(G5715,G2964,G3053);
  nand GNAME5716(G5716,G5188,G3051);
  nand GNAME5717(G5717,G58888,G3047);
  nand GNAME5718(G5718,G5710,G59042);
  nand GNAME5719(G5719,G5706,G58872);
  nand GNAME5720(G5720,G5701,G2966);
  nand GNAME5721(G5721,G2967,G3053);
  nand GNAME5722(G5722,G5210,G3051);
  nand GNAME5723(G5723,G58889,G3047);
  nand GNAME5724(G5724,G5710,G59041);
  nand GNAME5725(G5725,G5706,G58873);
  nand GNAME5726(G5726,G5701,G2968);
  nand GNAME5727(G5727,G2969,G3053);
  nand GNAME5728(G5728,G5219,G3051);
  nand GNAME5729(G5729,G58890,G3047);
  nand GNAME5730(G5730,G5710,G59040);
  nand GNAME5731(G5731,G5706,G58874);
  nand GNAME5732(G5732,G5701,G2970);
  nand GNAME5733(G5733,G2971,G3053);
  nand GNAME5734(G5734,G5228,G3051);
  nand GNAME5735(G5735,G58891,G3047);
  nand GNAME5736(G5736,G5710,G59039);
  nand GNAME5737(G5737,G5706,G58875);
  nand GNAME5738(G5738,G5701,G2972);
  nand GNAME5739(G5739,G2973,G3053);
  nand GNAME5740(G5740,G5237,G3051);
  nand GNAME5741(G5741,G58892,G3047);
  nand GNAME5742(G5742,G5710,G59038);
  nand GNAME5743(G5743,G5706,G58876);
  nand GNAME5744(G5744,G5701,G2974);
  nand GNAME5745(G5745,G2975,G3053);
  nand GNAME5746(G5746,G5246,G3051);
  nand GNAME5747(G5747,G58893,G3047);
  nand GNAME5748(G5748,G5710,G59037);
  nand GNAME5749(G5749,G5706,G58877);
  nand GNAME5750(G5750,G5701,G2976);
  nand GNAME5751(G5751,G2977,G3053);
  nand GNAME5752(G5752,G5255,G3051);
  nand GNAME5753(G5753,G58894,G3047);
  nand GNAME5754(G5754,G5710,G59036);
  nand GNAME5755(G5755,G5706,G58878);
  nand GNAME5756(G5756,G5701,G2978);
  nand GNAME5757(G5757,G2979,G3053);
  nand GNAME5758(G5758,G5264,G3051);
  not GNAME5759(G5759,G3054);
  nand GNAME5760(G5760,G58977,G5759);
  nand GNAME5761(G5761,G2836,G3057);
  nand GNAME5762(G5762,G5760,G5761);
  nand GNAME5763(G5763,G3054,G3055);
  and GNAME5764(G5764,G5763,G3803);
  nand GNAME5765(G5765,G3057,G3054,G3055);
  nand GNAME5766(G5766,G3058,G3059);
  nand GNAME5767(G5767,G5765,G5766);
  and GNAME5768(G5768,G3054,G58977);
  nor GNAME5769(G5769,G5768,G2805,G3059);
  or GNAME5770(G5770,G3058,G5769);
  nand GNAME5771(G5771,G5770,G2913);
  nand GNAME5772(G5772,G58887,G3056);
  nand GNAME5773(G5773,G5771,G59035);
  nand GNAME5774(G5774,G5767,G58871);
  nand GNAME5775(G5775,G5762,G2962);
  nand GNAME5776(G5776,G2964,G3060);
  nand GNAME5777(G5777,G5188,G3058);
  nand GNAME5778(G5778,G58888,G3056);
  nand GNAME5779(G5779,G5771,G59034);
  nand GNAME5780(G5780,G5767,G58872);
  nand GNAME5781(G5781,G5762,G2966);
  nand GNAME5782(G5782,G2967,G3060);
  nand GNAME5783(G5783,G5210,G3058);
  nand GNAME5784(G5784,G58889,G3056);
  nand GNAME5785(G5785,G5771,G59033);
  nand GNAME5786(G5786,G5767,G58873);
  nand GNAME5787(G5787,G5762,G2968);
  nand GNAME5788(G5788,G2969,G3060);
  nand GNAME5789(G5789,G5219,G3058);
  nand GNAME5790(G5790,G58890,G3056);
  nand GNAME5791(G5791,G5771,G59032);
  nand GNAME5792(G5792,G5767,G58874);
  nand GNAME5793(G5793,G5762,G2970);
  nand GNAME5794(G5794,G2971,G3060);
  nand GNAME5795(G5795,G5228,G3058);
  nand GNAME5796(G5796,G58891,G3056);
  nand GNAME5797(G5797,G5771,G59031);
  nand GNAME5798(G5798,G5767,G58875);
  nand GNAME5799(G5799,G5762,G2972);
  nand GNAME5800(G5800,G2973,G3060);
  nand GNAME5801(G5801,G5237,G3058);
  nand GNAME5802(G5802,G58892,G3056);
  nand GNAME5803(G5803,G5771,G59030);
  nand GNAME5804(G5804,G5767,G58876);
  nand GNAME5805(G5805,G5762,G2974);
  nand GNAME5806(G5806,G2975,G3060);
  nand GNAME5807(G5807,G5246,G3058);
  nand GNAME5808(G5808,G58893,G3056);
  nand GNAME5809(G5809,G5771,G59029);
  nand GNAME5810(G5810,G5767,G58877);
  nand GNAME5811(G5811,G5762,G2976);
  nand GNAME5812(G5812,G2977,G3060);
  nand GNAME5813(G5813,G5255,G3058);
  nand GNAME5814(G5814,G58894,G3056);
  nand GNAME5815(G5815,G5771,G59028);
  nand GNAME5816(G5816,G5767,G58878);
  nand GNAME5817(G5817,G5762,G2978);
  nand GNAME5818(G5818,G2979,G3060);
  nand GNAME5819(G5819,G5264,G3058);
  not GNAME5820(G5820,G3063);
  nand GNAME5821(G5821,G58977,G5820);
  nand GNAME5822(G5822,G2836,G3066);
  nand GNAME5823(G5823,G5821,G5822);
  nand GNAME5824(G5824,G3063,G3064);
  and GNAME5825(G5825,G5824,G3803);
  nand GNAME5826(G5826,G3066,G3063,G3064);
  nand GNAME5827(G5827,G3067,G3068);
  nand GNAME5828(G5828,G5826,G5827);
  and GNAME5829(G5829,G3063,G58977);
  nor GNAME5830(G5830,G5829,G2805,G3068);
  or GNAME5831(G5831,G3067,G5830);
  nand GNAME5832(G5832,G5831,G2913);
  nand GNAME5833(G5833,G58887,G3065);
  nand GNAME5834(G5834,G5832,G59027);
  nand GNAME5835(G5835,G5828,G58871);
  nand GNAME5836(G5836,G5823,G2962);
  nand GNAME5837(G5837,G2964,G3069);
  nand GNAME5838(G5838,G5188,G3067);
  nand GNAME5839(G5839,G58888,G3065);
  nand GNAME5840(G5840,G5832,G59026);
  nand GNAME5841(G5841,G5828,G58872);
  nand GNAME5842(G5842,G5823,G2966);
  nand GNAME5843(G5843,G2967,G3069);
  nand GNAME5844(G5844,G5210,G3067);
  nand GNAME5845(G5845,G58889,G3065);
  nand GNAME5846(G5846,G5832,G59025);
  nand GNAME5847(G5847,G5828,G58873);
  nand GNAME5848(G5848,G5823,G2968);
  nand GNAME5849(G5849,G2969,G3069);
  nand GNAME5850(G5850,G5219,G3067);
  nand GNAME5851(G5851,G58890,G3065);
  nand GNAME5852(G5852,G5832,G59024);
  nand GNAME5853(G5853,G5828,G58874);
  nand GNAME5854(G5854,G5823,G2970);
  nand GNAME5855(G5855,G2971,G3069);
  nand GNAME5856(G5856,G5228,G3067);
  nand GNAME5857(G5857,G58891,G3065);
  nand GNAME5858(G5858,G5832,G59023);
  nand GNAME5859(G5859,G5828,G58875);
  nand GNAME5860(G5860,G5823,G2972);
  nand GNAME5861(G5861,G2973,G3069);
  nand GNAME5862(G5862,G5237,G3067);
  nand GNAME5863(G5863,G58892,G3065);
  nand GNAME5864(G5864,G5832,G59022);
  nand GNAME5865(G5865,G5828,G58876);
  nand GNAME5866(G5866,G5823,G2974);
  nand GNAME5867(G5867,G2975,G3069);
  nand GNAME5868(G5868,G5246,G3067);
  nand GNAME5869(G5869,G58893,G3065);
  nand GNAME5870(G5870,G5832,G59021);
  nand GNAME5871(G5871,G5828,G58877);
  nand GNAME5872(G5872,G5823,G2976);
  nand GNAME5873(G5873,G2977,G3069);
  nand GNAME5874(G5874,G5255,G3067);
  nand GNAME5875(G5875,G58894,G3065);
  nand GNAME5876(G5876,G5832,G59020);
  nand GNAME5877(G5877,G5828,G58878);
  nand GNAME5878(G5878,G5823,G2978);
  nand GNAME5879(G5879,G2979,G3069);
  nand GNAME5880(G5880,G5264,G3067);
  not GNAME5881(G5881,G3070);
  nand GNAME5882(G5882,G58977,G5881);
  nand GNAME5883(G5883,G2836,G3073);
  nand GNAME5884(G5884,G5882,G5883);
  nand GNAME5885(G5885,G3070,G3071);
  and GNAME5886(G5886,G5885,G3803);
  nand GNAME5887(G5887,G3071,G3073);
  nand GNAME5888(G5888,G3074,G3075);
  nand GNAME5889(G5889,G5887,G5888);
  and GNAME5890(G5890,G3070,G58977);
  nor GNAME5891(G5891,G5890,G2805,G3075);
  or GNAME5892(G5892,G3074,G5891);
  nand GNAME5893(G5893,G5892,G2913);
  nand GNAME5894(G5894,G58887,G3072);
  nand GNAME5895(G5895,G5893,G59019);
  nand GNAME5896(G5896,G5889,G58871);
  nand GNAME5897(G5897,G5884,G2962);
  nand GNAME5898(G5898,G2964,G3076);
  nand GNAME5899(G5899,G5188,G3074);
  nand GNAME5900(G5900,G58888,G3072);
  nand GNAME5901(G5901,G5893,G59018);
  nand GNAME5902(G5902,G5889,G58872);
  nand GNAME5903(G5903,G5884,G2966);
  nand GNAME5904(G5904,G2967,G3076);
  nand GNAME5905(G5905,G5210,G3074);
  nand GNAME5906(G5906,G58889,G3072);
  nand GNAME5907(G5907,G5893,G59017);
  nand GNAME5908(G5908,G5889,G58873);
  nand GNAME5909(G5909,G5884,G2968);
  nand GNAME5910(G5910,G2969,G3076);
  nand GNAME5911(G5911,G5219,G3074);
  nand GNAME5912(G5912,G58890,G3072);
  nand GNAME5913(G5913,G5893,G59016);
  nand GNAME5914(G5914,G5889,G58874);
  nand GNAME5915(G5915,G5884,G2970);
  nand GNAME5916(G5916,G2971,G3076);
  nand GNAME5917(G5917,G5228,G3074);
  nand GNAME5918(G5918,G58891,G3072);
  nand GNAME5919(G5919,G5893,G59015);
  nand GNAME5920(G5920,G5889,G58875);
  nand GNAME5921(G5921,G5884,G2972);
  nand GNAME5922(G5922,G2973,G3076);
  nand GNAME5923(G5923,G5237,G3074);
  nand GNAME5924(G5924,G58892,G3072);
  nand GNAME5925(G5925,G5893,G59014);
  nand GNAME5926(G5926,G5889,G58876);
  nand GNAME5927(G5927,G5884,G2974);
  nand GNAME5928(G5928,G2975,G3076);
  nand GNAME5929(G5929,G5246,G3074);
  nand GNAME5930(G5930,G58893,G3072);
  nand GNAME5931(G5931,G5893,G59013);
  nand GNAME5932(G5932,G5889,G58877);
  nand GNAME5933(G5933,G5884,G2976);
  nand GNAME5934(G5934,G2977,G3076);
  nand GNAME5935(G5935,G5255,G3074);
  nand GNAME5936(G5936,G58894,G3072);
  nand GNAME5937(G5937,G5893,G59012);
  nand GNAME5938(G5938,G5889,G58878);
  nand GNAME5939(G5939,G5884,G2978);
  nand GNAME5940(G5940,G2979,G3076);
  nand GNAME5941(G5941,G5264,G3074);
  not GNAME5942(G5942,G3077);
  nand GNAME5943(G5943,G58977,G5942);
  nand GNAME5944(G5944,G2836,G3082);
  nand GNAME5945(G5945,G5943,G5944);
  nand GNAME5946(G5946,G3077,G3078);
  and GNAME5947(G5947,G5946,G3803);
  nand GNAME5948(G5948,G3082,G3077,G3078);
  nand GNAME5949(G5949,G3083,G3084);
  nand GNAME5950(G5950,G5948,G5949);
  and GNAME5951(G5951,G3077,G58977);
  nor GNAME5952(G5952,G5951,G2805,G3084);
  or GNAME5953(G5953,G3083,G5952);
  nand GNAME5954(G5954,G5953,G2913);
  nand GNAME5955(G5955,G58887,G3079);
  nand GNAME5956(G5956,G5954,G59011);
  nand GNAME5957(G5957,G5950,G58871);
  nand GNAME5958(G5958,G5945,G2962);
  nand GNAME5959(G5959,G2964,G3085);
  nand GNAME5960(G5960,G5188,G3083);
  nand GNAME5961(G5961,G58888,G3079);
  nand GNAME5962(G5962,G5954,G59010);
  nand GNAME5963(G5963,G5950,G58872);
  nand GNAME5964(G5964,G5945,G2966);
  nand GNAME5965(G5965,G2967,G3085);
  nand GNAME5966(G5966,G5210,G3083);
  nand GNAME5967(G5967,G58889,G3079);
  nand GNAME5968(G5968,G5954,G59009);
  nand GNAME5969(G5969,G5950,G58873);
  nand GNAME5970(G5970,G5945,G2968);
  nand GNAME5971(G5971,G2969,G3085);
  nand GNAME5972(G5972,G5219,G3083);
  nand GNAME5973(G5973,G58890,G3079);
  nand GNAME5974(G5974,G5954,G59008);
  nand GNAME5975(G5975,G5950,G58874);
  nand GNAME5976(G5976,G5945,G2970);
  nand GNAME5977(G5977,G2971,G3085);
  nand GNAME5978(G5978,G5228,G3083);
  nand GNAME5979(G5979,G58891,G3079);
  nand GNAME5980(G5980,G5954,G59007);
  nand GNAME5981(G5981,G5950,G58875);
  nand GNAME5982(G5982,G5945,G2972);
  nand GNAME5983(G5983,G2973,G3085);
  nand GNAME5984(G5984,G5237,G3083);
  nand GNAME5985(G5985,G58892,G3079);
  nand GNAME5986(G5986,G5954,G59006);
  nand GNAME5987(G5987,G5950,G58876);
  nand GNAME5988(G5988,G5945,G2974);
  nand GNAME5989(G5989,G2975,G3085);
  nand GNAME5990(G5990,G5246,G3083);
  nand GNAME5991(G5991,G58893,G3079);
  nand GNAME5992(G5992,G5954,G59005);
  nand GNAME5993(G5993,G5950,G58877);
  nand GNAME5994(G5994,G5945,G2976);
  nand GNAME5995(G5995,G2977,G3085);
  nand GNAME5996(G5996,G5255,G3083);
  nand GNAME5997(G5997,G58894,G3079);
  nand GNAME5998(G5998,G5954,G59004);
  nand GNAME5999(G5999,G5950,G58878);
  nand GNAME6000(G6000,G5945,G2978);
  nand GNAME6001(G6001,G2979,G3085);
  nand GNAME6002(G6002,G5264,G3083);
  not GNAME6003(G6003,G3086);
  nand GNAME6004(G6004,G58977,G6003);
  nand GNAME6005(G6005,G2836,G3089);
  nand GNAME6006(G6006,G6004,G6005);
  nand GNAME6007(G6007,G3086,G3087);
  and GNAME6008(G6008,G6007,G3803);
  nand GNAME6009(G6009,G3089,G3086,G3087);
  nand GNAME6010(G6010,G3090,G3091);
  nand GNAME6011(G6011,G6009,G6010);
  and GNAME6012(G6012,G3086,G58977);
  nor GNAME6013(G6013,G6012,G2805,G3091);
  or GNAME6014(G6014,G3090,G6013);
  nand GNAME6015(G6015,G6014,G2913);
  nand GNAME6016(G6016,G58887,G3088);
  nand GNAME6017(G6017,G6015,G59003);
  nand GNAME6018(G6018,G6011,G58871);
  nand GNAME6019(G6019,G6006,G2962);
  nand GNAME6020(G6020,G2964,G3092);
  nand GNAME6021(G6021,G5188,G3090);
  nand GNAME6022(G6022,G58888,G3088);
  nand GNAME6023(G6023,G6015,G59002);
  nand GNAME6024(G6024,G6011,G58872);
  nand GNAME6025(G6025,G6006,G2966);
  nand GNAME6026(G6026,G2967,G3092);
  nand GNAME6027(G6027,G5210,G3090);
  nand GNAME6028(G6028,G58889,G3088);
  nand GNAME6029(G6029,G6015,G59001);
  nand GNAME6030(G6030,G6011,G58873);
  nand GNAME6031(G6031,G6006,G2968);
  nand GNAME6032(G6032,G2969,G3092);
  nand GNAME6033(G6033,G5219,G3090);
  nand GNAME6034(G6034,G58890,G3088);
  nand GNAME6035(G6035,G6015,G59000);
  nand GNAME6036(G6036,G6011,G58874);
  nand GNAME6037(G6037,G6006,G2970);
  nand GNAME6038(G6038,G2971,G3092);
  nand GNAME6039(G6039,G5228,G3090);
  nand GNAME6040(G6040,G58891,G3088);
  nand GNAME6041(G6041,G6015,G58999);
  nand GNAME6042(G6042,G6011,G58875);
  nand GNAME6043(G6043,G6006,G2972);
  nand GNAME6044(G6044,G2973,G3092);
  nand GNAME6045(G6045,G5237,G3090);
  nand GNAME6046(G6046,G58892,G3088);
  nand GNAME6047(G6047,G6015,G58998);
  nand GNAME6048(G6048,G6011,G58876);
  nand GNAME6049(G6049,G6006,G2974);
  nand GNAME6050(G6050,G2975,G3092);
  nand GNAME6051(G6051,G5246,G3090);
  nand GNAME6052(G6052,G58893,G3088);
  nand GNAME6053(G6053,G6015,G58997);
  nand GNAME6054(G6054,G6011,G58877);
  nand GNAME6055(G6055,G6006,G2976);
  nand GNAME6056(G6056,G2977,G3092);
  nand GNAME6057(G6057,G5255,G3090);
  nand GNAME6058(G6058,G58894,G3088);
  nand GNAME6059(G6059,G6015,G58996);
  nand GNAME6060(G6060,G6011,G58878);
  nand GNAME6061(G6061,G6006,G2978);
  nand GNAME6062(G6062,G2979,G3092);
  nand GNAME6063(G6063,G5264,G3090);
  not GNAME6064(G6064,G3093);
  nand GNAME6065(G6065,G58977,G6064);
  nand GNAME6066(G6066,G2836,G3096);
  nand GNAME6067(G6067,G6065,G6066);
  nand GNAME6068(G6068,G3093,G3094);
  and GNAME6069(G6069,G6068,G3803);
  nand GNAME6070(G6070,G3096,G3093,G3094);
  nand GNAME6071(G6071,G3097,G3098);
  nand GNAME6072(G6072,G6070,G6071);
  and GNAME6073(G6073,G3093,G58977);
  nor GNAME6074(G6074,G6073,G2805,G3098);
  or GNAME6075(G6075,G3097,G6074);
  nand GNAME6076(G6076,G6075,G2913);
  nand GNAME6077(G6077,G58887,G3095);
  nand GNAME6078(G6078,G6076,G58995);
  nand GNAME6079(G6079,G6072,G58871);
  nand GNAME6080(G6080,G6067,G2962);
  nand GNAME6081(G6081,G2964,G3099);
  nand GNAME6082(G6082,G5188,G3097);
  nand GNAME6083(G6083,G58888,G3095);
  nand GNAME6084(G6084,G6076,G58994);
  nand GNAME6085(G6085,G6072,G58872);
  nand GNAME6086(G6086,G6067,G2966);
  nand GNAME6087(G6087,G2967,G3099);
  nand GNAME6088(G6088,G5210,G3097);
  nand GNAME6089(G6089,G58889,G3095);
  nand GNAME6090(G6090,G6076,G58993);
  nand GNAME6091(G6091,G6072,G58873);
  nand GNAME6092(G6092,G6067,G2968);
  nand GNAME6093(G6093,G2969,G3099);
  nand GNAME6094(G6094,G5219,G3097);
  nand GNAME6095(G6095,G58890,G3095);
  nand GNAME6096(G6096,G6076,G58992);
  nand GNAME6097(G6097,G6072,G58874);
  nand GNAME6098(G6098,G6067,G2970);
  nand GNAME6099(G6099,G2971,G3099);
  nand GNAME6100(G6100,G5228,G3097);
  nand GNAME6101(G6101,G58891,G3095);
  nand GNAME6102(G6102,G6076,G58991);
  nand GNAME6103(G6103,G6072,G58875);
  nand GNAME6104(G6104,G6067,G2972);
  nand GNAME6105(G6105,G2973,G3099);
  nand GNAME6106(G6106,G5237,G3097);
  nand GNAME6107(G6107,G58892,G3095);
  nand GNAME6108(G6108,G6076,G58990);
  nand GNAME6109(G6109,G6072,G58876);
  nand GNAME6110(G6110,G6067,G2974);
  nand GNAME6111(G6111,G2975,G3099);
  nand GNAME6112(G6112,G5246,G3097);
  nand GNAME6113(G6113,G58893,G3095);
  nand GNAME6114(G6114,G6076,G58989);
  nand GNAME6115(G6115,G6072,G58877);
  nand GNAME6116(G6116,G6067,G2976);
  nand GNAME6117(G6117,G2977,G3099);
  nand GNAME6118(G6118,G5255,G3097);
  nand GNAME6119(G6119,G58894,G3095);
  nand GNAME6120(G6120,G6076,G58988);
  nand GNAME6121(G6121,G6072,G58878);
  nand GNAME6122(G6122,G6067,G2978);
  nand GNAME6123(G6123,G2979,G3099);
  nand GNAME6124(G6124,G5264,G3097);
  not GNAME6125(G6125,G3100);
  nand GNAME6126(G6126,G58977,G6125);
  nand GNAME6127(G6127,G2836,G3103);
  nand GNAME6128(G6128,G6126,G6127);
  nand GNAME6129(G6129,G3100,G3101);
  and GNAME6130(G6130,G6129,G3803);
  nand GNAME6131(G6131,G3101,G3103);
  nand GNAME6132(G6132,G3104,G3105);
  nand GNAME6133(G6133,G6131,G6132);
  and GNAME6134(G6134,G3100,G58977);
  nor GNAME6135(G6135,G6134,G2805,G3104);
  or GNAME6136(G6136,G3105,G6135);
  nand GNAME6137(G6137,G6136,G2913);
  nand GNAME6138(G6138,G58887,G3102);
  nand GNAME6139(G6139,G6137,G58987);
  nand GNAME6140(G6140,G6133,G58871);
  nand GNAME6141(G6141,G6128,G2962);
  nand GNAME6142(G6142,G5188,G3105);
  nand GNAME6143(G6143,G2964,G3106);
  nand GNAME6144(G6144,G58888,G3102);
  nand GNAME6145(G6145,G6137,G58986);
  nand GNAME6146(G6146,G6133,G58872);
  nand GNAME6147(G6147,G6128,G2966);
  nand GNAME6148(G6148,G5210,G3105);
  nand GNAME6149(G6149,G2967,G3106);
  nand GNAME6150(G6150,G58889,G3102);
  nand GNAME6151(G6151,G6137,G58985);
  nand GNAME6152(G6152,G6133,G58873);
  nand GNAME6153(G6153,G6128,G2968);
  nand GNAME6154(G6154,G5219,G3105);
  nand GNAME6155(G6155,G2969,G3106);
  nand GNAME6156(G6156,G58890,G3102);
  nand GNAME6157(G6157,G6137,G58984);
  nand GNAME6158(G6158,G6133,G58874);
  nand GNAME6159(G6159,G6128,G2970);
  nand GNAME6160(G6160,G5228,G3105);
  nand GNAME6161(G6161,G2971,G3106);
  nand GNAME6162(G6162,G58891,G3102);
  nand GNAME6163(G6163,G6137,G58983);
  nand GNAME6164(G6164,G6133,G58875);
  nand GNAME6165(G6165,G6128,G2972);
  nand GNAME6166(G6166,G5237,G3105);
  nand GNAME6167(G6167,G2973,G3106);
  nand GNAME6168(G6168,G58892,G3102);
  nand GNAME6169(G6169,G6137,G58982);
  nand GNAME6170(G6170,G6133,G58876);
  nand GNAME6171(G6171,G6128,G2974);
  nand GNAME6172(G6172,G5246,G3105);
  nand GNAME6173(G6173,G2975,G3106);
  nand GNAME6174(G6174,G58893,G3102);
  nand GNAME6175(G6175,G6137,G58981);
  nand GNAME6176(G6176,G6133,G58877);
  nand GNAME6177(G6177,G6128,G2976);
  nand GNAME6178(G6178,G5255,G3105);
  nand GNAME6179(G6179,G2977,G3106);
  nand GNAME6180(G6180,G58894,G3102);
  nand GNAME6181(G6181,G6137,G58980);
  nand GNAME6182(G6182,G6133,G58878);
  nand GNAME6183(G6183,G6128,G2978);
  nand GNAME6184(G6184,G5264,G3105);
  nand GNAME6185(G6185,G2979,G3106);
  nand GNAME6186(G6186,G3108,G2797,G2802);
  or GNAME6187(G6187,G59346,G59347);
  nand GNAME6188(G6188,G2804,G6186);
  nand GNAME6189(G6189,G2792,G2789);
  nand GNAME6190(G6190,G2817,G3109);
  nand GNAME6191(G6191,G1590,G58978);
  nand GNAME6192(G6192,G2838,G3958,G3980);
  nand GNAME6193(G6193,G58976,G20108,G2805);
  nand GNAME6194(G6194,G2790,G6193);
  or GNAME6195(G6195,G3109,G3801);
  nand GNAME6196(G6196,G20108,G2910);
  nand GNAME6197(G6197,G6196,G6194,G6195);
  nand GNAME6198(G6198,G3111,G2752,G58979);
  nand GNAME6199(G6199,G6198,G3807);
  nand GNAME6200(G6200,G3813,G3110);
  nand GNAME6201(G6201,G6200,G58978);
  nand GNAME6202(G6202,G3110,G6199);
  nand GNAME6203(G6203,G2842,G2752,G58978);
  nand GNAME6204(G6204,G2790,G2943);
  or GNAME6205(G6205,G2837,G3110);
  or GNAME6206(G6206,G58941,G58943);
  nand GNAME6207(G6207,G6206,G3774);
  nand GNAME6208(G6208,G2751,G59349);
  nand GNAME6209(G6209,G2809,G34);
  nand GNAME6210(G6210,G59349,G3113,G6209);
  or GNAME6211(G6211,G2752,G2808);
  nand GNAME6212(G6212,G2752,G58941);
  or GNAME6213(G6213,G1590,G33);
  nand GNAME6214(G6214,G2815,G58941);
  nand GNAME6215(G6215,G2751,G6208);
  nand GNAME6216(G6216,G58943,G3112,G6215);
  nand GNAME6217(G6217,G6216,G2820);
  or GNAME6218(G6218,G3113,G2815,G2751);
  nand GNAME6219(G6219,G3787,G58940);
  nand GNAME6220(G6220,G59311,G3114);
  nand GNAME6221(G6221,G59310,G3115);
  nand GNAME6222(G6222,G3787,G58939);
  nand GNAME6223(G6223,G59311,G3115);
  nand GNAME6224(G6224,G59312,G3114);
  nand GNAME6225(G6225,G3787,G58938);
  nand GNAME6226(G6226,G59312,G3115);
  nand GNAME6227(G6227,G59313,G3114);
  nand GNAME6228(G6228,G3787,G58937);
  nand GNAME6229(G6229,G59313,G3115);
  nand GNAME6230(G6230,G59314,G3114);
  nand GNAME6231(G6231,G3787,G58936);
  nand GNAME6232(G6232,G59314,G3115);
  nand GNAME6233(G6233,G59315,G3114);
  nand GNAME6234(G6234,G3787,G58935);
  nand GNAME6235(G6235,G59315,G3115);
  nand GNAME6236(G6236,G59316,G3114);
  nand GNAME6237(G6237,G3787,G58934);
  nand GNAME6238(G6238,G59316,G3115);
  nand GNAME6239(G6239,G59317,G3114);
  nand GNAME6240(G6240,G3787,G58933);
  nand GNAME6241(G6241,G59317,G3115);
  nand GNAME6242(G6242,G59318,G3114);
  nand GNAME6243(G6243,G3787,G58932);
  nand GNAME6244(G6244,G59318,G3115);
  nand GNAME6245(G6245,G59319,G3114);
  nand GNAME6246(G6246,G3787,G58931);
  nand GNAME6247(G6247,G59319,G3115);
  nand GNAME6248(G6248,G59320,G3114);
  nand GNAME6249(G6249,G3787,G58930);
  nand GNAME6250(G6250,G59320,G3115);
  nand GNAME6251(G6251,G59321,G3114);
  nand GNAME6252(G6252,G3787,G58929);
  nand GNAME6253(G6253,G59321,G3115);
  nand GNAME6254(G6254,G59322,G3114);
  nand GNAME6255(G6255,G3787,G58928);
  nand GNAME6256(G6256,G59322,G3115);
  nand GNAME6257(G6257,G59323,G3114);
  nand GNAME6258(G6258,G3787,G58927);
  nand GNAME6259(G6259,G59323,G3115);
  nand GNAME6260(G6260,G59324,G3114);
  nand GNAME6261(G6261,G3787,G58926);
  nand GNAME6262(G6262,G59324,G3115);
  nand GNAME6263(G6263,G59325,G3114);
  nand GNAME6264(G6264,G3787,G58925);
  nand GNAME6265(G6265,G59325,G3115);
  nand GNAME6266(G6266,G59326,G3114);
  nand GNAME6267(G6267,G3787,G58924);
  nand GNAME6268(G6268,G59326,G3115);
  nand GNAME6269(G6269,G59327,G3114);
  nand GNAME6270(G6270,G3787,G58923);
  nand GNAME6271(G6271,G59327,G3115);
  nand GNAME6272(G6272,G59328,G3114);
  nand GNAME6273(G6273,G3787,G58922);
  nand GNAME6274(G6274,G59328,G3115);
  nand GNAME6275(G6275,G59329,G3114);
  nand GNAME6276(G6276,G3787,G58921);
  nand GNAME6277(G6277,G59329,G3115);
  nand GNAME6278(G6278,G59330,G3114);
  nand GNAME6279(G6279,G3787,G58920);
  nand GNAME6280(G6280,G59330,G3115);
  nand GNAME6281(G6281,G59331,G3114);
  nand GNAME6282(G6282,G3787,G58919);
  nand GNAME6283(G6283,G59331,G3115);
  nand GNAME6284(G6284,G59332,G3114);
  nand GNAME6285(G6285,G3787,G58918);
  nand GNAME6286(G6286,G59332,G3115);
  nand GNAME6287(G6287,G59333,G3114);
  nand GNAME6288(G6288,G3787,G58917);
  nand GNAME6289(G6289,G59333,G3115);
  nand GNAME6290(G6290,G59334,G3114);
  nand GNAME6291(G6291,G3787,G58916);
  nand GNAME6292(G6292,G59334,G3115);
  nand GNAME6293(G6293,G59335,G3114);
  nand GNAME6294(G6294,G3787,G58915);
  nand GNAME6295(G6295,G59335,G3115);
  nand GNAME6296(G6296,G59336,G3114);
  nand GNAME6297(G6297,G3787,G58914);
  nand GNAME6298(G6298,G59336,G3115);
  nand GNAME6299(G6299,G59337,G3114);
  nand GNAME6300(G6300,G3787,G58913);
  nand GNAME6301(G6301,G59337,G3115);
  nand GNAME6302(G6302,G59338,G3114);
  nand GNAME6303(G6303,G3787,G58912);
  nand GNAME6304(G6304,G59338,G3115);
  nand GNAME6305(G6305,G59339,G3114);
  nand GNAME6306(G6306,G3787,G58911);
  nand GNAME6307(G6307,G59339,G3115);
  nand GNAME6308(G6308,G59340,G3114);
  nand GNAME6309(G6309,G59092,G3118);
  nand GNAME6310(G6310,G59084,G3121);
  nand GNAME6311(G6311,G59076,G3122);
  nand GNAME6312(G6312,G59068,G3124);
  nand GNAME6313(G6313,G59060,G3125);
  nand GNAME6314(G6314,G59052,G3127);
  nand GNAME6315(G6315,G59044,G3128);
  nand GNAME6316(G6316,G59036,G3130);
  nand GNAME6317(G6317,G59028,G3132);
  nand GNAME6318(G6318,G59020,G3133);
  nand GNAME6319(G6319,G59012,G3134);
  nand GNAME6320(G6320,G59004,G3135);
  nand GNAME6321(G6321,G58996,G3136);
  nand GNAME6322(G6322,G58988,G3137);
  nand GNAME6323(G6323,G58980,G3138);
  nand GNAME6324(G6324,G59100,G3139);
  nand GNAME6325(G6325,G59093,G3118);
  nand GNAME6326(G6326,G59085,G3121);
  nand GNAME6327(G6327,G59077,G3122);
  nand GNAME6328(G6328,G59069,G3124);
  nand GNAME6329(G6329,G59061,G3125);
  nand GNAME6330(G6330,G59053,G3127);
  nand GNAME6331(G6331,G59045,G3128);
  nand GNAME6332(G6332,G59037,G3130);
  nand GNAME6333(G6333,G59029,G3132);
  nand GNAME6334(G6334,G59021,G3133);
  nand GNAME6335(G6335,G59013,G3134);
  nand GNAME6336(G6336,G59005,G3135);
  nand GNAME6337(G6337,G58997,G3136);
  nand GNAME6338(G6338,G58989,G3137);
  nand GNAME6339(G6339,G58981,G3138);
  nand GNAME6340(G6340,G59101,G3139);
  nand GNAME6341(G6341,G59094,G3118);
  nand GNAME6342(G6342,G59086,G3121);
  nand GNAME6343(G6343,G59078,G3122);
  nand GNAME6344(G6344,G59070,G3124);
  nand GNAME6345(G6345,G59062,G3125);
  nand GNAME6346(G6346,G59054,G3127);
  nand GNAME6347(G6347,G59046,G3128);
  nand GNAME6348(G6348,G59038,G3130);
  nand GNAME6349(G6349,G59030,G3132);
  nand GNAME6350(G6350,G59022,G3133);
  nand GNAME6351(G6351,G59014,G3134);
  nand GNAME6352(G6352,G59006,G3135);
  nand GNAME6353(G6353,G58998,G3136);
  nand GNAME6354(G6354,G58990,G3137);
  nand GNAME6355(G6355,G58982,G3138);
  nand GNAME6356(G6356,G59102,G3139);
  nand GNAME6357(G6357,G59095,G3118);
  nand GNAME6358(G6358,G59087,G3121);
  nand GNAME6359(G6359,G59079,G3122);
  nand GNAME6360(G6360,G59071,G3124);
  nand GNAME6361(G6361,G59063,G3125);
  nand GNAME6362(G6362,G59055,G3127);
  nand GNAME6363(G6363,G59047,G3128);
  nand GNAME6364(G6364,G59039,G3130);
  nand GNAME6365(G6365,G59031,G3132);
  nand GNAME6366(G6366,G59023,G3133);
  nand GNAME6367(G6367,G59015,G3134);
  nand GNAME6368(G6368,G59007,G3135);
  nand GNAME6369(G6369,G58999,G3136);
  nand GNAME6370(G6370,G58991,G3137);
  nand GNAME6371(G6371,G58983,G3138);
  nand GNAME6372(G6372,G59103,G3139);
  nand GNAME6373(G6373,G59096,G3118);
  nand GNAME6374(G6374,G59088,G3121);
  nand GNAME6375(G6375,G59080,G3122);
  nand GNAME6376(G6376,G59072,G3124);
  nand GNAME6377(G6377,G59064,G3125);
  nand GNAME6378(G6378,G59056,G3127);
  nand GNAME6379(G6379,G59048,G3128);
  nand GNAME6380(G6380,G59040,G3130);
  nand GNAME6381(G6381,G59032,G3132);
  nand GNAME6382(G6382,G59024,G3133);
  nand GNAME6383(G6383,G59016,G3134);
  nand GNAME6384(G6384,G59008,G3135);
  nand GNAME6385(G6385,G59000,G3136);
  nand GNAME6386(G6386,G58992,G3137);
  nand GNAME6387(G6387,G58984,G3138);
  nand GNAME6388(G6388,G59104,G3139);
  nand GNAME6389(G6389,G59105,G3139);
  nand GNAME6390(G6390,G59097,G3118);
  nand GNAME6391(G6391,G59089,G3121);
  nand GNAME6392(G6392,G59081,G3122);
  nand GNAME6393(G6393,G59073,G3124);
  nand GNAME6394(G6394,G59065,G3125);
  nand GNAME6395(G6395,G59057,G3127);
  nand GNAME6396(G6396,G59049,G3128);
  nand GNAME6397(G6397,G59041,G3130);
  nand GNAME6398(G6398,G59033,G3132);
  nand GNAME6399(G6399,G59025,G3133);
  nand GNAME6400(G6400,G59017,G3134);
  nand GNAME6401(G6401,G59009,G3135);
  nand GNAME6402(G6402,G59001,G3136);
  nand GNAME6403(G6403,G58993,G3137);
  nand GNAME6404(G6404,G58985,G3138);
  nand GNAME6405(G6405,G59106,G3139);
  nand GNAME6406(G6406,G59098,G3118);
  nand GNAME6407(G6407,G59090,G3121);
  nand GNAME6408(G6408,G59082,G3122);
  nand GNAME6409(G6409,G59074,G3124);
  nand GNAME6410(G6410,G59066,G3125);
  nand GNAME6411(G6411,G59058,G3127);
  nand GNAME6412(G6412,G59050,G3128);
  nand GNAME6413(G6413,G59042,G3130);
  nand GNAME6414(G6414,G59034,G3132);
  nand GNAME6415(G6415,G59026,G3133);
  nand GNAME6416(G6416,G59018,G3134);
  nand GNAME6417(G6417,G59010,G3135);
  nand GNAME6418(G6418,G59002,G3136);
  nand GNAME6419(G6419,G58994,G3137);
  nand GNAME6420(G6420,G58986,G3138);
  nand GNAME6421(G6421,G59107,G3139);
  nand GNAME6422(G6422,G59099,G3118);
  nand GNAME6423(G6423,G59091,G3121);
  nand GNAME6424(G6424,G59083,G3122);
  nand GNAME6425(G6425,G59075,G3124);
  nand GNAME6426(G6426,G59067,G3125);
  nand GNAME6427(G6427,G59059,G3127);
  nand GNAME6428(G6428,G59051,G3128);
  nand GNAME6429(G6429,G59043,G3130);
  nand GNAME6430(G6430,G59035,G3132);
  nand GNAME6431(G6431,G59027,G3133);
  nand GNAME6432(G6432,G59019,G3134);
  nand GNAME6433(G6433,G59011,G3135);
  nand GNAME6434(G6434,G59003,G3136);
  nand GNAME6435(G6435,G58995,G3137);
  nand GNAME6436(G6436,G58987,G3138);
  not GNAME6437(G6437,G3140);
  nand GNAME6438(G6438,G59092,G3142);
  nand GNAME6439(G6439,G59084,G3143);
  nand GNAME6440(G6440,G59076,G3144);
  nand GNAME6441(G6441,G59068,G3146);
  nand GNAME6442(G6442,G59060,G3147);
  nand GNAME6443(G6443,G59052,G3148);
  nand GNAME6444(G6444,G59044,G3149);
  nand GNAME6445(G6445,G59036,G3151);
  nand GNAME6446(G6446,G59028,G3152);
  nand GNAME6447(G6447,G59020,G3153);
  nand GNAME6448(G6448,G59012,G3154);
  nand GNAME6449(G6449,G59004,G3156);
  nand GNAME6450(G6450,G58996,G3157);
  nand GNAME6451(G6451,G58988,G3158);
  nand GNAME6452(G6452,G58980,G3159);
  nand GNAME6453(G6453,G59100,G3160);
  nand GNAME6454(G6454,G59093,G3142);
  nand GNAME6455(G6455,G59085,G3143);
  nand GNAME6456(G6456,G59077,G3144);
  nand GNAME6457(G6457,G59069,G3146);
  nand GNAME6458(G6458,G59061,G3147);
  nand GNAME6459(G6459,G59053,G3148);
  nand GNAME6460(G6460,G59045,G3149);
  nand GNAME6461(G6461,G59037,G3151);
  nand GNAME6462(G6462,G59029,G3152);
  nand GNAME6463(G6463,G59021,G3153);
  nand GNAME6464(G6464,G59013,G3154);
  nand GNAME6465(G6465,G59005,G3156);
  nand GNAME6466(G6466,G58997,G3157);
  nand GNAME6467(G6467,G58989,G3158);
  nand GNAME6468(G6468,G58981,G3159);
  nand GNAME6469(G6469,G59101,G3160);
  nand GNAME6470(G6470,G59094,G3142);
  nand GNAME6471(G6471,G59086,G3143);
  nand GNAME6472(G6472,G59078,G3144);
  nand GNAME6473(G6473,G59070,G3146);
  nand GNAME6474(G6474,G59062,G3147);
  nand GNAME6475(G6475,G59054,G3148);
  nand GNAME6476(G6476,G59046,G3149);
  nand GNAME6477(G6477,G59038,G3151);
  nand GNAME6478(G6478,G59030,G3152);
  nand GNAME6479(G6479,G59022,G3153);
  nand GNAME6480(G6480,G59014,G3154);
  nand GNAME6481(G6481,G59006,G3156);
  nand GNAME6482(G6482,G58998,G3157);
  nand GNAME6483(G6483,G58990,G3158);
  nand GNAME6484(G6484,G58982,G3159);
  nand GNAME6485(G6485,G59102,G3160);
  nand GNAME6486(G6486,G59095,G3142);
  nand GNAME6487(G6487,G59087,G3143);
  nand GNAME6488(G6488,G59079,G3144);
  nand GNAME6489(G6489,G59071,G3146);
  nand GNAME6490(G6490,G59063,G3147);
  nand GNAME6491(G6491,G59055,G3148);
  nand GNAME6492(G6492,G59047,G3149);
  nand GNAME6493(G6493,G59039,G3151);
  nand GNAME6494(G6494,G59031,G3152);
  nand GNAME6495(G6495,G59023,G3153);
  nand GNAME6496(G6496,G59015,G3154);
  nand GNAME6497(G6497,G59007,G3156);
  nand GNAME6498(G6498,G58999,G3157);
  nand GNAME6499(G6499,G58991,G3158);
  nand GNAME6500(G6500,G58983,G3159);
  nand GNAME6501(G6501,G59103,G3160);
  nand GNAME6502(G6502,G59096,G3142);
  nand GNAME6503(G6503,G59088,G3143);
  nand GNAME6504(G6504,G59080,G3144);
  nand GNAME6505(G6505,G59072,G3146);
  nand GNAME6506(G6506,G59064,G3147);
  nand GNAME6507(G6507,G59056,G3148);
  nand GNAME6508(G6508,G59048,G3149);
  nand GNAME6509(G6509,G59040,G3151);
  nand GNAME6510(G6510,G59032,G3152);
  nand GNAME6511(G6511,G59024,G3153);
  nand GNAME6512(G6512,G59016,G3154);
  nand GNAME6513(G6513,G59008,G3156);
  nand GNAME6514(G6514,G59000,G3157);
  nand GNAME6515(G6515,G58992,G3158);
  nand GNAME6516(G6516,G58984,G3159);
  nand GNAME6517(G6517,G59104,G3160);
  nand GNAME6518(G6518,G59105,G3160);
  nand GNAME6519(G6519,G59097,G3142);
  nand GNAME6520(G6520,G59089,G3143);
  nand GNAME6521(G6521,G59081,G3144);
  nand GNAME6522(G6522,G59073,G3146);
  nand GNAME6523(G6523,G59065,G3147);
  nand GNAME6524(G6524,G59057,G3148);
  nand GNAME6525(G6525,G59049,G3149);
  nand GNAME6526(G6526,G59041,G3151);
  nand GNAME6527(G6527,G59033,G3152);
  nand GNAME6528(G6528,G59025,G3153);
  nand GNAME6529(G6529,G59017,G3154);
  nand GNAME6530(G6530,G59009,G3156);
  nand GNAME6531(G6531,G59001,G3157);
  nand GNAME6532(G6532,G58993,G3158);
  nand GNAME6533(G6533,G58985,G3159);
  nand GNAME6534(G6534,G59106,G3160);
  nand GNAME6535(G6535,G59098,G3142);
  nand GNAME6536(G6536,G59090,G3143);
  nand GNAME6537(G6537,G59082,G3144);
  nand GNAME6538(G6538,G59074,G3146);
  nand GNAME6539(G6539,G59066,G3147);
  nand GNAME6540(G6540,G59058,G3148);
  nand GNAME6541(G6541,G59050,G3149);
  nand GNAME6542(G6542,G59042,G3151);
  nand GNAME6543(G6543,G59034,G3152);
  nand GNAME6544(G6544,G59026,G3153);
  nand GNAME6545(G6545,G59018,G3154);
  nand GNAME6546(G6546,G59010,G3156);
  nand GNAME6547(G6547,G59002,G3157);
  nand GNAME6548(G6548,G58994,G3158);
  nand GNAME6549(G6549,G58986,G3159);
  nand GNAME6550(G6550,G59107,G3160);
  nand GNAME6551(G6551,G59099,G3142);
  nand GNAME6552(G6552,G59091,G3143);
  nand GNAME6553(G6553,G59083,G3144);
  nand GNAME6554(G6554,G59075,G3146);
  nand GNAME6555(G6555,G59067,G3147);
  nand GNAME6556(G6556,G59059,G3148);
  nand GNAME6557(G6557,G59051,G3149);
  nand GNAME6558(G6558,G59043,G3151);
  nand GNAME6559(G6559,G59035,G3152);
  nand GNAME6560(G6560,G59027,G3153);
  nand GNAME6561(G6561,G59019,G3154);
  nand GNAME6562(G6562,G59011,G3156);
  nand GNAME6563(G6563,G59003,G3157);
  nand GNAME6564(G6564,G58995,G3158);
  nand GNAME6565(G6565,G58987,G3159);
  nand GNAME6566(G6566,G59092,G2990);
  nand GNAME6567(G6567,G59084,G3001);
  nand GNAME6568(G6568,G59076,G3009);
  nand GNAME6569(G6569,G59068,G3019);
  nand GNAME6570(G6570,G59060,G3028);
  nand GNAME6571(G6571,G59052,G3035);
  nand GNAME6572(G6572,G59044,G3042);
  nand GNAME6573(G6573,G59036,G3053);
  nand GNAME6574(G6574,G59028,G3060);
  nand GNAME6575(G6575,G59020,G3069);
  nand GNAME6576(G6576,G59012,G3076);
  nand GNAME6577(G6577,G59004,G3085);
  nand GNAME6578(G6578,G58996,G3092);
  nand GNAME6579(G6579,G58988,G3099);
  nand GNAME6580(G6580,G58980,G3106);
  nand GNAME6581(G6581,G59100,G2963);
  nand GNAME6582(G6582,G3600,G3601,G3602,G3603);
  nand GNAME6583(G6583,G59093,G2990);
  nand GNAME6584(G6584,G59085,G3001);
  nand GNAME6585(G6585,G59077,G3009);
  nand GNAME6586(G6586,G59069,G3019);
  nand GNAME6587(G6587,G59061,G3028);
  nand GNAME6588(G6588,G59053,G3035);
  nand GNAME6589(G6589,G59045,G3042);
  nand GNAME6590(G6590,G59037,G3053);
  nand GNAME6591(G6591,G59029,G3060);
  nand GNAME6592(G6592,G59021,G3069);
  nand GNAME6593(G6593,G59013,G3076);
  nand GNAME6594(G6594,G59005,G3085);
  nand GNAME6595(G6595,G58997,G3092);
  nand GNAME6596(G6596,G58989,G3099);
  nand GNAME6597(G6597,G58981,G3106);
  nand GNAME6598(G6598,G59101,G2963);
  nand GNAME6599(G6599,G3604,G3605,G3606,G3607);
  nand GNAME6600(G6600,G59094,G2990);
  nand GNAME6601(G6601,G59086,G3001);
  nand GNAME6602(G6602,G59078,G3009);
  nand GNAME6603(G6603,G59070,G3019);
  nand GNAME6604(G6604,G59062,G3028);
  nand GNAME6605(G6605,G59054,G3035);
  nand GNAME6606(G6606,G59046,G3042);
  nand GNAME6607(G6607,G59038,G3053);
  nand GNAME6608(G6608,G59030,G3060);
  nand GNAME6609(G6609,G59022,G3069);
  nand GNAME6610(G6610,G59014,G3076);
  nand GNAME6611(G6611,G59006,G3085);
  nand GNAME6612(G6612,G58998,G3092);
  nand GNAME6613(G6613,G58990,G3099);
  nand GNAME6614(G6614,G58982,G3106);
  nand GNAME6615(G6615,G59102,G2963);
  nand GNAME6616(G6616,G3608,G3609,G3610,G3611);
  nand GNAME6617(G6617,G59095,G2990);
  nand GNAME6618(G6618,G59087,G3001);
  nand GNAME6619(G6619,G59079,G3009);
  nand GNAME6620(G6620,G59071,G3019);
  nand GNAME6621(G6621,G59063,G3028);
  nand GNAME6622(G6622,G59055,G3035);
  nand GNAME6623(G6623,G59047,G3042);
  nand GNAME6624(G6624,G59039,G3053);
  nand GNAME6625(G6625,G59031,G3060);
  nand GNAME6626(G6626,G59023,G3069);
  nand GNAME6627(G6627,G59015,G3076);
  nand GNAME6628(G6628,G59007,G3085);
  nand GNAME6629(G6629,G58999,G3092);
  nand GNAME6630(G6630,G58991,G3099);
  nand GNAME6631(G6631,G58983,G3106);
  nand GNAME6632(G6632,G59103,G2963);
  nand GNAME6633(G6633,G3612,G3613,G3614,G3615);
  nand GNAME6634(G6634,G59096,G2990);
  nand GNAME6635(G6635,G59088,G3001);
  nand GNAME6636(G6636,G59080,G3009);
  nand GNAME6637(G6637,G59072,G3019);
  nand GNAME6638(G6638,G59064,G3028);
  nand GNAME6639(G6639,G59056,G3035);
  nand GNAME6640(G6640,G59048,G3042);
  nand GNAME6641(G6641,G59040,G3053);
  nand GNAME6642(G6642,G59032,G3060);
  nand GNAME6643(G6643,G59024,G3069);
  nand GNAME6644(G6644,G59016,G3076);
  nand GNAME6645(G6645,G59008,G3085);
  nand GNAME6646(G6646,G59000,G3092);
  nand GNAME6647(G6647,G58992,G3099);
  nand GNAME6648(G6648,G58984,G3106);
  nand GNAME6649(G6649,G59104,G2963);
  nand GNAME6650(G6650,G3616,G3617,G3618,G3619);
  nand GNAME6651(G6651,G59105,G2963);
  nand GNAME6652(G6652,G59097,G2990);
  nand GNAME6653(G6653,G59089,G3001);
  nand GNAME6654(G6654,G59081,G3009);
  nand GNAME6655(G6655,G59073,G3019);
  nand GNAME6656(G6656,G59065,G3028);
  nand GNAME6657(G6657,G59057,G3035);
  nand GNAME6658(G6658,G59049,G3042);
  nand GNAME6659(G6659,G59041,G3053);
  nand GNAME6660(G6660,G59033,G3060);
  nand GNAME6661(G6661,G59025,G3069);
  nand GNAME6662(G6662,G59017,G3076);
  nand GNAME6663(G6663,G59009,G3085);
  nand GNAME6664(G6664,G59001,G3092);
  nand GNAME6665(G6665,G58993,G3099);
  nand GNAME6666(G6666,G58985,G3106);
  nand GNAME6667(G6667,G3620,G3621,G3622,G3623);
  nand GNAME6668(G6668,G59106,G2963);
  nand GNAME6669(G6669,G59098,G2990);
  nand GNAME6670(G6670,G59090,G3001);
  nand GNAME6671(G6671,G59082,G3009);
  nand GNAME6672(G6672,G59074,G3019);
  nand GNAME6673(G6673,G59066,G3028);
  nand GNAME6674(G6674,G59058,G3035);
  nand GNAME6675(G6675,G59050,G3042);
  nand GNAME6676(G6676,G59042,G3053);
  nand GNAME6677(G6677,G59034,G3060);
  nand GNAME6678(G6678,G59026,G3069);
  nand GNAME6679(G6679,G59018,G3076);
  nand GNAME6680(G6680,G59010,G3085);
  nand GNAME6681(G6681,G59002,G3092);
  nand GNAME6682(G6682,G58994,G3099);
  nand GNAME6683(G6683,G58986,G3106);
  nand GNAME6684(G6684,G3624,G3625,G3626,G3627);
  nand GNAME6685(G6685,G59107,G2963);
  nand GNAME6686(G6686,G59099,G2990);
  nand GNAME6687(G6687,G59091,G3001);
  nand GNAME6688(G6688,G59083,G3009);
  nand GNAME6689(G6689,G59075,G3019);
  nand GNAME6690(G6690,G59067,G3028);
  nand GNAME6691(G6691,G59059,G3035);
  nand GNAME6692(G6692,G59051,G3042);
  nand GNAME6693(G6693,G59043,G3053);
  nand GNAME6694(G6694,G59035,G3060);
  nand GNAME6695(G6695,G59027,G3069);
  nand GNAME6696(G6696,G59019,G3076);
  nand GNAME6697(G6697,G59011,G3085);
  nand GNAME6698(G6698,G59003,G3092);
  nand GNAME6699(G6699,G58995,G3099);
  nand GNAME6700(G6700,G58987,G3106);
  nand GNAME6701(G6701,G3628,G3629,G3630,G3631);
  nand GNAME6702(G6702,G59092,G3163);
  nand GNAME6703(G6703,G59084,G3166);
  nand GNAME6704(G6704,G59076,G3168);
  nand GNAME6705(G6705,G59068,G3171);
  nand GNAME6706(G6706,G59060,G3172);
  nand GNAME6707(G6707,G59052,G3173);
  nand GNAME6708(G6708,G59044,G3174);
  nand GNAME6709(G6709,G59036,G3176);
  nand GNAME6710(G6710,G59028,G3177);
  nand GNAME6711(G6711,G59020,G3178);
  nand GNAME6712(G6712,G59012,G3179);
  nand GNAME6713(G6713,G59004,G3181);
  nand GNAME6714(G6714,G58996,G3182);
  nand GNAME6715(G6715,G58988,G3183);
  nand GNAME6716(G6716,G58980,G3184);
  nand GNAME6717(G6717,G59100,G3185);
  nand GNAME6718(G6718,G3632,G3633,G3634,G3635);
  nand GNAME6719(G6719,G59093,G3163);
  nand GNAME6720(G6720,G59085,G3166);
  nand GNAME6721(G6721,G59077,G3168);
  nand GNAME6722(G6722,G59069,G3171);
  nand GNAME6723(G6723,G59061,G3172);
  nand GNAME6724(G6724,G59053,G3173);
  nand GNAME6725(G6725,G59045,G3174);
  nand GNAME6726(G6726,G59037,G3176);
  nand GNAME6727(G6727,G59029,G3177);
  nand GNAME6728(G6728,G59021,G3178);
  nand GNAME6729(G6729,G59013,G3179);
  nand GNAME6730(G6730,G59005,G3181);
  nand GNAME6731(G6731,G58997,G3182);
  nand GNAME6732(G6732,G58989,G3183);
  nand GNAME6733(G6733,G58981,G3184);
  nand GNAME6734(G6734,G59101,G3185);
  nand GNAME6735(G6735,G3636,G3637,G3638,G3639);
  nand GNAME6736(G6736,G59094,G3163);
  nand GNAME6737(G6737,G59086,G3166);
  nand GNAME6738(G6738,G59078,G3168);
  nand GNAME6739(G6739,G59070,G3171);
  nand GNAME6740(G6740,G59062,G3172);
  nand GNAME6741(G6741,G59054,G3173);
  nand GNAME6742(G6742,G59046,G3174);
  nand GNAME6743(G6743,G59038,G3176);
  nand GNAME6744(G6744,G59030,G3177);
  nand GNAME6745(G6745,G59022,G3178);
  nand GNAME6746(G6746,G59014,G3179);
  nand GNAME6747(G6747,G59006,G3181);
  nand GNAME6748(G6748,G58998,G3182);
  nand GNAME6749(G6749,G58990,G3183);
  nand GNAME6750(G6750,G58982,G3184);
  nand GNAME6751(G6751,G59102,G3185);
  nand GNAME6752(G6752,G3640,G3641,G3642,G3643);
  nand GNAME6753(G6753,G59095,G3163);
  nand GNAME6754(G6754,G59087,G3166);
  nand GNAME6755(G6755,G59079,G3168);
  nand GNAME6756(G6756,G59071,G3171);
  nand GNAME6757(G6757,G59063,G3172);
  nand GNAME6758(G6758,G59055,G3173);
  nand GNAME6759(G6759,G59047,G3174);
  nand GNAME6760(G6760,G59039,G3176);
  nand GNAME6761(G6761,G59031,G3177);
  nand GNAME6762(G6762,G59023,G3178);
  nand GNAME6763(G6763,G59015,G3179);
  nand GNAME6764(G6764,G59007,G3181);
  nand GNAME6765(G6765,G58999,G3182);
  nand GNAME6766(G6766,G58991,G3183);
  nand GNAME6767(G6767,G58983,G3184);
  nand GNAME6768(G6768,G59103,G3185);
  nand GNAME6769(G6769,G3644,G3645,G3646,G3647);
  nand GNAME6770(G6770,G59096,G3163);
  nand GNAME6771(G6771,G59088,G3166);
  nand GNAME6772(G6772,G59080,G3168);
  nand GNAME6773(G6773,G59072,G3171);
  nand GNAME6774(G6774,G59064,G3172);
  nand GNAME6775(G6775,G59056,G3173);
  nand GNAME6776(G6776,G59048,G3174);
  nand GNAME6777(G6777,G59040,G3176);
  nand GNAME6778(G6778,G59032,G3177);
  nand GNAME6779(G6779,G59024,G3178);
  nand GNAME6780(G6780,G59016,G3179);
  nand GNAME6781(G6781,G59008,G3181);
  nand GNAME6782(G6782,G59000,G3182);
  nand GNAME6783(G6783,G58992,G3183);
  nand GNAME6784(G6784,G58984,G3184);
  nand GNAME6785(G6785,G59104,G3185);
  nand GNAME6786(G6786,G3648,G3649,G3650,G3651);
  nand GNAME6787(G6787,G59105,G3185);
  nand GNAME6788(G6788,G59097,G3163);
  nand GNAME6789(G6789,G59089,G3166);
  nand GNAME6790(G6790,G59081,G3168);
  nand GNAME6791(G6791,G59073,G3171);
  nand GNAME6792(G6792,G59065,G3172);
  nand GNAME6793(G6793,G59057,G3173);
  nand GNAME6794(G6794,G59049,G3174);
  nand GNAME6795(G6795,G59041,G3176);
  nand GNAME6796(G6796,G59033,G3177);
  nand GNAME6797(G6797,G59025,G3178);
  nand GNAME6798(G6798,G59017,G3179);
  nand GNAME6799(G6799,G59009,G3181);
  nand GNAME6800(G6800,G59001,G3182);
  nand GNAME6801(G6801,G58993,G3183);
  nand GNAME6802(G6802,G58985,G3184);
  nand GNAME6803(G6803,G3652,G3653,G3654,G3655);
  nand GNAME6804(G6804,G59106,G3185);
  nand GNAME6805(G6805,G59098,G3163);
  nand GNAME6806(G6806,G59090,G3166);
  nand GNAME6807(G6807,G59082,G3168);
  nand GNAME6808(G6808,G59074,G3171);
  nand GNAME6809(G6809,G59066,G3172);
  nand GNAME6810(G6810,G59058,G3173);
  nand GNAME6811(G6811,G59050,G3174);
  nand GNAME6812(G6812,G59042,G3176);
  nand GNAME6813(G6813,G59034,G3177);
  nand GNAME6814(G6814,G59026,G3178);
  nand GNAME6815(G6815,G59018,G3179);
  nand GNAME6816(G6816,G59010,G3181);
  nand GNAME6817(G6817,G59002,G3182);
  nand GNAME6818(G6818,G58994,G3183);
  nand GNAME6819(G6819,G58986,G3184);
  nand GNAME6820(G6820,G3656,G3657,G3658,G3659);
  nand GNAME6821(G6821,G59107,G3185);
  nand GNAME6822(G6822,G59099,G3163);
  nand GNAME6823(G6823,G59091,G3166);
  nand GNAME6824(G6824,G59083,G3168);
  nand GNAME6825(G6825,G59075,G3171);
  nand GNAME6826(G6826,G59067,G3172);
  nand GNAME6827(G6827,G59059,G3173);
  nand GNAME6828(G6828,G59051,G3174);
  nand GNAME6829(G6829,G59043,G3176);
  nand GNAME6830(G6830,G59035,G3177);
  nand GNAME6831(G6831,G59027,G3178);
  nand GNAME6832(G6832,G59019,G3179);
  nand GNAME6833(G6833,G59011,G3181);
  nand GNAME6834(G6834,G59003,G3182);
  nand GNAME6835(G6835,G58995,G3183);
  nand GNAME6836(G6836,G58987,G3184);
  nand GNAME6837(G6837,G3660,G3661,G3662,G3663);
  nand GNAME6838(G6838,G3808,G3785,G3794);
  or GNAME6839(G6839,G3239,G3240);
  nand GNAME6840(G6840,G2827,G21265);
  nand GNAME6841(G6841,G6839,G20481);
  nand GNAME6842(G6842,G6838,G59127);
  nand GNAME6843(G6843,G20219,G3187);
  nand GNAME6844(G6844,G59318,G3189);
  nand GNAME6845(G6845,G2827,G21266);
  nand GNAME6846(G6846,G6839,G20516);
  nand GNAME6847(G6847,G6838,G59126);
  nand GNAME6848(G6848,G20176,G3187);
  nand GNAME6849(G6849,G59317,G3189);
  nand GNAME6850(G6850,G2827,G20506);
  nand GNAME6851(G6851,G6839,G20506);
  nand GNAME6852(G6852,G6838,G59125);
  nand GNAME6853(G6853,G20177,G3187);
  nand GNAME6854(G6854,G59316,G3189);
  nand GNAME6855(G6855,G2827,G20448);
  nand GNAME6856(G6856,G6839,G20448);
  nand GNAME6857(G6857,G6838,G59124);
  nand GNAME6858(G6858,G20143,G3187);
  nand GNAME6859(G6859,G59315,G3189);
  nand GNAME6860(G6860,G2827,G20520);
  nand GNAME6861(G6861,G6839,G20520);
  nand GNAME6862(G6862,G6838,G59123);
  nand GNAME6863(G6863,G20178,G3187);
  nand GNAME6864(G6864,G59314,G3189);
  nand GNAME6865(G6865,G2827,G20523);
  nand GNAME6866(G6866,G6839,G20523);
  nand GNAME6867(G6867,G6838,G59122);
  nand GNAME6868(G6868,G20179,G3187);
  nand GNAME6869(G6869,G59313,G3189);
  nand GNAME6870(G6870,G6839,G20508);
  nand GNAME6871(G6871,G6838,G59149);
  nand GNAME6872(G6872,G20210,G3187);
  nand GNAME6873(G6873,G59340,G3189);
  nand GNAME6874(G6874,G2827,G21267);
  nand GNAME6875(G6875,G6839,G20447);
  nand GNAME6876(G6876,G6838,G59148);
  nand GNAME6877(G6877,G20142,G3187);
  nand GNAME6878(G6878,G59339,G3189);
  nand GNAME6879(G6879,G2827,G20507);
  nand GNAME6880(G6880,G6839,G20507);
  nand GNAME6881(G6881,G6838,G59121);
  nand GNAME6882(G6882,G59312,G3189);
  nand GNAME6883(G6883,G20180,G3187);
  nand GNAME6884(G6884,G2827,G21268);
  nand GNAME6885(G6885,G6839,G20495);
  nand GNAME6886(G6886,G6838,G59147);
  nand GNAME6887(G6887,G20196,G3187);
  nand GNAME6888(G6888,G59338,G3189);
  nand GNAME6889(G6889,G2827,G21269);
  nand GNAME6890(G6890,G6839,G20496);
  nand GNAME6891(G6891,G6838,G59146);
  nand GNAME6892(G6892,G20197,G3187);
  nand GNAME6893(G6893,G59337,G3189);
  nand GNAME6894(G6894,G2827,G21270);
  nand GNAME6895(G6895,G6839,G20497);
  nand GNAME6896(G6896,G6838,G59145);
  nand GNAME6897(G6897,G20198,G3187);
  nand GNAME6898(G6898,G59336,G3189);
  nand GNAME6899(G6899,G2827,G21271);
  nand GNAME6900(G6900,G6839,G20498);
  nand GNAME6901(G6901,G6838,G59144);
  nand GNAME6902(G6902,G20199,G3187);
  nand GNAME6903(G6903,G59335,G3189);
  nand GNAME6904(G6904,G2827,G21272);
  nand GNAME6905(G6905,G6839,G20499);
  nand GNAME6906(G6906,G6838,G59143);
  nand GNAME6907(G6907,G20200,G3187);
  nand GNAME6908(G6908,G59334,G3189);
  nand GNAME6909(G6909,G2827,G21273);
  nand GNAME6910(G6910,G6839,G20537);
  nand GNAME6911(G6911,G6838,G59142);
  nand GNAME6912(G6912,G20201,G3187);
  nand GNAME6913(G6913,G59333,G3189);
  nand GNAME6914(G6914,G2827,G21274);
  nand GNAME6915(G6915,G6839,G20540);
  nand GNAME6916(G6916,G6838,G59141);
  nand GNAME6917(G6917,G20202,G3187);
  nand GNAME6918(G6918,G59332,G3189);
  nand GNAME6919(G6919,G2827,G21275);
  nand GNAME6920(G6920,G6839,G20543);
  nand GNAME6921(G6921,G6838,G59140);
  nand GNAME6922(G6922,G20203,G3187);
  nand GNAME6923(G6923,G59331,G3189);
  nand GNAME6924(G6924,G2827,G21276);
  nand GNAME6925(G6925,G6839,G20546);
  nand GNAME6926(G6926,G6838,G59139);
  nand GNAME6927(G6927,G20204,G3187);
  nand GNAME6928(G6928,G59330,G3189);
  nand GNAME6929(G6929,G2827,G21277);
  nand GNAME6930(G6930,G6839,G20549);
  nand GNAME6931(G6931,G6838,G59138);
  nand GNAME6932(G6932,G20205,G3187);
  nand GNAME6933(G6933,G59329,G3189);
  nand GNAME6934(G6934,G2827,G20446);
  nand GNAME6935(G6935,G6839,G20446);
  nand GNAME6936(G6936,G6838,G59120);
  nand GNAME6937(G6937,G59311,G3189);
  nand GNAME6938(G6938,G20141,G3187);
  nand GNAME6939(G6939,G2827,G21278);
  nand GNAME6940(G6940,G6839,G20555);
  nand GNAME6941(G6941,G6838,G59137);
  nand GNAME6942(G6942,G20206,G3187);
  nand GNAME6943(G6943,G59328,G3189);
  nand GNAME6944(G6944,G2827,G21279);
  nand GNAME6945(G6945,G6839,G20558);
  nand GNAME6946(G6946,G6838,G59136);
  nand GNAME6947(G6947,G20207,G3187);
  nand GNAME6948(G6948,G59327,G3189);
  nand GNAME6949(G6949,G2827,G21280);
  nand GNAME6950(G6950,G6839,G20561);
  nand GNAME6951(G6951,G6838,G59135);
  nand GNAME6952(G6952,G20208,G3187);
  nand GNAME6953(G6953,G59326,G3189);
  nand GNAME6954(G6954,G2827,G21293);
  nand GNAME6955(G6955,G6839,G20500);
  nand GNAME6956(G6956,G6838,G59134);
  nand GNAME6957(G6957,G20236,G3187);
  nand GNAME6958(G6958,G59325,G3189);
  nand GNAME6959(G6959,G2827,G21230);
  nand GNAME6960(G6960,G6839,G20501);
  nand GNAME6961(G6961,G6838,G59133);
  nand GNAME6962(G6962,G20239,G3187);
  nand GNAME6963(G6963,G59324,G3189);
  nand GNAME6964(G6964,G2827,G21295);
  nand GNAME6965(G6965,G6839,G20445);
  nand GNAME6966(G6966,G6838,G59132);
  nand GNAME6967(G6967,G20211,G3187);
  nand GNAME6968(G6968,G59323,G3189);
  nand GNAME6969(G6969,G2827,G21296);
  nand GNAME6970(G6970,G6839,G20502);
  nand GNAME6971(G6971,G6838,G59131);
  nand GNAME6972(G6972,G20243,G3187);
  nand GNAME6973(G6973,G59322,G3189);
  nand GNAME6974(G6974,G2827,G21297);
  nand GNAME6975(G6975,G6839,G20503);
  nand GNAME6976(G6976,G6838,G59130);
  nand GNAME6977(G6977,G20246,G3187);
  nand GNAME6978(G6978,G59321,G3189);
  nand GNAME6979(G6979,G2827,G21298);
  nand GNAME6980(G6980,G6839,G20504);
  nand GNAME6981(G6981,G6838,G59129);
  nand GNAME6982(G6982,G20212,G3187);
  nand GNAME6983(G6983,G59320,G3189);
  nand GNAME6984(G6984,G2827,G21299);
  nand GNAME6985(G6985,G6839,G20444);
  nand GNAME6986(G6986,G6838,G59128);
  nand GNAME6987(G6987,G20140,G3187);
  nand GNAME6988(G6988,G59319,G3189);
  nand GNAME6989(G6989,G2827,G20552);
  nand GNAME6990(G6990,G6839,G20552);
  nand GNAME6991(G6991,G6838,G59119);
  nand GNAME6992(G6992,G20233,G3187);
  nand GNAME6993(G6993,G59310,G3189);
  nand GNAME6994(G6994,G2827,G20505);
  nand GNAME6995(G6995,G6839,G20505);
  nand GNAME6996(G6996,G6838,G59118);
  nand GNAME6997(G6997,G20209,G3187);
  nand GNAME6998(G6998,G59309,G3189);
  nand GNAME6999(G6999,G59092,G5271);
  nand GNAME7000(G7000,G59084,G5332);
  nand GNAME7001(G7001,G59076,G5393);
  nand GNAME7002(G7002,G59068,G5454);
  nand GNAME7003(G7003,G59060,G5515);
  nand GNAME7004(G7004,G59052,G5576);
  nand GNAME7005(G7005,G59044,G5637);
  nand GNAME7006(G7006,G59036,G5698);
  nand GNAME7007(G7007,G59028,G5759);
  nand GNAME7008(G7008,G59020,G5820);
  nand GNAME7009(G7009,G59012,G5881);
  nand GNAME7010(G7010,G59004,G5942);
  nand GNAME7011(G7011,G58996,G6003);
  nand GNAME7012(G7012,G58988,G6064);
  nand GNAME7013(G7013,G58980,G6125);
  nand GNAME7014(G7014,G59100,G5189);
  nand GNAME7015(G7015,G3673,G3674,G3675,G3676);
  nand GNAME7016(G7016,G59092,G3217);
  nand GNAME7017(G7017,G59084,G3219);
  nand GNAME7018(G7018,G59076,G3221);
  nand GNAME7019(G7019,G59068,G3224);
  nand GNAME7020(G7020,G59060,G3225);
  nand GNAME7021(G7021,G59052,G3226);
  nand GNAME7022(G7022,G59044,G3227);
  nand GNAME7023(G7023,G59036,G3229);
  nand GNAME7024(G7024,G59028,G3230);
  nand GNAME7025(G7025,G59020,G3231);
  nand GNAME7026(G7026,G59012,G3232);
  nand GNAME7027(G7027,G59004,G3234);
  nand GNAME7028(G7028,G58996,G3235);
  nand GNAME7029(G7029,G58988,G3236);
  nand GNAME7030(G7030,G58980,G3237);
  nand GNAME7031(G7031,G59100,G3238);
  nand GNAME7032(G7032,G3669,G3670,G3671,G3672);
  nand GNAME7033(G7033,G59092,G3193);
  nand GNAME7034(G7034,G59084,G3196);
  nand GNAME7035(G7035,G59076,G3197);
  nand GNAME7036(G7036,G59068,G3199);
  nand GNAME7037(G7037,G59060,G3201);
  nand GNAME7038(G7038,G59052,G3202);
  nand GNAME7039(G7039,G59044,G3203);
  nand GNAME7040(G7040,G59036,G3205);
  nand GNAME7041(G7041,G59028,G3206);
  nand GNAME7042(G7042,G59020,G3208);
  nand GNAME7043(G7043,G59012,G3209);
  nand GNAME7044(G7044,G59004,G3210);
  nand GNAME7045(G7045,G58996,G3211);
  nand GNAME7046(G7046,G58988,G3212);
  nand GNAME7047(G7047,G58980,G3213);
  nand GNAME7048(G7048,G59100,G3214);
  nand GNAME7049(G7049,G3665,G3666,G3667,G3668);
  nand GNAME7050(G7050,G3187,G20438);
  nand GNAME7051(G7051,G7049,G2827);
  nand GNAME7052(G7052,G7032,G3239);
  nand GNAME7053(G7053,G7015,G3240);
  nand GNAME7054(G7054,G59093,G5271);
  nand GNAME7055(G7055,G59085,G5332);
  nand GNAME7056(G7056,G59077,G5393);
  nand GNAME7057(G7057,G59069,G5454);
  nand GNAME7058(G7058,G59061,G5515);
  nand GNAME7059(G7059,G59053,G5576);
  nand GNAME7060(G7060,G59045,G5637);
  nand GNAME7061(G7061,G59037,G5698);
  nand GNAME7062(G7062,G59029,G5759);
  nand GNAME7063(G7063,G59021,G5820);
  nand GNAME7064(G7064,G59013,G5881);
  nand GNAME7065(G7065,G59005,G5942);
  nand GNAME7066(G7066,G58997,G6003);
  nand GNAME7067(G7067,G58989,G6064);
  nand GNAME7068(G7068,G58981,G6125);
  nand GNAME7069(G7069,G59101,G5189);
  nand GNAME7070(G7070,G3685,G3686,G3687,G3688);
  nand GNAME7071(G7071,G59093,G3217);
  nand GNAME7072(G7072,G59085,G3219);
  nand GNAME7073(G7073,G59077,G3221);
  nand GNAME7074(G7074,G59069,G3224);
  nand GNAME7075(G7075,G59061,G3225);
  nand GNAME7076(G7076,G59053,G3226);
  nand GNAME7077(G7077,G59045,G3227);
  nand GNAME7078(G7078,G59037,G3229);
  nand GNAME7079(G7079,G59029,G3230);
  nand GNAME7080(G7080,G59021,G3231);
  nand GNAME7081(G7081,G59013,G3232);
  nand GNAME7082(G7082,G59005,G3234);
  nand GNAME7083(G7083,G58997,G3235);
  nand GNAME7084(G7084,G58989,G3236);
  nand GNAME7085(G7085,G58981,G3237);
  nand GNAME7086(G7086,G59101,G3238);
  nand GNAME7087(G7087,G3681,G3682,G3683,G3684);
  nand GNAME7088(G7088,G59093,G3193);
  nand GNAME7089(G7089,G59085,G3196);
  nand GNAME7090(G7090,G59077,G3197);
  nand GNAME7091(G7091,G59069,G3199);
  nand GNAME7092(G7092,G59061,G3201);
  nand GNAME7093(G7093,G59053,G3202);
  nand GNAME7094(G7094,G59045,G3203);
  nand GNAME7095(G7095,G59037,G3205);
  nand GNAME7096(G7096,G59029,G3206);
  nand GNAME7097(G7097,G59021,G3208);
  nand GNAME7098(G7098,G59013,G3209);
  nand GNAME7099(G7099,G59005,G3210);
  nand GNAME7100(G7100,G58997,G3211);
  nand GNAME7101(G7101,G58989,G3212);
  nand GNAME7102(G7102,G58981,G3213);
  nand GNAME7103(G7103,G59101,G3214);
  nand GNAME7104(G7104,G3677,G3678,G3679,G3680);
  nand GNAME7105(G7105,G3187,G20436);
  nand GNAME7106(G7106,G7104,G2827);
  nand GNAME7107(G7107,G7087,G3239);
  nand GNAME7108(G7108,G7070,G3240);
  nand GNAME7109(G7109,G59094,G5271);
  nand GNAME7110(G7110,G59086,G5332);
  nand GNAME7111(G7111,G59078,G5393);
  nand GNAME7112(G7112,G59070,G5454);
  nand GNAME7113(G7113,G59062,G5515);
  nand GNAME7114(G7114,G59054,G5576);
  nand GNAME7115(G7115,G59046,G5637);
  nand GNAME7116(G7116,G59038,G5698);
  nand GNAME7117(G7117,G59030,G5759);
  nand GNAME7118(G7118,G59022,G5820);
  nand GNAME7119(G7119,G59014,G5881);
  nand GNAME7120(G7120,G59006,G5942);
  nand GNAME7121(G7121,G58998,G6003);
  nand GNAME7122(G7122,G58990,G6064);
  nand GNAME7123(G7123,G58982,G6125);
  nand GNAME7124(G7124,G59102,G5189);
  nand GNAME7125(G7125,G3697,G3698,G3699,G3700);
  nand GNAME7126(G7126,G59094,G3217);
  nand GNAME7127(G7127,G59086,G3219);
  nand GNAME7128(G7128,G59078,G3221);
  nand GNAME7129(G7129,G59070,G3224);
  nand GNAME7130(G7130,G59062,G3225);
  nand GNAME7131(G7131,G59054,G3226);
  nand GNAME7132(G7132,G59046,G3227);
  nand GNAME7133(G7133,G59038,G3229);
  nand GNAME7134(G7134,G59030,G3230);
  nand GNAME7135(G7135,G59022,G3231);
  nand GNAME7136(G7136,G59014,G3232);
  nand GNAME7137(G7137,G59006,G3234);
  nand GNAME7138(G7138,G58998,G3235);
  nand GNAME7139(G7139,G58990,G3236);
  nand GNAME7140(G7140,G58982,G3237);
  nand GNAME7141(G7141,G59102,G3238);
  nand GNAME7142(G7142,G3693,G3694,G3695,G3696);
  nand GNAME7143(G7143,G59094,G3193);
  nand GNAME7144(G7144,G59086,G3196);
  nand GNAME7145(G7145,G59078,G3197);
  nand GNAME7146(G7146,G59070,G3199);
  nand GNAME7147(G7147,G59062,G3201);
  nand GNAME7148(G7148,G59054,G3202);
  nand GNAME7149(G7149,G59046,G3203);
  nand GNAME7150(G7150,G59038,G3205);
  nand GNAME7151(G7151,G59030,G3206);
  nand GNAME7152(G7152,G59022,G3208);
  nand GNAME7153(G7153,G59014,G3209);
  nand GNAME7154(G7154,G59006,G3210);
  nand GNAME7155(G7155,G58998,G3211);
  nand GNAME7156(G7156,G58990,G3212);
  nand GNAME7157(G7157,G58982,G3213);
  nand GNAME7158(G7158,G59102,G3214);
  nand GNAME7159(G7159,G3689,G3690,G3691,G3692);
  nand GNAME7160(G7160,G3187,G20439);
  nand GNAME7161(G7161,G7159,G2827);
  nand GNAME7162(G7162,G7142,G3239);
  nand GNAME7163(G7163,G7125,G3240);
  nand GNAME7164(G7164,G59095,G3217);
  nand GNAME7165(G7165,G59087,G3219);
  nand GNAME7166(G7166,G59079,G3221);
  nand GNAME7167(G7167,G59071,G3224);
  nand GNAME7168(G7168,G59063,G3225);
  nand GNAME7169(G7169,G59055,G3226);
  nand GNAME7170(G7170,G59047,G3227);
  nand GNAME7171(G7171,G59039,G3229);
  nand GNAME7172(G7172,G59031,G3230);
  nand GNAME7173(G7173,G59023,G3231);
  nand GNAME7174(G7174,G59015,G3232);
  nand GNAME7175(G7175,G59007,G3234);
  nand GNAME7176(G7176,G58999,G3235);
  nand GNAME7177(G7177,G58991,G3236);
  nand GNAME7178(G7178,G58983,G3237);
  nand GNAME7179(G7179,G59103,G3238);
  nand GNAME7180(G7180,G3709,G3710,G3711,G3712);
  nand GNAME7181(G7181,G59095,G3193);
  nand GNAME7182(G7182,G59087,G3196);
  nand GNAME7183(G7183,G59079,G3197);
  nand GNAME7184(G7184,G59071,G3199);
  nand GNAME7185(G7185,G59063,G3201);
  nand GNAME7186(G7186,G59055,G3202);
  nand GNAME7187(G7187,G59047,G3203);
  nand GNAME7188(G7188,G59039,G3205);
  nand GNAME7189(G7189,G59031,G3206);
  nand GNAME7190(G7190,G59023,G3208);
  nand GNAME7191(G7191,G59015,G3209);
  nand GNAME7192(G7192,G59007,G3210);
  nand GNAME7193(G7193,G58999,G3211);
  nand GNAME7194(G7194,G58991,G3212);
  nand GNAME7195(G7195,G58983,G3213);
  nand GNAME7196(G7196,G59103,G3214);
  nand GNAME7197(G7197,G3705,G3706,G3707,G3708);
  nand GNAME7198(G7198,G59095,G5271);
  nand GNAME7199(G7199,G59087,G5332);
  nand GNAME7200(G7200,G59079,G5393);
  nand GNAME7201(G7201,G59071,G5454);
  nand GNAME7202(G7202,G59063,G5515);
  nand GNAME7203(G7203,G59055,G5576);
  nand GNAME7204(G7204,G59047,G5637);
  nand GNAME7205(G7205,G59039,G5698);
  nand GNAME7206(G7206,G59031,G5759);
  nand GNAME7207(G7207,G59023,G5820);
  nand GNAME7208(G7208,G59015,G5881);
  nand GNAME7209(G7209,G59007,G5942);
  nand GNAME7210(G7210,G58999,G6003);
  nand GNAME7211(G7211,G58991,G6064);
  nand GNAME7212(G7212,G58983,G6125);
  nand GNAME7213(G7213,G59103,G5189);
  nand GNAME7214(G7214,G3701,G3702,G3703,G3704);
  or GNAME7215(G7215,G3886,G7985);
  nand GNAME7216(G7216,G3187,G20443);
  nand GNAME7217(G7217,G7214,G3240);
  nand GNAME7218(G7218,G7197,G2827);
  nand GNAME7219(G7219,G7180,G3239);
  nand GNAME7220(G7220,G59096,G3217);
  nand GNAME7221(G7221,G59088,G3219);
  nand GNAME7222(G7222,G59080,G3221);
  nand GNAME7223(G7223,G59072,G3224);
  nand GNAME7224(G7224,G59064,G3225);
  nand GNAME7225(G7225,G59056,G3226);
  nand GNAME7226(G7226,G59048,G3227);
  nand GNAME7227(G7227,G59040,G3229);
  nand GNAME7228(G7228,G59032,G3230);
  nand GNAME7229(G7229,G59024,G3231);
  nand GNAME7230(G7230,G59016,G3232);
  nand GNAME7231(G7231,G59008,G3234);
  nand GNAME7232(G7232,G59000,G3235);
  nand GNAME7233(G7233,G58992,G3236);
  nand GNAME7234(G7234,G58984,G3237);
  nand GNAME7235(G7235,G59104,G3238);
  nand GNAME7236(G7236,G3721,G3722,G3723,G3724);
  nand GNAME7237(G7237,G59096,G3193);
  nand GNAME7238(G7238,G59088,G3196);
  nand GNAME7239(G7239,G59080,G3197);
  nand GNAME7240(G7240,G59072,G3199);
  nand GNAME7241(G7241,G59064,G3201);
  nand GNAME7242(G7242,G59056,G3202);
  nand GNAME7243(G7243,G59048,G3203);
  nand GNAME7244(G7244,G59040,G3205);
  nand GNAME7245(G7245,G59032,G3206);
  nand GNAME7246(G7246,G59024,G3208);
  nand GNAME7247(G7247,G59016,G3209);
  nand GNAME7248(G7248,G59008,G3210);
  nand GNAME7249(G7249,G59000,G3211);
  nand GNAME7250(G7250,G58992,G3212);
  nand GNAME7251(G7251,G58984,G3213);
  nand GNAME7252(G7252,G59104,G3214);
  nand GNAME7253(G7253,G3717,G3718,G3719,G3720);
  nand GNAME7254(G7254,G59096,G5271);
  nand GNAME7255(G7255,G59088,G5332);
  nand GNAME7256(G7256,G59080,G5393);
  nand GNAME7257(G7257,G59072,G5454);
  nand GNAME7258(G7258,G59064,G5515);
  nand GNAME7259(G7259,G59056,G5576);
  nand GNAME7260(G7260,G59048,G5637);
  nand GNAME7261(G7261,G59040,G5698);
  nand GNAME7262(G7262,G59032,G5759);
  nand GNAME7263(G7263,G59024,G5820);
  nand GNAME7264(G7264,G59016,G5881);
  nand GNAME7265(G7265,G59008,G5942);
  nand GNAME7266(G7266,G59000,G6003);
  nand GNAME7267(G7267,G58992,G6064);
  nand GNAME7268(G7268,G58984,G6125);
  nand GNAME7269(G7269,G59104,G5189);
  nand GNAME7270(G7270,G3713,G3714,G3715,G3716);
  nand GNAME7271(G7271,G3187,G20441);
  nand GNAME7272(G7272,G7270,G3240);
  nand GNAME7273(G7273,G7253,G2827);
  nand GNAME7274(G7274,G7236,G3239);
  nand GNAME7275(G7275,G2784,G59109);
  nand GNAME7276(G7276,G59105,G3238);
  nand GNAME7277(G7277,G59097,G3217);
  nand GNAME7278(G7278,G59089,G3219);
  nand GNAME7279(G7279,G59081,G3221);
  nand GNAME7280(G7280,G59073,G3224);
  nand GNAME7281(G7281,G59065,G3225);
  nand GNAME7282(G7282,G59057,G3226);
  nand GNAME7283(G7283,G59049,G3227);
  nand GNAME7284(G7284,G59041,G3229);
  nand GNAME7285(G7285,G59033,G3230);
  nand GNAME7286(G7286,G59025,G3231);
  nand GNAME7287(G7287,G59017,G3232);
  nand GNAME7288(G7288,G59009,G3234);
  nand GNAME7289(G7289,G59001,G3235);
  nand GNAME7290(G7290,G58993,G3236);
  nand GNAME7291(G7291,G58985,G3237);
  nand GNAME7292(G7292,G3733,G3734,G3735,G3736);
  nand GNAME7293(G7293,G59105,G3214);
  nand GNAME7294(G7294,G59097,G3193);
  nand GNAME7295(G7295,G59089,G3196);
  nand GNAME7296(G7296,G59081,G3197);
  nand GNAME7297(G7297,G59073,G3199);
  nand GNAME7298(G7298,G59065,G3201);
  nand GNAME7299(G7299,G59057,G3202);
  nand GNAME7300(G7300,G59049,G3203);
  nand GNAME7301(G7301,G59041,G3205);
  nand GNAME7302(G7302,G59033,G3206);
  nand GNAME7303(G7303,G59025,G3208);
  nand GNAME7304(G7304,G59017,G3209);
  nand GNAME7305(G7305,G59009,G3210);
  nand GNAME7306(G7306,G59001,G3211);
  nand GNAME7307(G7307,G58993,G3212);
  nand GNAME7308(G7308,G58985,G3213);
  nand GNAME7309(G7309,G3729,G3730,G3731,G3732);
  nand GNAME7310(G7310,G59105,G5189);
  nand GNAME7311(G7311,G59097,G5271);
  nand GNAME7312(G7312,G59089,G5332);
  nand GNAME7313(G7313,G59081,G5393);
  nand GNAME7314(G7314,G59073,G5454);
  nand GNAME7315(G7315,G59065,G5515);
  nand GNAME7316(G7316,G59057,G5576);
  nand GNAME7317(G7317,G59049,G5637);
  nand GNAME7318(G7318,G59041,G5698);
  nand GNAME7319(G7319,G59033,G5759);
  nand GNAME7320(G7320,G59025,G5820);
  nand GNAME7321(G7321,G59017,G5881);
  nand GNAME7322(G7322,G59009,G5942);
  nand GNAME7323(G7323,G59001,G6003);
  nand GNAME7324(G7324,G58993,G6064);
  nand GNAME7325(G7325,G58985,G6125);
  nand GNAME7326(G7326,G3725,G3726,G3727,G3728);
  nand GNAME7327(G7327,G3187,G20442);
  nand GNAME7328(G7328,G7326,G3240);
  nand GNAME7329(G7329,G7309,G2827);
  nand GNAME7330(G7330,G7292,G3239);
  nand GNAME7331(G7331,G2784,G59110);
  nand GNAME7332(G7332,G59106,G3238);
  nand GNAME7333(G7333,G59098,G3217);
  nand GNAME7334(G7334,G59090,G3219);
  nand GNAME7335(G7335,G59082,G3221);
  nand GNAME7336(G7336,G59074,G3224);
  nand GNAME7337(G7337,G59066,G3225);
  nand GNAME7338(G7338,G59058,G3226);
  nand GNAME7339(G7339,G59050,G3227);
  nand GNAME7340(G7340,G59042,G3229);
  nand GNAME7341(G7341,G59034,G3230);
  nand GNAME7342(G7342,G59026,G3231);
  nand GNAME7343(G7343,G59018,G3232);
  nand GNAME7344(G7344,G59010,G3234);
  nand GNAME7345(G7345,G59002,G3235);
  nand GNAME7346(G7346,G58994,G3236);
  nand GNAME7347(G7347,G58986,G3237);
  nand GNAME7348(G7348,G3746,G3747,G3748,G3749);
  nand GNAME7349(G7349,G59106,G3214);
  nand GNAME7350(G7350,G59098,G3193);
  nand GNAME7351(G7351,G59090,G3196);
  nand GNAME7352(G7352,G59082,G3197);
  nand GNAME7353(G7353,G59074,G3199);
  nand GNAME7354(G7354,G59066,G3201);
  nand GNAME7355(G7355,G59058,G3202);
  nand GNAME7356(G7356,G59050,G3203);
  nand GNAME7357(G7357,G59042,G3205);
  nand GNAME7358(G7358,G59034,G3206);
  nand GNAME7359(G7359,G59026,G3208);
  nand GNAME7360(G7360,G59018,G3209);
  nand GNAME7361(G7361,G59010,G3210);
  nand GNAME7362(G7362,G59002,G3211);
  nand GNAME7363(G7363,G58994,G3212);
  nand GNAME7364(G7364,G58986,G3213);
  nand GNAME7365(G7365,G3742,G3743,G3744,G3745);
  nand GNAME7366(G7366,G59106,G5189);
  nand GNAME7367(G7367,G59098,G5271);
  nand GNAME7368(G7368,G59090,G5332);
  nand GNAME7369(G7369,G59082,G5393);
  nand GNAME7370(G7370,G59074,G5454);
  nand GNAME7371(G7371,G59066,G5515);
  nand GNAME7372(G7372,G59058,G5576);
  nand GNAME7373(G7373,G59050,G5637);
  nand GNAME7374(G7374,G59042,G5698);
  nand GNAME7375(G7375,G59034,G5759);
  nand GNAME7376(G7376,G59026,G5820);
  nand GNAME7377(G7377,G59018,G5881);
  nand GNAME7378(G7378,G59010,G5942);
  nand GNAME7379(G7379,G59002,G6003);
  nand GNAME7380(G7380,G58994,G6064);
  nand GNAME7381(G7381,G58986,G6125);
  nand GNAME7382(G7382,G3738,G3739,G3740,G3741);
  nand GNAME7383(G7383,G3187,G20437);
  nand GNAME7384(G7384,G7382,G3240);
  nand GNAME7385(G7385,G7365,G2827);
  nand GNAME7386(G7386,G7348,G3239);
  nand GNAME7387(G7387,G2784,G59111);
  nand GNAME7388(G7388,G59107,G3238);
  nand GNAME7389(G7389,G59099,G3217);
  nand GNAME7390(G7390,G59091,G3219);
  nand GNAME7391(G7391,G59083,G3221);
  nand GNAME7392(G7392,G59075,G3224);
  nand GNAME7393(G7393,G59067,G3225);
  nand GNAME7394(G7394,G59059,G3226);
  nand GNAME7395(G7395,G59051,G3227);
  nand GNAME7396(G7396,G59043,G3229);
  nand GNAME7397(G7397,G59035,G3230);
  nand GNAME7398(G7398,G59027,G3231);
  nand GNAME7399(G7399,G59019,G3232);
  nand GNAME7400(G7400,G59011,G3234);
  nand GNAME7401(G7401,G59003,G3235);
  nand GNAME7402(G7402,G58995,G3236);
  nand GNAME7403(G7403,G58987,G3237);
  nand GNAME7404(G7404,G3759,G3760,G3761,G3762);
  nand GNAME7405(G7405,G59107,G3214);
  nand GNAME7406(G7406,G59099,G3193);
  nand GNAME7407(G7407,G59091,G3196);
  nand GNAME7408(G7408,G59083,G3197);
  nand GNAME7409(G7409,G59075,G3199);
  nand GNAME7410(G7410,G59067,G3201);
  nand GNAME7411(G7411,G59059,G3202);
  nand GNAME7412(G7412,G59051,G3203);
  nand GNAME7413(G7413,G59043,G3205);
  nand GNAME7414(G7414,G59035,G3206);
  nand GNAME7415(G7415,G59027,G3208);
  nand GNAME7416(G7416,G59019,G3209);
  nand GNAME7417(G7417,G59011,G3210);
  nand GNAME7418(G7418,G59003,G3211);
  nand GNAME7419(G7419,G58995,G3212);
  nand GNAME7420(G7420,G58987,G3213);
  nand GNAME7421(G7421,G3755,G3756,G3757,G3758);
  nand GNAME7422(G7422,G59107,G5189);
  nand GNAME7423(G7423,G59099,G5271);
  nand GNAME7424(G7424,G59091,G5332);
  nand GNAME7425(G7425,G59083,G5393);
  nand GNAME7426(G7426,G59075,G5454);
  nand GNAME7427(G7427,G59067,G5515);
  nand GNAME7428(G7428,G59059,G5576);
  nand GNAME7429(G7429,G59051,G5637);
  nand GNAME7430(G7430,G59043,G5698);
  nand GNAME7431(G7431,G59035,G5759);
  nand GNAME7432(G7432,G59027,G5820);
  nand GNAME7433(G7433,G59019,G5881);
  nand GNAME7434(G7434,G59011,G5942);
  nand GNAME7435(G7435,G59003,G6003);
  nand GNAME7436(G7436,G58995,G6064);
  nand GNAME7437(G7437,G58987,G6125);
  nand GNAME7438(G7438,G3751,G3752,G3753,G3754);
  nand GNAME7439(G7439,G3187,G20440);
  nand GNAME7440(G7440,G7438,G3240);
  nand GNAME7441(G7441,G7421,G2827);
  nand GNAME7442(G7442,G7404,G3239);
  nand GNAME7443(G7443,G2784,G59112);
  nand GNAME7444(G7444,G2801,G3240,G58979,G2785,G3903);
  nand GNAME7445(G7445,G59105,G2859);
  or GNAME7446(G7446,G2790,G3920,G2753);
  nand GNAME7447(G7447,G2787,G58979,G2801,G7990);
  nand GNAME7448(G7448,G59106,G2859);
  nand GNAME7449(G7449,G2784,G3835);
  nand GNAME7450(G7450,G2794,G2890);
  nand GNAME7451(G7451,G3765,G7835,G7970,G2895,G3243);
  nand GNAME7452(G7452,G7451,G58979);
  nand GNAME7453(G7453,G59107,G2859);
  nand GNAME7454(G7454,G2855,G2863);
  nand GNAME7455(G7455,G3852,G2856);
  nand GNAME7456(G7456,G2783,G3954);
  nand GNAME7457(G7457,G7456,G7454,G7455);
  nand GNAME7458(G7458,G2749,G2795);
  nand GNAME7459(G7459,G2746,G2785);
  nand GNAME7460(G7460,G7459,G3786);
  nand GNAME7461(G7461,G7460,G2890);
  nand GNAME7462(G7462,G7458,G2830);
  nand GNAME7463(G7463,G2856,G2897);
  nand GNAME7464(G7464,G2795,G7457);
  nand GNAME7465(G7465,G2824,G2827);
  nand GNAME7466(G7466,G3766,G2898,G7464,G7465);
  nand GNAME7467(G7467,G7466,G58979);
  or GNAME7468(G7468,G2902,G2790);
  nand GNAME7469(G7469,G3810,G7444,G7468,G3244);
  nand GNAME7470(G7470,G3799,G3782);
  nand GNAME7471(G7471,G7470,G20219);
  nand GNAME7472(G7472,G7469,G59127);
  nand GNAME7473(G7473,G3783,G59159);
  nand GNAME7474(G7474,G2791,G59318);
  nand GNAME7475(G7475,G7470,G20176);
  nand GNAME7476(G7476,G7469,G59126);
  nand GNAME7477(G7477,G3783,G59158);
  nand GNAME7478(G7478,G2791,G59317);
  nand GNAME7479(G7479,G7470,G20177);
  nand GNAME7480(G7480,G7469,G59125);
  nand GNAME7481(G7481,G3783,G59157);
  nand GNAME7482(G7482,G2791,G59316);
  nand GNAME7483(G7483,G7470,G20143);
  nand GNAME7484(G7484,G7469,G59124);
  nand GNAME7485(G7485,G3783,G59156);
  nand GNAME7486(G7486,G2791,G59315);
  nand GNAME7487(G7487,G7470,G20178);
  nand GNAME7488(G7488,G7469,G59123);
  nand GNAME7489(G7489,G3783,G59155);
  nand GNAME7490(G7490,G2791,G59314);
  nand GNAME7491(G7491,G58979,G2874);
  nand GNAME7492(G7492,G7491,G2866);
  nand GNAME7493(G7493,G7492,G59108);
  nand GNAME7494(G7494,G7470,G20179);
  nand GNAME7495(G7495,G7469,G59122);
  nand GNAME7496(G7496,G3783,G59154);
  nand GNAME7497(G7497,G2791,G59313);
  nand GNAME7498(G7498,G7469,G59149);
  nand GNAME7499(G7499,G3783,G59181);
  nand GNAME7500(G7500,G2836,G20210);
  nand GNAME7501(G7501,G2791,G59340);
  nand GNAME7502(G7502,G7470,G20142);
  nand GNAME7503(G7503,G7469,G59148);
  nand GNAME7504(G7504,G3783,G59180);
  nand GNAME7505(G7505,G2791,G59339);
  nand GNAME7506(G7506,G6582,G2867);
  nand GNAME7507(G7507,G4833,G4834);
  nand GNAME7508(G7508,G7507,G58979);
  nand GNAME7509(G7509,G3186,G3241);
  or GNAME7510(G7510,G2905,G2790);
  nand GNAME7511(G7511,G7510,G3245,G7509,G3800,G4323);
  nand GNAME7512(G7512,G7511,G59109);
  nand GNAME7513(G7513,G7470,G20180);
  nand GNAME7514(G7514,G7469,G59121);
  nand GNAME7515(G7515,G3783,G59153);
  nand GNAME7516(G7516,G2791,G59312);
  nand GNAME7517(G7517,G7470,G20196);
  nand GNAME7518(G7518,G7469,G59147);
  nand GNAME7519(G7519,G3783,G59179);
  nand GNAME7520(G7520,G2791,G59338);
  nand GNAME7521(G7521,G6599,G2867);
  nand GNAME7522(G7522,G7470,G20197);
  nand GNAME7523(G7523,G7469,G59146);
  nand GNAME7524(G7524,G3783,G59178);
  nand GNAME7525(G7525,G2791,G59337);
  nand GNAME7526(G7526,G6616,G2867);
  nand GNAME7527(G7527,G7470,G20198);
  nand GNAME7528(G7528,G7469,G59145);
  nand GNAME7529(G7529,G3783,G59177);
  nand GNAME7530(G7530,G2791,G59336);
  nand GNAME7531(G7531,G6633,G2867);
  nand GNAME7532(G7532,G7470,G20199);
  nand GNAME7533(G7533,G7469,G59144);
  nand GNAME7534(G7534,G3783,G59176);
  nand GNAME7535(G7535,G2791,G59335);
  nand GNAME7536(G7536,G6650,G2867);
  nand GNAME7537(G7537,G7470,G20200);
  nand GNAME7538(G7538,G7469,G59143);
  nand GNAME7539(G7539,G3783,G59175);
  nand GNAME7540(G7540,G2791,G59334);
  nand GNAME7541(G7541,G6667,G2867);
  nand GNAME7542(G7542,G7470,G20201);
  nand GNAME7543(G7543,G7469,G59142);
  nand GNAME7544(G7544,G3783,G59174);
  nand GNAME7545(G7545,G2791,G59333);
  nand GNAME7546(G7546,G6684,G2867);
  nand GNAME7547(G7547,G7470,G20202);
  nand GNAME7548(G7548,G7469,G59141);
  nand GNAME7549(G7549,G3783,G59173);
  nand GNAME7550(G7550,G2791,G59332);
  nand GNAME7551(G7551,G6701,G2867);
  nand GNAME7552(G7552,G7470,G20203);
  nand GNAME7553(G7553,G7469,G59140);
  nand GNAME7554(G7554,G3783,G59172);
  nand GNAME7555(G7555,G2791,G59331);
  nand GNAME7556(G7556,G7470,G20204);
  nand GNAME7557(G7557,G7469,G59139);
  nand GNAME7558(G7558,G3783,G59171);
  nand GNAME7559(G7559,G2791,G59330);
  nand GNAME7560(G7560,G7470,G20205);
  nand GNAME7561(G7561,G7469,G59138);
  nand GNAME7562(G7562,G3783,G59170);
  nand GNAME7563(G7563,G2791,G59329);
  nand GNAME7564(G7564,G7511,G59110);
  nand GNAME7565(G7565,G7470,G20141);
  nand GNAME7566(G7566,G7469,G59120);
  nand GNAME7567(G7567,G3783,G59152);
  nand GNAME7568(G7568,G2791,G59311);
  nand GNAME7569(G7569,G7470,G20206);
  nand GNAME7570(G7570,G7469,G59137);
  nand GNAME7571(G7571,G3783,G59169);
  nand GNAME7572(G7572,G2791,G59328);
  nand GNAME7573(G7573,G7470,G20207);
  nand GNAME7574(G7574,G7469,G59136);
  nand GNAME7575(G7575,G3783,G59168);
  nand GNAME7576(G7576,G2791,G59327);
  nand GNAME7577(G7577,G7470,G20208);
  nand GNAME7578(G7578,G7469,G59135);
  nand GNAME7579(G7579,G3783,G59167);
  nand GNAME7580(G7580,G2791,G59326);
  nand GNAME7581(G7581,G7470,G20236);
  nand GNAME7582(G7582,G7469,G59134);
  nand GNAME7583(G7583,G3783,G59166);
  nand GNAME7584(G7584,G2791,G59325);
  nand GNAME7585(G7585,G7470,G20239);
  nand GNAME7586(G7586,G7469,G59133);
  nand GNAME7587(G7587,G3783,G59165);
  nand GNAME7588(G7588,G2791,G59324);
  nand GNAME7589(G7589,G7470,G20211);
  nand GNAME7590(G7590,G7469,G59132);
  nand GNAME7591(G7591,G3783,G59164);
  nand GNAME7592(G7592,G2791,G59323);
  nand GNAME7593(G7593,G7470,G20243);
  nand GNAME7594(G7594,G7469,G59131);
  nand GNAME7595(G7595,G3783,G59163);
  nand GNAME7596(G7596,G2791,G59322);
  nand GNAME7597(G7597,G7470,G20246);
  nand GNAME7598(G7598,G7469,G59130);
  nand GNAME7599(G7599,G3783,G59162);
  nand GNAME7600(G7600,G2791,G59321);
  nand GNAME7601(G7601,G7470,G20212);
  nand GNAME7602(G7602,G7469,G59129);
  nand GNAME7603(G7603,G3783,G59161);
  nand GNAME7604(G7604,G2791,G59320);
  nand GNAME7605(G7605,G7470,G20140);
  nand GNAME7606(G7606,G7469,G59128);
  nand GNAME7607(G7607,G3783,G59160);
  nand GNAME7608(G7608,G2791,G59319);
  nand GNAME7609(G7609,G7511,G59111);
  nand GNAME7610(G7610,G7470,G20233);
  nand GNAME7611(G7611,G7469,G59119);
  nand GNAME7612(G7612,G3783,G59151);
  nand GNAME7613(G7613,G2791,G59310);
  nand GNAME7614(G7614,G7511,G59112);
  nand GNAME7615(G7615,G7470,G20209);
  nand GNAME7616(G7616,G7469,G59118);
  nand GNAME7617(G7617,G3783,G59150);
  nand GNAME7618(G7618,G2791,G59309);
  nand GNAME7619(G7619,G2786,G7973,G7974);
  or GNAME7620(G7620,G3954,G2826);
  nand GNAME7621(G7621,G3886,G2794);
  nand GNAME7622(G7622,G3767,G3243,G7975,G7976);
  nand GNAME7623(G7623,G7622,G58979);
  nand GNAME7624(G7624,G2804,G3241);
  nand GNAME7625(G7625,G58979,G2899);
  nand GNAME7626(G7626,G3812,G7624,G7625,G3245);
  nand GNAME7627(G7627,G4224,G3956);
  nand GNAME7628(G7628,G7627,G59286);
  nand GNAME7629(G7629,G7626,G59127);
  nand GNAME7630(G7630,G59254,G3247);
  nand GNAME7631(G7631,G2836,G59159);
  nand GNAME7632(G7632,G2859,G21434);
  nand GNAME7633(G7633,G7627,G59285);
  nand GNAME7634(G7634,G7626,G59126);
  nand GNAME7635(G7635,G59253,G3247);
  nand GNAME7636(G7636,G2836,G59158);
  nand GNAME7637(G7637,G2859,G21435);
  nand GNAME7638(G7638,G7627,G59284);
  nand GNAME7639(G7639,G7626,G59125);
  nand GNAME7640(G7640,G59252,G3247);
  nand GNAME7641(G7641,G2836,G59157);
  nand GNAME7642(G7642,G2859,G21436);
  nand GNAME7643(G7643,G7627,G59283);
  nand GNAME7644(G7644,G7626,G59124);
  nand GNAME7645(G7645,G59251,G3247);
  nand GNAME7646(G7646,G2836,G59156);
  nand GNAME7647(G7647,G2859,G21437);
  nand GNAME7648(G7648,G7627,G59282);
  nand GNAME7649(G7649,G7626,G59123);
  nand GNAME7650(G7650,G59250,G3247);
  nand GNAME7651(G7651,G2836,G59155);
  nand GNAME7652(G7652,G2859,G21438);
  nand GNAME7653(G7653,G7627,G59281);
  nand GNAME7654(G7654,G7626,G59122);
  nand GNAME7655(G7655,G59249,G3247);
  nand GNAME7656(G7656,G2836,G59154);
  nand GNAME7657(G7657,G2859,G21439);
  nand GNAME7658(G7658,G7627,G59308);
  nand GNAME7659(G7659,G7626,G59149);
  nand GNAME7660(G7660,G59276,G3247);
  nand GNAME7661(G7661,G2836,G59181);
  nand GNAME7662(G7662,G7627,G59307);
  nand GNAME7663(G7663,G7626,G59148);
  nand GNAME7664(G7664,G59275,G3247);
  nand GNAME7665(G7665,G2836,G59180);
  nand GNAME7666(G7666,G2859,G21442);
  nand GNAME7667(G7667,G20108,G3241);
  nand GNAME7668(G7668,G3244,G3994,G7667);
  nand GNAME7669(G7669,G7668,G59109);
  nand GNAME7670(G7670,G7627,G59280);
  nand GNAME7671(G7671,G7626,G59121);
  nand GNAME7672(G7672,G59248,G3247);
  nand GNAME7673(G7673,G2836,G59153);
  nand GNAME7674(G7674,G2859,G21440);
  nand GNAME7675(G7675,G2816,G7882);
  nand GNAME7676(G7676,G2944,G2943);
  nand GNAME7677(G7677,G2805,G59114);
  nand GNAME7678(G7678,G7627,G59306);
  nand GNAME7679(G7679,G7626,G59147);
  nand GNAME7680(G7680,G59274,G3247);
  nand GNAME7681(G7681,G2836,G59179);
  nand GNAME7682(G7682,G2859,G21393);
  nand GNAME7683(G7683,G7627,G59305);
  nand GNAME7684(G7684,G7626,G59146);
  nand GNAME7685(G7685,G59273,G3247);
  nand GNAME7686(G7686,G2836,G59178);
  nand GNAME7687(G7687,G2859,G21392);
  nand GNAME7688(G7688,G7627,G59304);
  nand GNAME7689(G7689,G7626,G59145);
  nand GNAME7690(G7690,G59272,G3247);
  nand GNAME7691(G7691,G2836,G59177);
  nand GNAME7692(G7692,G2859,G21444);
  nand GNAME7693(G7693,G7627,G59303);
  nand GNAME7694(G7694,G7626,G59144);
  nand GNAME7695(G7695,G59271,G3247);
  nand GNAME7696(G7696,G2836,G59176);
  nand GNAME7697(G7697,G2859,G21391);
  nand GNAME7698(G7698,G7627,G59302);
  nand GNAME7699(G7699,G7626,G59143);
  nand GNAME7700(G7700,G59270,G3247);
  nand GNAME7701(G7701,G2836,G59175);
  nand GNAME7702(G7702,G2859,G21390);
  nand GNAME7703(G7703,G7627,G59301);
  nand GNAME7704(G7704,G7626,G59142);
  nand GNAME7705(G7705,G59269,G3247);
  nand GNAME7706(G7706,G2836,G59174);
  nand GNAME7707(G7707,G2859,G21468);
  nand GNAME7708(G7708,G7627,G59300);
  nand GNAME7709(G7709,G7626,G59141);
  nand GNAME7710(G7710,G59268,G3247);
  nand GNAME7711(G7711,G2836,G59173);
  nand GNAME7712(G7712,G2859,G21469);
  nand GNAME7713(G7713,G7627,G59299);
  nand GNAME7714(G7714,G7626,G59140);
  nand GNAME7715(G7715,G59267,G3247);
  nand GNAME7716(G7716,G2836,G59172);
  nand GNAME7717(G7717,G2859,G21470);
  nand GNAME7718(G7718,G7627,G59298);
  nand GNAME7719(G7719,G7626,G59139);
  nand GNAME7720(G7720,G59266,G3247);
  nand GNAME7721(G7721,G2836,G59171);
  nand GNAME7722(G7722,G2859,G21471);
  nand GNAME7723(G7723,G7627,G59297);
  nand GNAME7724(G7724,G7626,G59138);
  nand GNAME7725(G7725,G59265,G3247);
  nand GNAME7726(G7726,G2836,G59170);
  nand GNAME7727(G7727,G2859,G21472);
  nand GNAME7728(G7728,G7668,G59110);
  nand GNAME7729(G7729,G7627,G59279);
  nand GNAME7730(G7730,G7626,G59120);
  nand GNAME7731(G7731,G59247,G3247);
  nand GNAME7732(G7732,G2836,G59152);
  nand GNAME7733(G7733,G2859,G21443);
  nand GNAME7734(G7734,G7895,G2943);
  nand GNAME7735(G7735,G2816,G5069);
  nand GNAME7736(G7736,G2805,G59115);
  nand GNAME7737(G7737,G7627,G59296);
  nand GNAME7738(G7738,G7626,G59137);
  nand GNAME7739(G7739,G59264,G3247);
  nand GNAME7740(G7740,G2836,G59169);
  nand GNAME7741(G7741,G2859,G21474);
  nand GNAME7742(G7742,G7627,G59295);
  nand GNAME7743(G7743,G7626,G59136);
  nand GNAME7744(G7744,G59263,G3247);
  nand GNAME7745(G7745,G2836,G59168);
  nand GNAME7746(G7746,G2859,G21475);
  nand GNAME7747(G7747,G7627,G59294);
  nand GNAME7748(G7748,G7626,G59135);
  nand GNAME7749(G7749,G59262,G3247);
  nand GNAME7750(G7750,G2836,G59167);
  nand GNAME7751(G7751,G2859,G21476);
  nand GNAME7752(G7752,G7627,G59293);
  nand GNAME7753(G7753,G7626,G59134);
  nand GNAME7754(G7754,G59261,G3247);
  nand GNAME7755(G7755,G2836,G59166);
  nand GNAME7756(G7756,G2859,G21446);
  nand GNAME7757(G7757,G7627,G59292);
  nand GNAME7758(G7758,G7626,G59133);
  nand GNAME7759(G7759,G59260,G3247);
  nand GNAME7760(G7760,G2836,G59165);
  nand GNAME7761(G7761,G2859,G21447);
  nand GNAME7762(G7762,G7627,G59291);
  nand GNAME7763(G7763,G7626,G59132);
  nand GNAME7764(G7764,G59259,G3247);
  nand GNAME7765(G7765,G2836,G59164);
  nand GNAME7766(G7766,G2859,G21448);
  nand GNAME7767(G7767,G7627,G59290);
  nand GNAME7768(G7768,G7626,G59131);
  nand GNAME7769(G7769,G59258,G3247);
  nand GNAME7770(G7770,G2836,G59163);
  nand GNAME7771(G7771,G2859,G21449);
  nand GNAME7772(G7772,G7627,G59289);
  nand GNAME7773(G7773,G7626,G59130);
  nand GNAME7774(G7774,G59257,G3247);
  nand GNAME7775(G7775,G2836,G59162);
  nand GNAME7776(G7776,G2859,G21450);
  nand GNAME7777(G7777,G7627,G59288);
  nand GNAME7778(G7778,G7626,G59129);
  nand GNAME7779(G7779,G59256,G3247);
  nand GNAME7780(G7780,G2836,G59161);
  nand GNAME7781(G7781,G2859,G21451);
  nand GNAME7782(G7782,G7627,G59287);
  nand GNAME7783(G7783,G7626,G59128);
  nand GNAME7784(G7784,G59255,G3247);
  nand GNAME7785(G7785,G2836,G59160);
  nand GNAME7786(G7786,G2859,G21452);
  nand GNAME7787(G7787,G7668,G59111);
  nand GNAME7788(G7788,G7627,G59278);
  nand GNAME7789(G7789,G7626,G59119);
  nand GNAME7790(G7790,G59246,G3247);
  nand GNAME7791(G7791,G2836,G59151);
  nand GNAME7792(G7792,G2859,G21445);
  nand GNAME7793(G7793,G3253,G2816);
  nand GNAME7794(G7794,G7889,G2943);
  nand GNAME7795(G7795,G2805,G59116);
  nand GNAME7796(G7796,G7668,G59112);
  nand GNAME7797(G7797,G7627,G59277);
  nand GNAME7798(G7798,G7626,G59118);
  nand GNAME7799(G7799,G59245,G3247);
  nand GNAME7800(G7800,G2836,G59150);
  nand GNAME7801(G7801,G2859,G21453);
  nand GNAME7802(G7802,G5099,G2943);
  nand GNAME7803(G7803,G2816,G5047);
  nand GNAME7804(G7804,G2805,G59117);
  not GNAME7805(G7805,G3248);
  or GNAME7806(G7806,G2837,G7985);
  nand GNAME7807(G7807,G7214,G7805);
  nand GNAME7808(G7808,G7270,G7805);
  nand GNAME7809(G7809,G59109,G58976);
  nand GNAME7810(G7810,G2783,G3920);
  nand GNAME7811(G7811,G7810,G3793);
  nand GNAME7812(G7812,G7811,G3111);
  nand GNAME7813(G7813,G7326,G7805);
  nand GNAME7814(G7814,G59110,G58976);
  nand GNAME7815(G7815,G2783,G7977,G7978);
  nand GNAME7816(G7816,G7382,G7805);
  nand GNAME7817(G7817,G7438,G7805);
  nand GNAME7818(G7818,G3793,G3249);
  nand GNAME7819(G7819,G20804,G3250);
  nand GNAME7820(G7820,G58978,G2118);
  nand GNAME7821(G7821,G3250,G20818);
  nand GNAME7822(G7822,G58978,G21388);
  nand GNAME7823(G7823,G3250,G20819);
  nand GNAME7824(G7824,G58978,G21389);
  nand GNAME7825(G7825,G3250,G20820);
  nand GNAME7826(G7826,G58978,G21386);
  nand GNAME7827(G7827,G3250,G20817);
  nand GNAME7828(G7828,G58978,G21387);
  nand GNAME7829(G7829,G3250,G20805);
  nand GNAME7830(G7830,G2785,G3249);
  nand GNAME7831(G7831,G2837,G7830);
  nand GNAME7832(G7832,G58942,G6212,G6213);
  nand GNAME7833(G7833,G59349,G3113,G58943);
  nand GNAME7834(G7834,G58942,G1590,G6217);
  nand GNAME7835(G7835,G2785,G3186);
  nand GNAME7836(G7836,G7984,G59355);
  nand GNAME7837(G7837,G3772,G3961);
  nand GNAME7838(G7838,G59354,G7984);
  nand GNAME7839(G7839,G3772,G3962);
  nand GNAME7840(G7840,G3787,G59351);
  nand GNAME7841(G7841,G2814,G59355);
  or GNAME7842(G7842,G59352,G3787);
  nand GNAME7843(G7843,G3787,G59350);
  nand GNAME7844(G7844,G59349,G3773);
  or GNAME7845(G7845,G3773,G3990);
  nand GNAME7846(G7846,G2810,G35);
  nand GNAME7847(G7847,G3964,G59348);
  nand GNAME7848(G7848,G2784,G3852);
  nand GNAME7849(G7849,G2799,G3886);
  not GNAME7850(G7850,G3252);
  nand GNAME7851(G7851,G3787,G59345);
  or GNAME7852(G7852,G59354,G3787);
  nand GNAME7853(G7853,G7988,G59344);
  nand GNAME7854(G7854,G2832,G59309);
  nand GNAME7855(G7855,G2783,G2786,G2785);
  nand GNAME7856(G7856,G3835,G2786,G2749);
  nand GNAME7857(G7857,G2786,G2897);
  nand GNAME7858(G7858,G4844,G3903);
  nand GNAME7859(G7859,G2795,G4836,G3954);
  nand GNAME7860(G7860,G2748,G3869);
  nand GNAME7861(G7861,G2817,G2816);
  nand GNAME7862(G7862,G58978,G2754,G2790);
  nand GNAME7863(G7863,G2920,G58979,G20108);
  nand GNAME7864(G7864,G59117,G5043);
  nand GNAME7865(G7865,G2841,G59118);
  nand GNAME7866(G7866,G3285,G59118);
  nand GNAME7867(G7867,G7865,G7866);
  or GNAME7868(G7868,G59117,G58977);
  nand GNAME7869(G7869,G2816,G59117);
  or GNAME7870(G7870,G3285,G59119);
  or GNAME7871(G7871,G2841,G21592);
  nand GNAME7872(G7872,G2923,G3804);
  nand GNAME7873(G7873,G2922,G5054);
  nand GNAME7874(G7874,G5058,G3402);
  or GNAME7875(G7875,G5058,G3402);
  not GNAME7876(G7876,G3253);
  or GNAME7877(G7877,G2926,G2925);
  nand GNAME7878(G7878,G2925,G2926);
  not GNAME7879(G7879,G3254);
  or GNAME7880(G7880,G3776,G3775);
  nand GNAME7881(G7881,G3775,G3776);
  not GNAME7882(G7882,G3255);
  or GNAME7883(G7883,G2755,G3777);
  nand GNAME7884(G7884,G3777,G5119);
  or GNAME7885(G7885,G5097,G3778);
  nand GNAME7886(G7886,G3778,G5097);
  nand GNAME7887(G7887,G5122,G3403);
  or GNAME7888(G7888,G5122,G3403);
  not GNAME7889(G7889,G3256);
  or GNAME7890(G7890,G2759,G3777);
  nand GNAME7891(G7891,G3777,G5137);
  nand GNAME7892(G7892,G5163,G5166);
  nand GNAME7893(G7893,G2939,G7892);
  nand GNAME7894(G7894,G5141,G5163,G5166);
  not GNAME7895(G7895,G3267);
  nand GNAME7896(G7896,G2795,G59110);
  nand GNAME7897(G7897,G2764,G3869);
  not GNAME7898(G7898,G3258);
  nand GNAME7899(G7899,G5147,G59110);
  nand GNAME7900(G7900,G2764,G3779);
  not GNAME7901(G7901,G3257);
  or GNAME7902(G7902,G2764,G3777);
  nand GNAME7903(G7903,G3777,G5158);
  or GNAME7904(G7904,G2771,G3780);
  nand GNAME7905(G7905,G3780,G5173);
  or GNAME7906(G7906,G2771,G3777);
  nand GNAME7907(G7907,G3777,G5185);
  nand GNAME7908(G7908,G3777,G2865,G2793,G20523);
  or GNAME7909(G7909,G7985,G3777);
  nand GNAME7910(G7910,G6190,G58979);
  nand GNAME7911(G7911,G2790,G6191);
  or GNAME7912(G7912,G2790,G3110);
  nand GNAME7913(G7913,G3110,G6197);
  nand GNAME7914(G7914,G3964,G58945);
  nand GNAME7915(G7915,G2810,G6207);
  nand GNAME7916(G7916,G2810,G3774,G6206);
  nand GNAME7917(G7917,G3964,G58944);
  nand GNAME7918(G7918,G2807,G6210);
  nand GNAME7919(G7919,G58942,G6208,G58943);
  or GNAME7920(G7920,G2809,G2751,G58942,G59349);
  nand GNAME7921(G7921,G2809,G3112,G58941);
  nand GNAME7922(G7922,G3787,G58910);
  nand GNAME7923(G7923,G2814,G59344);
  nand GNAME7924(G7924,G3787,G58909);
  nand GNAME7925(G7925,G2814,G59343);
  nand GNAME7926(G7926,G3787,G58908);
  nand GNAME7927(G7927,G2814,G59342);
  nand GNAME7928(G7928,G3787,G58907);
  nand GNAME7929(G7929,G2814,G59341);
  nand GNAME7930(G7930,G2764,G59111);
  nand GNAME7931(G7931,G2759,G59110);
  not GNAME7932(G7932,G3259);
  nand GNAME7933(G7933,G2759,G59109);
  nand GNAME7934(G7934,G59111,G2765);
  or GNAME7935(G7935,G59346,G2764);
  nand GNAME7936(G7936,G59346,G7867,G5069);
  or GNAME7937(G7937,G59346,G2759);
  nand GNAME7938(G7938,G59346,G7867,G3253);
  or GNAME7939(G7939,G59346,G2755);
  nand GNAME7940(G7940,G5115,G59346);
  nand GNAME7941(G7941,G3781,G20523,G2865);
  or GNAME7942(G7942,G7985,G3781);
  or GNAME7943(G7943,G2771,G3781);
  nand GNAME7944(G7944,G3781,G5182);
  or GNAME7945(G7945,G2764,G3781);
  nand GNAME7946(G7946,G3781,G5154);
  or GNAME7947(G7947,G2759,G3781);
  nand GNAME7948(G7948,G3781,G5133);
  or GNAME7949(G7949,G2755,G3781);
  nand GNAME7950(G7950,G3781,G5114);
  nand GNAME7951(G7951,G2817,G59308);
  nand GNAME7952(G7952,G58978,G59149);
  nand GNAME7953(G7953,G3869,G59148);
  nand GNAME7954(G7954,G2795,G6718);
  nand GNAME7955(G7955,G3869,G59147);
  nand GNAME7956(G7956,G2795,G6735);
  nand GNAME7957(G7957,G3869,G59146);
  nand GNAME7958(G7958,G2795,G6752);
  nand GNAME7959(G7959,G3869,G59145);
  nand GNAME7960(G7960,G2795,G6769);
  nand GNAME7961(G7961,G3869,G59144);
  nand GNAME7962(G7962,G2795,G6786);
  nand GNAME7963(G7963,G3869,G59143);
  nand GNAME7964(G7964,G2795,G6803);
  nand GNAME7965(G7965,G3869,G59142);
  nand GNAME7966(G7966,G2795,G6820);
  nand GNAME7967(G7967,G3869,G59141);
  nand GNAME7968(G7968,G2795,G6837);
  nand GNAME7969(G7969,G3954,G3920);
  nand GNAME7970(G7970,G2749,G2863);
  nand GNAME7971(G7971,G2795,G3954);
  nand GNAME7972(G7972,G2787,G3869);
  nand GNAME7973(G7973,G2785,G3835);
  nand GNAME7974(G7974,G2783,G2749);
  nand GNAME7975(G7975,G2799,G2890);
  nand GNAME7976(G7976,G3852,G3937);
  nand GNAME7977(G7977,G2785,G3852);
  nand GNAME7978(G7978,G2799,G3954);
  nand GNAME7979(G7979,G59111,G58976);
  nand GNAME7980(G7980,G2837,G7815);
  nand GNAME7981(G7981,G59112,G58976);
  nand GNAME7982(G7982,G2837,G7811);
  not GNAME7983(G7983,G2806);
  not GNAME7984(G7984,G3772);
  not GNAME7985(G7985,G59108);
  not GNAME7986(G7986,G2947);
  not GNAME7987(G7987,G2911);
  not GNAME7988(G7988,G2832);
  not GNAME7989(G7989,G2797);
  not GNAME7990(G7990,G3188);
  or GNAME7991(G7991,G8076,G14027);
  or GNAME7992(G7992,G14000,G8092);
  nand GNAME7993(G7993,G14000,G8092);
  or GNAME7994(G7994,G14279,G13999);
  nand GNAME7995(G7995,G13999,G14279);
  or GNAME7996(G7996,G13998,G8093);
  nand GNAME7997(G7997,G13998,G8093);
  or GNAME7998(G7998,G14278,G13997);
  nand GNAME7999(G7999,G13997,G14278);
  or GNAME8000(G8000,G13996,G8094);
  nand GNAME8001(G8001,G13996,G8094);
  or GNAME8002(G8002,G14277,G13995);
  nand GNAME8003(G8003,G13995,G14277);
  or GNAME8004(G8004,G13994,G8095);
  nand GNAME8005(G8005,G13994,G8095);
  or GNAME8006(G8006,G15287,G13993);
  nand GNAME8007(G8007,G13993,G15287);
  or GNAME8008(G8008,G15286,G8082);
  nand GNAME8009(G8009,G8082,G15286);
  nand GNAME8010(G8010,G8066,G15283);
  or GNAME8011(G8011,G15283,G8066);
  nand GNAME8012(G8012,G8084,G8032);
  nand GNAME8013(G8013,G8083,G14297);
  or GNAME8014(G8014,G15280,G2085);
  nand GNAME8015(G8015,G2085,G15280);
  or GNAME8016(G8016,G14276,G8085);
  nand GNAME8017(G8017,G8085,G14276);
  nand GNAME8018(G8018,G14025,G8064);
  nand GNAME8019(G8019,G14028,G14296);
  nand GNAME8020(G8020,G14023,G14024);
  or GNAME8021(G8021,G14024,G14023);
  nand GNAME8022(G8022,G14022,G8086);
  or GNAME8023(G8023,G8086,G14022);
  nand GNAME8024(G8024,G2086,G14293);
  or GNAME8025(G8025,G14293,G2086);
  nand GNAME8026(G8026,G14018,G14020);
  or GNAME8027(G8027,G14020,G14018);
  nand GNAME8028(G8028,G14019,G8087);
  or GNAME8029(G8029,G8087,G14019);
  or GNAME8030(G8030,G14017,G14016);
  nand GNAME8031(G8031,G14016,G14017);
  not GNAME8032(G8032,G8083);
  nor GNAME8033(G8033,G8034,G15285);
  and GNAME8034(G8034,G8082,G15286);
  or GNAME8035(G8035,G15284,G13992);
  nor GNAME8036(G8036,G8037,G15282);
  and GNAME8037(G8037,G15283,G13991);
  or GNAME8038(G8038,G15281,G13990);
  or GNAME8039(G8039,G13994,G13993);
  nand GNAME8040(G8040,G8041,G15287);
  nand GNAME8041(G8041,G13993,G13994);
  or GNAME8042(G8042,G13996,G13995);
  nand GNAME8043(G8043,G8044,G14277);
  nand GNAME8044(G8044,G13995,G13996);
  or GNAME8045(G8045,G13998,G13997);
  nand GNAME8046(G8046,G8047,G14278);
  nand GNAME8047(G8047,G13997,G13998);
  or GNAME8048(G8048,G14000,G13999);
  nand GNAME8049(G8049,G8050,G14279);
  nand GNAME8050(G8050,G13999,G14000);
  or GNAME8051(G8051,G14002,G14001);
  nand GNAME8052(G8052,G8053,G14280);
  nand GNAME8053(G8053,G14001,G14002);
  or GNAME8054(G8054,G14004,G14003);
  nand GNAME8055(G8055,G8056,G14281);
  nand GNAME8056(G8056,G14003,G14004);
  or GNAME8057(G8057,G14006,G14005);
  nand GNAME8058(G8058,G8059,G14282);
  nand GNAME8059(G8059,G14005,G14006);
  nand GNAME8060(G8060,G14307,G14283);
  nand GNAME8061(G8061,G8062,G14008);
  or GNAME8062(G8062,G14283,G14307);
  not GNAME8063(G8063,G14015);
  not GNAME8064(G8064,G14028);
  nand GNAME8065(G8065,G8084,G8069);
  not GNAME8066(G8066,G13991);
  not GNAME8067(G8067,G14010);
  not GNAME8068(G8068,G14012);
  nand GNAME8069(G8069,G14298,G14299);
  and GNAME8070(G8070,G8063,G14289);
  and GNAME8071(G8071,G14287,G14012);
  and GNAME8072(G8072,G14285,G14010);
  and GNAME8073(G8073,G2106,G2105);
  and GNAME8074(G8074,G2110,G2109);
  and GNAME8075(G8075,G2114,G2113);
  and GNAME8076(G8076,G14299,G15863);
  and GNAME8077(G8077,G7993,G7992);
  and GNAME8078(G8078,G7997,G7996);
  and GNAME8079(G8079,G8001,G8000);
  and GNAME8080(G8080,G8005,G8004);
  and GNAME8081(G8081,G8009,G8008);
  nand GNAME8082(G8082,G8040,G8039);
  nand GNAME8083(G8083,G8069,G15863);
  not GNAME8084(G8084,G14297);
  nand GNAME8085(G8085,G13989,G15280);
  and GNAME8086(G8086,G14024,G14295);
  and GNAME8087(G8087,G14020,G14292);
  and GNAME8088(G8088,G2104,G2103);
  and GNAME8089(G8089,G2108,G2107);
  and GNAME8090(G8090,G2112,G2111);
  and GNAME8091(G8091,G2116,G2115);
  and GNAME8092(G8092,G7995,G7994);
  and GNAME8093(G8093,G7999,G7998);
  and GNAME8094(G8094,G8003,G8002);
  and GNAME8095(G8095,G8007,G8006);
  nand GNAME8096(G8096,G2088,G2087);
  nand GNAME8097(G8097,G2090,G2089);
  nand GNAME8098(G8098,G2092,G2091);
  nand GNAME8099(G8099,G2094,G2093);
  nand GNAME8100(G8100,G2096,G2095);
  nand GNAME8101(G8101,G2098,G2097);
  nand GNAME8102(G8102,G2100,G2099);
  nand GNAME8103(G8103,G2102,G2101);
  nand GNAME8104(G8104,G7991,G2117);
  nand GNAME8105(G8105,G8011,G8010);
  nand GNAME8106(G8106,G8013,G8012);
  nand GNAME8107(G8107,G8015,G8014);
  nand GNAME8108(G8108,G8017,G8016);
  nand GNAME8109(G8109,G8019,G8018);
  nand GNAME8110(G8110,G8021,G8020);
  nand GNAME8111(G8111,G8023,G8022);
  nand GNAME8112(G8112,G8025,G8024);
  nand GNAME8113(G8113,G8027,G8026);
  nand GNAME8114(G8114,G8029,G8028);
  nor GNAME8115(G8115,G59795,G13982);
  nor GNAME8116(G8116,G59795,G8768);
  nand GNAME8117(G8117,G9533,G9534,G9535,G9536);
  nand GNAME8118(G8118,G9537,G9538,G9539,G9540);
  nand GNAME8119(G8119,G9541,G9542,G9543,G9544);
  nand GNAME8120(G8120,G9545,G9546,G9547,G9548);
  nand GNAME8121(G8121,G9549,G9550,G9551,G9552);
  nand GNAME8122(G8122,G9553,G9554,G9555,G9556);
  nand GNAME8123(G8123,G9557,G9558,G9559,G9560);
  nand GNAME8124(G8124,G9561,G9562,G9563,G9564);
  nand GNAME8125(G8125,G9565,G9566,G9567,G9568);
  nand GNAME8126(G8126,G9569,G9570,G9571,G9572);
  nand GNAME8127(G8127,G9573,G9574,G9575,G9576);
  nand GNAME8128(G8128,G9577,G9578,G9579,G9580);
  nand GNAME8129(G8129,G9581,G9582,G9583,G9584);
  nand GNAME8130(G8130,G9585,G9586,G9587,G9588);
  nand GNAME8131(G8131,G9589,G9590,G9591,G9592);
  nand GNAME8132(G8132,G9593,G9594,G9595,G9596);
  nand GNAME8133(G8133,G13828,G8814);
  nand GNAME8134(G8134,G13816,G13817);
  or GNAME8135(G8135,G8134,G13802);
  nand GNAME8136(G8136,G13818,G9245,G13817);
  nand GNAME8137(G8137,G9248,G13819,G13820);
  nand GNAME8138(G8138,G9248,G13821,G13822);
  nand GNAME8139(G8139,G9248,G13823,G13824);
  nand GNAME8140(G8140,G9248,G13825,G13826);
  and GNAME8141(G8141,G13012,G13802);
  and GNAME8142(G8142,G13067,G13802);
  and GNAME8143(G8143,G13122,G13802);
  nand GNAME8144(G8144,G13803,G13804);
  nand GNAME8145(G8145,G13805,G13806);
  nand GNAME8146(G8146,G13811,G13809,G13810);
  nand GNAME8147(G8147,G13976,G13977,G8814,G13813);
  nand GNAME8148(G8148,G13978,G13979,G8814,G13814);
  nand GNAME8149(G8149,G13655,G13656,G13657,G13658);
  nand GNAME8150(G8150,G13662,G13663,G13661,G13659,G13660);
  nand GNAME8151(G8151,G13678,G13679,G13677,G13675,G13676);
  nand GNAME8152(G8152,G13683,G13684,G13682,G13680,G13681);
  nand GNAME8153(G8153,G13688,G13689,G13687,G13685,G13686);
  nand GNAME8154(G8154,G13693,G13694,G13692,G13690,G13691);
  nand GNAME8155(G8155,G13698,G13699,G13697,G13695,G13696);
  nand GNAME8156(G8156,G13703,G13704,G13702,G13700,G13701);
  nand GNAME8157(G8157,G13708,G13709,G13707,G13705,G13706);
  nand GNAME8158(G8158,G13713,G13714,G13712,G13710,G13711);
  nand GNAME8159(G8159,G13718,G13719,G13717,G13715,G13716);
  nand GNAME8160(G8160,G13723,G13724,G13722,G13720,G13721);
  nand GNAME8161(G8161,G13737,G13738,G13736,G13734,G13735);
  nand GNAME8162(G8162,G13742,G13743,G13741,G13739,G13740);
  nand GNAME8163(G8163,G13747,G13748,G13746,G13744,G13745);
  nand GNAME8164(G8164,G13752,G13753,G13751,G13749,G13750);
  nand GNAME8165(G8165,G13757,G13758,G13756,G13754,G13755);
  nand GNAME8166(G8166,G13762,G13763,G13761,G13759,G13760);
  nand GNAME8167(G8167,G13767,G13768,G13766,G13764,G13765);
  nand GNAME8168(G8168,G13772,G13773,G13771,G13769,G13770);
  nand GNAME8169(G8169,G13777,G13778,G13776,G13774,G13775);
  nand GNAME8170(G8170,G13782,G13783,G13781,G13779,G13780);
  nand GNAME8171(G8171,G13628,G13629,G13627,G13625,G13626);
  nand GNAME8172(G8172,G13633,G13634,G13632,G13630,G13631);
  nand GNAME8173(G8173,G13638,G13639,G13637,G13635,G13636);
  nand GNAME8174(G8174,G13643,G13644,G13642,G13640,G13641);
  nand GNAME8175(G8175,G13648,G13649,G13647,G13645,G13646);
  nand GNAME8176(G8176,G13653,G13654,G13652,G13650,G13651);
  nand GNAME8177(G8177,G9765,G13666,G13672,G13673,G13668);
  nand GNAME8178(G8178,G9766,G13725,G13731,G13732,G13727);
  nand GNAME8179(G8179,G9767,G13784,G13790,G13791,G13786);
  nand GNAME8180(G8180,G9768,G13793,G13799,G13800,G13795);
  and GNAME8181(G8181,G8125,G8856);
  and GNAME8182(G8182,G8126,G8856);
  and GNAME8183(G8183,G8127,G8856);
  and GNAME8184(G8184,G8128,G8856);
  and GNAME8185(G8185,G8129,G8856);
  and GNAME8186(G8186,G8130,G8856);
  and GNAME8187(G8187,G8131,G8856);
  and GNAME8188(G8188,G8132,G8856);
  nand GNAME8189(G8189,G8872,G9239,G9991,G9796,G9809);
  nand GNAME8190(G8190,G9797,G9991,G13620,G9243);
  nand GNAME8191(G8191,G13495,G13496,G13497,G13498);
  nand GNAME8192(G8192,G13502,G13503,G13501,G13499,G13500);
  nand GNAME8193(G8193,G13517,G13518,G13516,G13514,G13515);
  nand GNAME8194(G8194,G13522,G13523,G13521,G13519,G13520);
  nand GNAME8195(G8195,G13527,G13528,G13526,G13524,G13525);
  nand GNAME8196(G8196,G13532,G13533,G13531,G13529,G13530);
  nand GNAME8197(G8197,G13537,G13538,G13536,G13534,G13535);
  nand GNAME8198(G8198,G13542,G13543,G13541,G13539,G13540);
  nand GNAME8199(G8199,G13547,G13548,G13546,G13544,G13545);
  nand GNAME8200(G8200,G13549,G13550,G13551,G13552);
  nand GNAME8201(G8201,G13553,G13554,G13555,G13556);
  nand GNAME8202(G8202,G13557,G13558,G13559,G13560);
  nand GNAME8203(G8203,G13566,G13567,G13568,G13569);
  nand GNAME8204(G8204,G13570,G13571,G13572,G13573);
  nand GNAME8205(G8205,G13574,G13575,G13576,G13577);
  nand GNAME8206(G8206,G13578,G13579,G13580,G13581);
  nand GNAME8207(G8207,G13582,G13583,G13584,G13585);
  nand GNAME8208(G8208,G13586,G13587,G13588,G13589);
  nand GNAME8209(G8209,G13590,G13591,G13592,G13593);
  nand GNAME8210(G8210,G13594,G13595,G13596,G13597);
  nand GNAME8211(G8211,G13598,G13599,G13600,G13601);
  nand GNAME8212(G8212,G13602,G13603,G13604,G13605);
  nand GNAME8213(G8213,G13468,G13469,G13470,G13471);
  nand GNAME8214(G8214,G13472,G13473,G13474,G13475);
  nand GNAME8215(G8215,G13476,G13477,G13478,G13479);
  nand GNAME8216(G8216,G13480,G13481,G13482,G13483);
  nand GNAME8217(G8217,G13484,G13485,G13486,G13487);
  nand GNAME8218(G8218,G13493,G13494,G13492,G13490,G13491);
  nand GNAME8219(G8219,G13512,G13513,G13511,G13509,G13510);
  nand GNAME8220(G8220,G13564,G13565,G13563,G13561,G13562);
  nand GNAME8221(G8221,G13609,G13610,G13608,G13606,G13607);
  nand GNAME8222(G8222,G13614,G13615,G13613,G13611,G13612);
  and GNAME8223(G8223,G13029,G8864);
  and GNAME8224(G8224,G13084,G8864);
  and GNAME8225(G8225,G13139,G8864);
  and GNAME8226(G8226,G13177,G8864);
  and GNAME8227(G8227,G13233,G8864);
  and GNAME8228(G8228,G13289,G8864);
  and GNAME8229(G8229,G13345,G8864);
  and GNAME8230(G8230,G13401,G8864);
  and GNAME8231(G8231,G59549,G8856);
  and GNAME8232(G8232,G59550,G8856);
  and GNAME8233(G8233,G59551,G8856);
  and GNAME8234(G8234,G59552,G8856);
  and GNAME8235(G8235,G59553,G8856);
  nand GNAME8236(G8236,G13442,G9795,G13441);
  nand GNAME8237(G8237,G9239,G9761,G9953,G9799,G9807);
  nand GNAME8238(G8238,G9797,G13441,G13449,G13450);
  nand GNAME8239(G8239,G13047,G13048,G13049,G13050);
  nand GNAME8240(G8240,G13102,G13103,G13104,G13105);
  nand GNAME8241(G8241,G13157,G13158,G13159,G13160);
  nand GNAME8242(G8242,G13215,G13216,G13214,G13212,G13213);
  nand GNAME8243(G8243,G13271,G13272,G13270,G13268,G13269);
  nand GNAME8244(G8244,G9734,G13325,G9791,G13324);
  nand GNAME8245(G8245,G9747,G9782,G9185,G13380,G13381);
  nand GNAME8246(G8246,G9760,G9791,G9805,G13436,G13437);
  nand GNAME8247(G8247,G12867,G12868,G12869,G12870);
  nand GNAME8248(G8248,G12874,G12875,G12873,G12871,G12872);
  nand GNAME8249(G8249,G12884,G12885,G12883,G12881,G12882);
  nand GNAME8250(G8250,G12889,G12890,G12888,G12886,G12887);
  nand GNAME8251(G8251,G12894,G12895,G12893,G12891,G12892);
  nand GNAME8252(G8252,G12899,G12900,G12898,G12896,G12897);
  nand GNAME8253(G8253,G12904,G12905,G12903,G12901,G12902);
  nand GNAME8254(G8254,G12909,G12910,G12908,G12906,G12907);
  nand GNAME8255(G8255,G12914,G12915,G12913,G12911,G12912);
  nand GNAME8256(G8256,G12919,G12920,G12918,G12916,G12917);
  nand GNAME8257(G8257,G12924,G12925,G12923,G12921,G12922);
  nand GNAME8258(G8258,G12929,G12930,G12928,G12926,G12927);
  nand GNAME8259(G8259,G12939,G12940,G12938,G12936,G12937);
  nand GNAME8260(G8260,G12944,G12945,G12943,G12941,G12942);
  nand GNAME8261(G8261,G12949,G12950,G12948,G12946,G12947);
  nand GNAME8262(G8262,G12954,G12955,G12953,G12951,G12952);
  nand GNAME8263(G8263,G12959,G12960,G12958,G12956,G12957);
  nand GNAME8264(G8264,G12964,G12965,G12963,G12961,G12962);
  nand GNAME8265(G8265,G12969,G12970,G12968,G12966,G12967);
  nand GNAME8266(G8266,G12974,G12975,G12973,G12971,G12972);
  nand GNAME8267(G8267,G12979,G12980,G12978,G12976,G12977);
  nand GNAME8268(G8268,G12984,G12985,G12983,G12981,G12982);
  nand GNAME8269(G8269,G12840,G12841,G12839,G12837,G12838);
  nand GNAME8270(G8270,G12845,G12846,G12844,G12842,G12843);
  nand GNAME8271(G8271,G12850,G12851,G12849,G12847,G12848);
  nand GNAME8272(G8272,G12855,G12856,G12854,G12852,G12853);
  nand GNAME8273(G8273,G12860,G12861,G12859,G12857,G12858);
  nand GNAME8274(G8274,G12865,G12866,G12864,G12862,G12863);
  nand GNAME8275(G8275,G12879,G12880,G12878,G12876,G12877);
  nand GNAME8276(G8276,G12934,G12935,G12933,G12931,G12932);
  nand GNAME8277(G8277,G12989,G12990,G12988,G12986,G12987);
  nand GNAME8278(G8278,G9661,G12993,G12991,G12992);
  and GNAME8279(G8279,G9866,G59598);
  and GNAME8280(G8280,G9866,G59589);
  and GNAME8281(G8281,G9866,G59588);
  and GNAME8282(G8282,G9866,G59587);
  and GNAME8283(G8283,G9866,G59586);
  and GNAME8284(G8284,G9866,G59585);
  and GNAME8285(G8285,G9866,G59584);
  and GNAME8286(G8286,G9866,G59583);
  and GNAME8287(G8287,G9866,G59582);
  and GNAME8288(G8288,G9866,G59581);
  and GNAME8289(G8289,G9866,G59580);
  and GNAME8290(G8290,G9866,G59579);
  and GNAME8291(G8291,G9866,G59578);
  and GNAME8292(G8292,G9866,G59577);
  and GNAME8293(G8293,G9866,G59576);
  and GNAME8294(G8294,G9866,G59575);
  and GNAME8295(G8295,G9866,G59574);
  and GNAME8296(G8296,G9866,G59573);
  and GNAME8297(G8297,G9866,G59572);
  and GNAME8298(G8298,G9866,G59571);
  and GNAME8299(G8299,G9866,G59570);
  and GNAME8300(G8300,G9866,G59569);
  and GNAME8301(G8301,G9866,G59568);
  and GNAME8302(G8302,G9866,G59567);
  and GNAME8303(G8303,G8792,G12579);
  and GNAME8304(G8304,G8792,G12596);
  and GNAME8305(G8305,G8792,G12613);
  and GNAME8306(G8306,G8792,G12630);
  and GNAME8307(G8307,G8792,G12647);
  and GNAME8308(G8308,G8792,G12664);
  and GNAME8309(G8309,G8792,G12681);
  and GNAME8310(G8310,G8792,G12698);
  nand GNAME8311(G8311,G12305,G12303,G12304);
  nand GNAME8312(G8312,G12302,G12300,G12301);
  nand GNAME8313(G8313,G12299,G12297,G12298);
  nand GNAME8314(G8314,G12296,G12294,G12295);
  nand GNAME8315(G8315,G12293,G12291,G12292);
  nand GNAME8316(G8316,G12290,G12288,G12289);
  nand GNAME8317(G8317,G12287,G12285,G12286);
  nand GNAME8318(G8318,G12284,G12282,G12283);
  nand GNAME8319(G8319,G12281,G12279,G12280);
  nand GNAME8320(G8320,G12278,G12276,G12277);
  nand GNAME8321(G8321,G12275,G12273,G12274);
  nand GNAME8322(G8322,G12272,G12270,G12271);
  nand GNAME8323(G8323,G12269,G12267,G12268);
  nand GNAME8324(G8324,G12266,G12264,G12265);
  nand GNAME8325(G8325,G12263,G12261,G12262);
  nand GNAME8326(G8326,G12260,G12258,G12259);
  nand GNAME8327(G8327,G12257,G12255,G12256);
  nand GNAME8328(G8328,G12254,G12252,G12253);
  nand GNAME8329(G8329,G12251,G12249,G12250);
  nand GNAME8330(G8330,G12248,G12246,G12247);
  nand GNAME8331(G8331,G12245,G12243,G12244);
  nand GNAME8332(G8332,G12242,G12240,G12241);
  nand GNAME8333(G8333,G12239,G12237,G12238);
  nand GNAME8334(G8334,G12236,G12234,G12235);
  nand GNAME8335(G8335,G12233,G12231,G12232);
  nand GNAME8336(G8336,G12230,G12228,G12229);
  nand GNAME8337(G8337,G12227,G12225,G12226);
  nand GNAME8338(G8338,G12224,G12222,G12223);
  nand GNAME8339(G8339,G12221,G12219,G12220);
  nand GNAME8340(G8340,G12218,G12216,G12217);
  nand GNAME8341(G8341,G9786,G12215,G13831,G13917,G13918);
  nand GNAME8342(G8342,G9785,G12211,G13829,G13830);
  nand GNAME8343(G8343,G13915,G13916,G12203,G12208);
  and GNAME8344(G8344,G9961,G59395);
  and GNAME8345(G8345,G9961,G59396);
  and GNAME8346(G8346,G9961,G59397);
  and GNAME8347(G8347,G9961,G59398);
  and GNAME8348(G8348,G9961,G59399);
  and GNAME8349(G8349,G9961,G59400);
  and GNAME8350(G8350,G9961,G59401);
  and GNAME8351(G8351,G9961,G59402);
  and GNAME8352(G8352,G9961,G59403);
  and GNAME8353(G8353,G9961,G59404);
  and GNAME8354(G8354,G9961,G59405);
  and GNAME8355(G8355,G9961,G59406);
  and GNAME8356(G8356,G9961,G59407);
  and GNAME8357(G8357,G9961,G59408);
  and GNAME8358(G8358,G9961,G59409);
  and GNAME8359(G8359,G9961,G59410);
  and GNAME8360(G8360,G9961,G59411);
  and GNAME8361(G8361,G9961,G59412);
  and GNAME8362(G8362,G9961,G59413);
  and GNAME8363(G8363,G9961,G59414);
  and GNAME8364(G8364,G9961,G59415);
  and GNAME8365(G8365,G9961,G59416);
  and GNAME8366(G8366,G9961,G59417);
  and GNAME8367(G8367,G9961,G59418);
  and GNAME8368(G8368,G9961,G59419);
  and GNAME8369(G8369,G9961,G59420);
  and GNAME8370(G8370,G9961,G59421);
  and GNAME8371(G8371,G9961,G59422);
  and GNAME8372(G8372,G9961,G59423);
  and GNAME8373(G8373,G9961,G59424);
  nand GNAME8374(G8374,G12202,G8909,G13984);
  nand GNAME8375(G8375,G9798,G9799,G12200,G12201);
  nand GNAME8376(G8376,G12199,G9811,G12198);
  nand GNAME8377(G8377,G13909,G13910,G9810,G9812);
  nand GNAME8378(G8378,G9531,G12179,G12177,G12178);
  nand GNAME8379(G8379,G9530,G12173,G12171,G12172);
  nand GNAME8380(G8380,G9529,G12167,G12165,G12166);
  nand GNAME8381(G8381,G9528,G12161,G12159,G12160);
  nand GNAME8382(G8382,G9527,G12155,G12153,G12154);
  nand GNAME8383(G8383,G9526,G12149,G12147,G12148);
  nand GNAME8384(G8384,G9525,G12143,G12141,G12142);
  nand GNAME8385(G8385,G9524,G12137,G12135,G12136);
  nand GNAME8386(G8386,G9523,G12118,G12116,G12117);
  nand GNAME8387(G8387,G9522,G12112,G12110,G12111);
  nand GNAME8388(G8388,G9521,G12106,G12104,G12105);
  nand GNAME8389(G8389,G9520,G12100,G12098,G12099);
  nand GNAME8390(G8390,G9519,G12094,G12092,G12093);
  nand GNAME8391(G8391,G9518,G12088,G12086,G12087);
  nand GNAME8392(G8392,G9517,G12082,G12080,G12081);
  nand GNAME8393(G8393,G9516,G12076,G12074,G12075);
  nand GNAME8394(G8394,G9515,G12057,G12055,G12056);
  nand GNAME8395(G8395,G9514,G12051,G12049,G12050);
  nand GNAME8396(G8396,G9513,G12045,G12043,G12044);
  nand GNAME8397(G8397,G9512,G12039,G12037,G12038);
  nand GNAME8398(G8398,G9511,G12033,G12031,G12032);
  nand GNAME8399(G8399,G9510,G12027,G12025,G12026);
  nand GNAME8400(G8400,G9509,G12021,G12019,G12020);
  nand GNAME8401(G8401,G9508,G12015,G12013,G12014);
  nand GNAME8402(G8402,G9507,G11996,G11994,G11995);
  nand GNAME8403(G8403,G9506,G11990,G11988,G11989);
  nand GNAME8404(G8404,G9505,G11984,G11982,G11983);
  nand GNAME8405(G8405,G9504,G11978,G11976,G11977);
  nand GNAME8406(G8406,G9503,G11972,G11970,G11971);
  nand GNAME8407(G8407,G9502,G11966,G11964,G11965);
  nand GNAME8408(G8408,G9501,G11960,G11958,G11959);
  nand GNAME8409(G8409,G9500,G11954,G11952,G11953);
  nand GNAME8410(G8410,G9499,G11935,G11933,G11934);
  nand GNAME8411(G8411,G9498,G11929,G11927,G11928);
  nand GNAME8412(G8412,G9497,G11923,G11921,G11922);
  nand GNAME8413(G8413,G9496,G11917,G11915,G11916);
  nand GNAME8414(G8414,G9495,G11911,G11909,G11910);
  nand GNAME8415(G8415,G9494,G11905,G11903,G11904);
  nand GNAME8416(G8416,G9493,G11899,G11897,G11898);
  nand GNAME8417(G8417,G9492,G11893,G11891,G11892);
  nand GNAME8418(G8418,G9491,G11874,G11872,G11873);
  nand GNAME8419(G8419,G9490,G11868,G11866,G11867);
  nand GNAME8420(G8420,G9489,G11862,G11860,G11861);
  nand GNAME8421(G8421,G9488,G11856,G11854,G11855);
  nand GNAME8422(G8422,G9487,G11850,G11848,G11849);
  nand GNAME8423(G8423,G9486,G11844,G11842,G11843);
  nand GNAME8424(G8424,G9485,G11838,G11836,G11837);
  nand GNAME8425(G8425,G9484,G11832,G11830,G11831);
  nand GNAME8426(G8426,G9483,G11813,G11811,G11812);
  nand GNAME8427(G8427,G9482,G11807,G11805,G11806);
  nand GNAME8428(G8428,G9481,G11801,G11799,G11800);
  nand GNAME8429(G8429,G9480,G11795,G11793,G11794);
  nand GNAME8430(G8430,G9479,G11789,G11787,G11788);
  nand GNAME8431(G8431,G9478,G11783,G11781,G11782);
  nand GNAME8432(G8432,G9477,G11777,G11775,G11776);
  nand GNAME8433(G8433,G9476,G11771,G11769,G11770);
  nand GNAME8434(G8434,G9475,G11752,G11750,G11751);
  nand GNAME8435(G8435,G9474,G11746,G11744,G11745);
  nand GNAME8436(G8436,G9473,G11740,G11738,G11739);
  nand GNAME8437(G8437,G9472,G11734,G11732,G11733);
  nand GNAME8438(G8438,G9471,G11728,G11726,G11727);
  nand GNAME8439(G8439,G9470,G11722,G11720,G11721);
  nand GNAME8440(G8440,G9469,G11716,G11714,G11715);
  nand GNAME8441(G8441,G9468,G11710,G11708,G11709);
  nand GNAME8442(G8442,G9467,G11691,G11689,G11690);
  nand GNAME8443(G8443,G9466,G11685,G11683,G11684);
  nand GNAME8444(G8444,G9465,G11679,G11677,G11678);
  nand GNAME8445(G8445,G9464,G11673,G11671,G11672);
  nand GNAME8446(G8446,G9463,G11667,G11665,G11666);
  nand GNAME8447(G8447,G9462,G11661,G11659,G11660);
  nand GNAME8448(G8448,G9461,G11655,G11653,G11654);
  nand GNAME8449(G8449,G9460,G11649,G11647,G11648);
  nand GNAME8450(G8450,G9459,G11630,G11628,G11629);
  nand GNAME8451(G8451,G9458,G11624,G11622,G11623);
  nand GNAME8452(G8452,G9457,G11618,G11616,G11617);
  nand GNAME8453(G8453,G9456,G11612,G11610,G11611);
  nand GNAME8454(G8454,G9455,G11606,G11604,G11605);
  nand GNAME8455(G8455,G9454,G11600,G11598,G11599);
  nand GNAME8456(G8456,G9453,G11594,G11592,G11593);
  nand GNAME8457(G8457,G9452,G11588,G11586,G11587);
  nand GNAME8458(G8458,G9451,G11569,G11567,G11568);
  nand GNAME8459(G8459,G9450,G11563,G11561,G11562);
  nand GNAME8460(G8460,G9449,G11557,G11555,G11556);
  nand GNAME8461(G8461,G9448,G11551,G11549,G11550);
  nand GNAME8462(G8462,G9447,G11545,G11543,G11544);
  nand GNAME8463(G8463,G9446,G11539,G11537,G11538);
  nand GNAME8464(G8464,G9445,G11533,G11531,G11532);
  nand GNAME8465(G8465,G9444,G11527,G11525,G11526);
  nand GNAME8466(G8466,G9443,G11508,G11506,G11507);
  nand GNAME8467(G8467,G9442,G11502,G11500,G11501);
  nand GNAME8468(G8468,G9441,G11496,G11494,G11495);
  nand GNAME8469(G8469,G9440,G11490,G11488,G11489);
  nand GNAME8470(G8470,G9439,G11484,G11482,G11483);
  nand GNAME8471(G8471,G9438,G11478,G11476,G11477);
  nand GNAME8472(G8472,G9437,G11472,G11470,G11471);
  nand GNAME8473(G8473,G9436,G11466,G11464,G11465);
  nand GNAME8474(G8474,G9435,G11447,G11445,G11446);
  nand GNAME8475(G8475,G9434,G11441,G11439,G11440);
  nand GNAME8476(G8476,G9433,G11435,G11433,G11434);
  nand GNAME8477(G8477,G9432,G11429,G11427,G11428);
  nand GNAME8478(G8478,G9431,G11423,G11421,G11422);
  nand GNAME8479(G8479,G9430,G11417,G11415,G11416);
  nand GNAME8480(G8480,G9429,G11411,G11409,G11410);
  nand GNAME8481(G8481,G9428,G11405,G11403,G11404);
  nand GNAME8482(G8482,G9427,G11386,G11384,G11385);
  nand GNAME8483(G8483,G9426,G11380,G11378,G11379);
  nand GNAME8484(G8484,G9425,G11374,G11372,G11373);
  nand GNAME8485(G8485,G9424,G11368,G11366,G11367);
  nand GNAME8486(G8486,G9423,G11362,G11360,G11361);
  nand GNAME8487(G8487,G9422,G11356,G11354,G11355);
  nand GNAME8488(G8488,G9421,G11350,G11348,G11349);
  nand GNAME8489(G8489,G9420,G11344,G11342,G11343);
  nand GNAME8490(G8490,G9419,G11325,G11323,G11324);
  nand GNAME8491(G8491,G9418,G11319,G11317,G11318);
  nand GNAME8492(G8492,G9417,G11313,G11311,G11312);
  nand GNAME8493(G8493,G9416,G11307,G11305,G11306);
  nand GNAME8494(G8494,G9415,G11301,G11299,G11300);
  nand GNAME8495(G8495,G9414,G11295,G11293,G11294);
  nand GNAME8496(G8496,G9413,G11289,G11287,G11288);
  nand GNAME8497(G8497,G9412,G11283,G11281,G11282);
  nand GNAME8498(G8498,G9411,G11264,G11262,G11263);
  nand GNAME8499(G8499,G9410,G11255,G11253,G11254);
  nand GNAME8500(G8500,G9409,G11246,G11244,G11245);
  nand GNAME8501(G8501,G9408,G11237,G11235,G11236);
  nand GNAME8502(G8502,G9407,G11228,G11226,G11227);
  nand GNAME8503(G8503,G9406,G11219,G11217,G11218);
  nand GNAME8504(G8504,G9405,G11210,G11208,G11209);
  nand GNAME8505(G8505,G9404,G11201,G11199,G11200);
  and GNAME8506(G8506,G11040,G59562);
  nand GNAME8507(G8507,G11076,G11074,G11075);
  nand GNAME8508(G8508,G11069,G11067,G11068);
  nand GNAME8509(G8509,G11058,G11056,G11057);
  nand GNAME8510(G8510,G9398,G11032,G11034,G11035);
  nand GNAME8511(G8511,G9397,G11026,G11028,G11029);
  nand GNAME8512(G8512,G9396,G11020,G11022,G11023);
  nand GNAME8513(G8513,G9395,G11014,G11016,G11017);
  nand GNAME8514(G8514,G9394,G11012,G11010,G11011);
  nand GNAME8515(G8515,G9393,G11006,G11004,G11005);
  nand GNAME8516(G8516,G9392,G11000,G10998,G10999);
  nand GNAME8517(G8517,G9391,G10994,G10992,G10993);
  nand GNAME8518(G8518,G9390,G10988,G10986,G10987);
  nand GNAME8519(G8519,G9389,G10982,G10980,G10981);
  nand GNAME8520(G8520,G9388,G10976,G10974,G10975);
  nand GNAME8521(G8521,G9387,G10970,G10968,G10969);
  nand GNAME8522(G8522,G9386,G10964,G10962,G10963);
  nand GNAME8523(G8523,G9385,G10958,G10956,G10957);
  nand GNAME8524(G8524,G9384,G10952,G10950,G10951);
  nand GNAME8525(G8525,G9383,G10946,G10944,G10945);
  nand GNAME8526(G8526,G9382,G10940,G10938,G10939);
  nand GNAME8527(G8527,G9381,G10934,G10932,G10933);
  nand GNAME8528(G8528,G9380,G10928,G10926,G10927);
  nand GNAME8529(G8529,G9379,G10922,G10920,G10921);
  nand GNAME8530(G8530,G9378,G10916,G10914,G10915);
  nand GNAME8531(G8531,G9377,G10910,G10908,G10909);
  nand GNAME8532(G8532,G9376,G10904,G10902,G10903);
  nand GNAME8533(G8533,G9375,G10898,G10896,G10897);
  nand GNAME8534(G8534,G9374,G10892,G10890,G10891);
  nand GNAME8535(G8535,G9373,G10886,G10884,G10885);
  nand GNAME8536(G8536,G9372,G10880,G10878,G10879);
  nand GNAME8537(G8537,G9371,G10874,G10872,G10873);
  nand GNAME8538(G8538,G9370,G10868,G10866,G10867);
  nand GNAME8539(G8539,G9369,G10862,G10860,G10861);
  nand GNAME8540(G8540,G9368,G10856,G10854,G10855);
  nand GNAME8541(G8541,G9367,G10850,G10848,G10849);
  nand GNAME8542(G8542,G10807,G10808,G10806,G10804,G10805);
  nand GNAME8543(G8543,G10802,G10803,G10801,G10799,G10800);
  nand GNAME8544(G8544,G10797,G10798,G10796,G10794,G10795);
  nand GNAME8545(G8545,G10792,G10793,G10791,G10789,G10790);
  nand GNAME8546(G8546,G10787,G10788,G10786,G10784,G10785);
  nand GNAME8547(G8547,G10782,G10783,G10781,G10779,G10780);
  nand GNAME8548(G8548,G10777,G10778,G10776,G10774,G10775);
  nand GNAME8549(G8549,G10772,G10773,G10771,G10769,G10770);
  nand GNAME8550(G8550,G10767,G10768,G10766,G10764,G10765);
  nand GNAME8551(G8551,G10762,G10763,G10761,G10759,G10760);
  nand GNAME8552(G8552,G10757,G10758,G10756,G10754,G10755);
  nand GNAME8553(G8553,G10752,G10753,G10751,G10749,G10750);
  nand GNAME8554(G8554,G10747,G10748,G10746,G10744,G10745);
  nand GNAME8555(G8555,G10742,G10743,G10741,G10739,G10740);
  nand GNAME8556(G8556,G10737,G10738,G10736,G10734,G10735);
  nand GNAME8557(G8557,G10732,G10733,G10731,G10729,G10730);
  nand GNAME8558(G8558,G10727,G10728,G10726,G10724,G10725);
  nand GNAME8559(G8559,G10722,G10723,G10721,G10719,G10720);
  nand GNAME8560(G8560,G10717,G10718,G10716,G10714,G10715);
  nand GNAME8561(G8561,G10712,G10713,G10711,G10709,G10710);
  nand GNAME8562(G8562,G10707,G10708,G10706,G10704,G10705);
  nand GNAME8563(G8563,G10702,G10703,G10701,G10699,G10700);
  nand GNAME8564(G8564,G10697,G10698,G10696,G10694,G10695);
  nand GNAME8565(G8565,G10692,G10693,G10691,G10689,G10690);
  nand GNAME8566(G8566,G10687,G10688,G10686,G10684,G10685);
  nand GNAME8567(G8567,G10682,G10683,G10681,G10679,G10680);
  nand GNAME8568(G8568,G10677,G10678,G10676,G10674,G10675);
  nand GNAME8569(G8569,G10672,G10673,G10671,G10669,G10670);
  nand GNAME8570(G8570,G10667,G10668,G10666,G10664,G10665);
  nand GNAME8571(G8571,G10662,G10663,G10661,G10659,G10660);
  nand GNAME8572(G8572,G10657,G10658,G10656,G10654,G10655);
  nand GNAME8573(G8573,G10652,G10653,G10651,G10649,G10650);
  nand GNAME8574(G8574,G10647,G10645,G10646);
  nand GNAME8575(G8575,G10644,G10642,G10643);
  nand GNAME8576(G8576,G10641,G10639,G10640);
  nand GNAME8577(G8577,G10638,G10636,G10637);
  nand GNAME8578(G8578,G10635,G10633,G10634);
  nand GNAME8579(G8579,G10632,G10630,G10631);
  nand GNAME8580(G8580,G10629,G10627,G10628);
  nand GNAME8581(G8581,G10626,G10624,G10625);
  nand GNAME8582(G8582,G10623,G10621,G10622);
  nand GNAME8583(G8583,G10620,G10618,G10619);
  nand GNAME8584(G8584,G10617,G10615,G10616);
  nand GNAME8585(G8585,G10614,G10612,G10613);
  nand GNAME8586(G8586,G10611,G10609,G10610);
  nand GNAME8587(G8587,G10608,G10606,G10607);
  nand GNAME8588(G8588,G10605,G10603,G10604);
  nand GNAME8589(G8589,G10602,G10600,G10601);
  nand GNAME8590(G8590,G10599,G10598,G10642);
  nand GNAME8591(G8591,G10597,G10596,G10639);
  nand GNAME8592(G8592,G10595,G10594,G10636);
  nand GNAME8593(G8593,G10593,G10592,G10633);
  nand GNAME8594(G8594,G10591,G10590,G10630);
  nand GNAME8595(G8595,G10589,G10588,G10627);
  nand GNAME8596(G8596,G10587,G10586,G10624);
  nand GNAME8597(G8597,G10623,G10584,G10585);
  nand GNAME8598(G8598,G10620,G10582,G10583);
  nand GNAME8599(G8599,G10617,G10580,G10581);
  nand GNAME8600(G8600,G10614,G10578,G10579);
  nand GNAME8601(G8601,G10611,G10576,G10577);
  nand GNAME8602(G8602,G10608,G10574,G10575);
  nand GNAME8603(G8603,G10605,G10572,G10573);
  nand GNAME8604(G8604,G10602,G10570,G10571);
  nand GNAME8605(G8605,G10567,G10565,G10566);
  nand GNAME8606(G8606,G10564,G10562,G10563);
  nand GNAME8607(G8607,G10561,G10559,G10560);
  nand GNAME8608(G8608,G10558,G10556,G10557);
  nand GNAME8609(G8609,G10555,G10553,G10554);
  nand GNAME8610(G8610,G10552,G10550,G10551);
  nand GNAME8611(G8611,G10549,G10547,G10548);
  nand GNAME8612(G8612,G10546,G10544,G10545);
  nand GNAME8613(G8613,G10543,G10541,G10542);
  nand GNAME8614(G8614,G10540,G10538,G10539);
  nand GNAME8615(G8615,G10537,G10535,G10536);
  nand GNAME8616(G8616,G10534,G10532,G10533);
  nand GNAME8617(G8617,G10531,G10529,G10530);
  nand GNAME8618(G8618,G10528,G10526,G10527);
  nand GNAME8619(G8619,G10525,G10523,G10524);
  nand GNAME8620(G8620,G10522,G10520,G10521);
  nand GNAME8621(G8621,G10519,G10517,G10518);
  nand GNAME8622(G8622,G10516,G10514,G10515);
  nand GNAME8623(G8623,G10513,G10511,G10512);
  nand GNAME8624(G8624,G10510,G10508,G10509);
  nand GNAME8625(G8625,G10507,G10505,G10506);
  nand GNAME8626(G8626,G10504,G10502,G10503);
  nand GNAME8627(G8627,G10501,G10499,G10500);
  nand GNAME8628(G8628,G10498,G10496,G10497);
  nand GNAME8629(G8629,G10495,G10493,G10494);
  nand GNAME8630(G8630,G10492,G10490,G10491);
  nand GNAME8631(G8631,G10489,G10487,G10488);
  nand GNAME8632(G8632,G10486,G10484,G10485);
  nand GNAME8633(G8633,G10483,G10481,G10482);
  nand GNAME8634(G8634,G10480,G10478,G10479);
  nand GNAME8635(G8635,G10477,G10475,G10476);
  and GNAME8636(G8636,G8873,G59693);
  nand GNAME8637(G8637,G10466,G10467,G10468,G10469);
  nand GNAME8638(G8638,G10462,G10463,G10464,G10465);
  nand GNAME8639(G8639,G10458,G10459,G10460,G10461);
  nand GNAME8640(G8640,G10454,G10455,G10456,G10457);
  nand GNAME8641(G8641,G10450,G10451,G10452,G10453);
  nand GNAME8642(G8642,G10446,G10447,G10448,G10449);
  nand GNAME8643(G8643,G10442,G10443,G10444,G10445);
  nand GNAME8644(G8644,G10438,G10439,G10440,G10441);
  nand GNAME8645(G8645,G10434,G10435,G10436,G10437);
  nand GNAME8646(G8646,G10430,G10431,G10432,G10433);
  nand GNAME8647(G8647,G10426,G10427,G10428,G10429);
  nand GNAME8648(G8648,G10422,G10423,G10424,G10425);
  nand GNAME8649(G8649,G10418,G10419,G10420,G10421);
  nand GNAME8650(G8650,G10414,G10415,G10416,G10417);
  nand GNAME8651(G8651,G10410,G10411,G10412,G10413);
  nand GNAME8652(G8652,G10406,G10407,G10408,G10409);
  nand GNAME8653(G8653,G10404,G10405,G10403,G10401,G10402);
  nand GNAME8654(G8654,G10399,G10400,G10398,G10396,G10397);
  nand GNAME8655(G8655,G10394,G10395,G10393,G10391,G10392);
  nand GNAME8656(G8656,G10389,G10390,G10388,G10386,G10387);
  nand GNAME8657(G8657,G10384,G10385,G10383,G10381,G10382);
  nand GNAME8658(G8658,G10379,G10380,G10378,G10376,G10377);
  nand GNAME8659(G8659,G10374,G10375,G10373,G10371,G10372);
  nand GNAME8660(G8660,G10369,G10370,G10368,G10366,G10367);
  nand GNAME8661(G8661,G10364,G10365,G10363,G10361,G10362);
  nand GNAME8662(G8662,G10359,G10360,G10358,G10356,G10357);
  nand GNAME8663(G8663,G10354,G10355,G10353,G10351,G10352);
  nand GNAME8664(G8664,G10349,G10350,G10348,G10346,G10347);
  nand GNAME8665(G8665,G10344,G10345,G10343,G10341,G10342);
  nand GNAME8666(G8666,G10339,G10340,G10338,G10336,G10337);
  nand GNAME8667(G8667,G10334,G10335,G10333,G10331,G10332);
  nand GNAME8668(G8668,G10330,G10328,G10329);
  nand GNAME8669(G8669,G10318,G10316,G10317);
  nand GNAME8670(G8670,G10315,G10313,G10314);
  nand GNAME8671(G8671,G10312,G10310,G10311);
  nand GNAME8672(G8672,G10309,G10307,G10308);
  nand GNAME8673(G8673,G10306,G10304,G10305);
  nand GNAME8674(G8674,G10303,G10301,G10302);
  nand GNAME8675(G8675,G10300,G10298,G10299);
  nand GNAME8676(G8676,G10297,G10295,G10296);
  nand GNAME8677(G8677,G10294,G10292,G10293);
  nand GNAME8678(G8678,G10291,G10289,G10290);
  nand GNAME8679(G8679,G10288,G10286,G10287);
  nand GNAME8680(G8680,G10285,G10283,G10284);
  nand GNAME8681(G8681,G10282,G10280,G10281);
  nand GNAME8682(G8682,G10279,G10277,G10278);
  nand GNAME8683(G8683,G10276,G10274,G10275);
  nand GNAME8684(G8684,G10273,G10271,G10272);
  nand GNAME8685(G8685,G10270,G10268,G10269);
  nand GNAME8686(G8686,G10267,G10265,G10266);
  nand GNAME8687(G8687,G10264,G10262,G10263);
  nand GNAME8688(G8688,G10261,G10259,G10260);
  nand GNAME8689(G8689,G10258,G10256,G10257);
  nand GNAME8690(G8690,G10255,G10253,G10254);
  nand GNAME8691(G8691,G10252,G10250,G10251);
  nand GNAME8692(G8692,G10249,G10247,G10248);
  nand GNAME8693(G8693,G10246,G10244,G10245);
  nand GNAME8694(G8694,G10243,G10241,G10242);
  nand GNAME8695(G8695,G10240,G10238,G10239);
  nand GNAME8696(G8696,G10237,G10235,G10236);
  nand GNAME8697(G8697,G10234,G10232,G10233);
  nand GNAME8698(G8698,G10231,G10229,G10230);
  nand GNAME8699(G8699,G10228,G10226,G10227);
  nand GNAME8700(G8700,G10224,G10225);
  nand GNAME8701(G8701,G9362,G10215,G10217,G10218);
  nand GNAME8702(G8702,G9361,G10209,G10211,G10212);
  nand GNAME8703(G8703,G10207,G9360,G10204,G10202,G10203);
  nand GNAME8704(G8704,G10201,G9359,G10198,G10196,G10197);
  nand GNAME8705(G8705,G9358,G10191,G10193,G10194);
  nand GNAME8706(G8706,G9357,G10185,G10187,G10188);
  nand GNAME8707(G8707,G9356,G10177,G10174,G10175,G10176);
  nand GNAME8708(G8708,G9355,G10171,G10168,G10169,G10170);
  nand GNAME8709(G8709,G9354,G10165,G10162,G10163,G10164);
  nand GNAME8710(G8710,G9353,G10159,G10156,G10157,G10160);
  nand GNAME8711(G8711,G9352,G10154,G10150,G10151,G10152);
  nand GNAME8712(G8712,G9351,G10148,G10144,G10145,G10146);
  nand GNAME8713(G8713,G9350,G10142,G10138,G10139,G10140);
  nand GNAME8714(G8714,G9349,G10136,G10132,G10133,G10134);
  nand GNAME8715(G8715,G9348,G10130,G10126,G10127,G10128);
  nand GNAME8716(G8716,G9347,G10124,G10120,G10121,G10122);
  nand GNAME8717(G8717,G9346,G10118,G10114,G10115,G10116);
  nand GNAME8718(G8718,G9345,G10112,G10108,G10109,G10110);
  nand GNAME8719(G8719,G9344,G10106,G10102,G10103,G10104);
  nand GNAME8720(G8720,G9343,G10100,G10096,G10097,G10098);
  nand GNAME8721(G8721,G9342,G10093,G10089,G10090);
  nand GNAME8722(G8722,G9341,G10087,G10083,G10084);
  nand GNAME8723(G8723,G9340,G10081,G10077,G10078);
  nand GNAME8724(G8724,G9339,G10075,G10071,G10072);
  nand GNAME8725(G8725,G9338,G10069,G10065,G10066);
  nand GNAME8726(G8726,G9337,G10063,G10059,G10060);
  nand GNAME8727(G8727,G9336,G10057,G10053,G10054);
  nand GNAME8728(G8728,G9335,G10051,G10047,G10048);
  nand GNAME8729(G8729,G9334,G10045,G10041,G10042);
  nand GNAME8730(G8730,G9333,G10039,G10035,G10036);
  nand GNAME8731(G8731,G9332,G10033,G10029,G10030);
  nand GNAME8732(G8732,G9331,G10027,G10023,G10024);
  nand GNAME8733(G8733,G10011,G9808,G8831);
  nand GNAME8734(G8734,G10010,G10008,G10009);
  nand GNAME8735(G8735,G10006,G9808,G8832);
  nand GNAME8736(G8736,G8832,G13850,G13851);
  nand GNAME8737(G8737,G10004,G10003);
  nand GNAME8738(G8738,G10001,G10002);
  nand GNAME8739(G8739,G9814,G13843,G13844);
  nand GNAME8740(G8740,G9814,G13839,G13840);
  nand GNAME8741(G8741,G9970,G9971);
  nand GNAME8742(G8742,G9962,G9961);
  and GNAME8743(G8743,G8780,G9849);
  nand GNAME8744(G8744,G13860,G13861,G11047,G11048);
  and GNAME8745(G8745,G8796,G9832);
  nand GNAME8746(G8746,G9299,G9300,G9301,G9302);
  and GNAME8747(G8747,G12184,G9104);
  not GNAME8748(G8748,G33);
  not GNAME8749(G8749,G1588);
  nand GNAME8750(G8750,G8891,G9832,G9849);
  not GNAME8751(G8751,G59426);
  not GNAME8752(G8752,G59561);
  and GNAME8753(G8753,G8768,G8761);
  and GNAME8754(G8754,G8756,G59561);
  and GNAME8755(G8755,G8753,G8754);
  not GNAME8756(G8756,G59560);
  and GNAME8757(G8757,G8752,G59560);
  and GNAME8758(G8758,G8753,G8757);
  and GNAME8759(G8759,G59561,G59560);
  and GNAME8760(G8760,G8753,G8759);
  not GNAME8761(G8761,G59559);
  nor GNAME8762(G8762,G59558,G8761);
  nor GNAME8763(G8763,G59561,G59560);
  and GNAME8764(G8764,G8762,G8763);
  and GNAME8765(G8765,G8754,G8762);
  and GNAME8766(G8766,G8757,G8762);
  and GNAME8767(G8767,G8759,G8762);
  not GNAME8768(G8768,G59558);
  and GNAME8769(G8769,G8761,G59558);
  and GNAME8770(G8770,G8763,G8769);
  and GNAME8771(G8771,G8754,G8769);
  and GNAME8772(G8772,G8757,G8769);
  nor GNAME8773(G8773,G9787,G9788);
  nor GNAME8774(G8774,G8761,G8768);
  and GNAME8775(G8775,G8763,G8774);
  and GNAME8776(G8776,G8754,G8774);
  and GNAME8777(G8777,G8757,G8774);
  and GNAME8778(G8778,G8759,G8774);
  and GNAME8779(G8779,G8753,G8763);
  nand GNAME8780(G8780,G9315,G9316,G9317,G9318);
  nand GNAME8781(G8781,G9319,G9320,G9321,G9322);
  nand GNAME8782(G8782,G9303,G9304,G9305,G9306);
  nand GNAME8783(G8783,G9307,G9308,G9309,G9310);
  and GNAME8784(G8784,G9917,G9900);
  and GNAME8785(G8785,G9883,G8745,G8792);
  and GNAME8786(G8786,G8852,G8746,G8784,G8785);
  not GNAME8787(G8787,G59428);
  and GNAME8788(G8788,G8786,G59428);
  not GNAME8789(G8789,G22263);
  and GNAME8790(G8790,G8814,G59426);
  nor GNAME8791(G8791,G9832,G8783);
  nand GNAME8792(G8792,G9291,G9292,G9293,G9294);
  and GNAME8793(G8793,G8791,G8782,G8852);
  nand GNAME8794(G8794,G8781,G9951,G9866,G8793);
  nor GNAME8795(G8795,G59427,G8787);
  nand GNAME8796(G8796,G9311,G9312,G9313,G9314);
  nor GNAME8797(G8797,G8782,G8796);
  nor GNAME8798(G8798,G8781,G9934,G9951);
  nand GNAME8799(G8799,G8797,G8798,G9900,G8792,G9832);
  and GNAME8800(G8800,G59428,G8790);
  not GNAME8801(G8801,G21598);
  and GNAME8802(G8802,G8814,G8751);
  nand GNAME8803(G8803,G8878,G9957);
  not GNAME8804(G8804,G59391);
  nand GNAME8805(G8805,G8817,G59391);
  not GNAME8806(G8806,G59392);
  or GNAME8807(G8807,G9960,G8812);
  and GNAME8808(G8808,G9964,G9805,G8852);
  and GNAME8809(G8809,G9803,G9967,G9968,G8808);
  and GNAME8810(G8810,G8834,G8802);
  and GNAME8811(G8811,G8806,G59391);
  and GNAME8812(G8812,G8804,G8806);
  and GNAME8813(G8813,G8787,G59426);
  not GNAME8814(G8814,G59427);
  nand GNAME8815(G8815,G8813,G59427);
  nor GNAME8816(G8816,G8907,G59425);
  not GNAME8817(G8817,G59390);
  nand GNAME8818(G8818,G9976,G8806);
  not GNAME8819(G8819,G59797);
  and GNAME8820(G8820,G59426,G9849);
  and GNAME8821(G8821,G9883,G8793);
  and GNAME8822(G8822,G8821,G8792,G8746);
  and GNAME8823(G8823,G8852,G9917);
  and GNAME8824(G8824,G8746,G9866);
  and GNAME8825(G8825,G8823,G8824,G9883,G8743,G8783);
  and GNAME8826(G8826,G8792,G8783);
  and GNAME8827(G8827,G8796,G9917);
  and GNAME8828(G8828,G8780,G8798,G8826,G8827);
  and GNAME8829(G8829,G9324,G9326,G9328,G9330);
  not GNAME8830(G8830,G59758);
  or GNAME8831(G8831,G13985,G59759,G59394);
  nand GNAME8832(G8832,G8829,G59759);
  and GNAME8833(G8833,G8819,G59427);
  not GNAME8834(G8834,G59425);
  and GNAME8835(G8835,G8749,G8819);
  nor GNAME8836(G8836,G10012,G8751);
  and GNAME8837(G8837,G10022,G8836);
  not GNAME8838(G8838,G9282);
  nor GNAME8839(G8839,G59426,G8787);
  and GNAME8840(G8840,G8842,G8839);
  and GNAME8841(G8841,G8797,G9977,G8835,G8836);
  nand GNAME8842(G8842,G9811,G9812,G10828,G13980);
  nand GNAME8843(G8843,G10014,G10015);
  not GNAME8844(G8844,G21670);
  not GNAME8845(G8845,G21997);
  not GNAME8846(G8846,G21631);
  not GNAME8847(G8847,G21936);
  not GNAME8848(G8848,G21723);
  not GNAME8849(G8849,G22042);
  not GNAME8850(G8850,G21699);
  not GNAME8851(G8851,G21995);
  nand GNAME8852(G8852,G9295,G9296,G9297,G9298);
  and GNAME8853(G8853,G9951,G9883);
  nor GNAME8854(G8854,G9805,G8783,G8852);
  nand GNAME8855(G8855,G8745,G8792,G8782,G8854);
  and GNAME8856(G8856,G59428,G8828);
  nand GNAME8857(G8857,G10223,G8790);
  nor GNAME8858(G8858,G8746,G8857);
  nor GNAME8859(G8859,G9951,G8857);
  and GNAME8860(G8860,G8782,G9832);
  nand GNAME8861(G8861,G9866,G9849,G8854,G8860);
  and GNAME8862(G8862,G13986,G9849);
  nand GNAME8863(G8863,G59428,G8862);
  and GNAME8864(G8864,G59428,G8825);
  nand GNAME8865(G8865,G10327,G8790);
  nor GNAME8866(G8866,G9805,G8865);
  nor GNAME8867(G8867,G9883,G8865);
  nor GNAME8868(G8868,G9866,G8865);
  nor GNAME8869(G8869,G9789,G8865);
  nor GNAME8870(G8870,G8887,G8865);
  and GNAME8871(G8871,G8796,G13986);
  nand GNAME8872(G8872,G9955,G9976,G59428);
  and GNAME8873(G8873,G8815,G10474);
  nor GNAME8874(G8874,G8873,G59428);
  nor GNAME8875(G8875,G8873,G8787);
  and GNAME8876(G8876,G8792,G8875);
  nand GNAME8877(G8877,G9955,G8800);
  nand GNAME8878(G8878,G8790,G8788,G22263);
  and GNAME8879(G8879,G10568,G10569);
  nor GNAME8880(G8880,G8879,G8796);
  nor GNAME8881(G8881,G8879,G9849);
  and GNAME8882(G8882,G10003,G10648);
  nor GNAME8883(G8883,G9243,G8882);
  nor GNAME8884(G8884,G8882,G9796);
  nor GNAME8885(G8885,G8882,G8787);
  nor GNAME8886(G8886,G8882,G9797);
  and GNAME8887(G8887,G9883,G9866);
  and GNAME8888(G8888,G9363,G8808,G10813,G10814);
  nor GNAME8889(G8889,G8906,G8751);
  and GNAME8890(G8890,G8825,G8889);
  nor GNAME8891(G8891,G9805,G9934,G8792);
  and GNAME8892(G8892,G10809,G13852,G13853);
  and GNAME8893(G8893,G10810,G10834);
  and GNAME8894(G8894,G8796,G9866);
  and GNAME8895(G8895,G9365,G8893,G10839,G8892);
  and GNAME8896(G8896,G9364,G9934,G9900,G8797);
  and GNAME8897(G8897,G8791,G8894,G9951,G8781,G8782);
  and GNAME8898(G8898,G10842,G10843);
  and GNAME8899(G8899,G8855,G8898);
  and GNAME8900(G8900,G9366,G8799,G8895);
  and GNAME8901(G8901,G10844,G8889);
  and GNAME8902(G8902,G11100,G10470);
  and GNAME8903(G8903,G10832,G8889);
  and GNAME8904(G8904,G10829,G8889);
  nor GNAME8905(G8905,G59426,G8906);
  and GNAME8906(G8906,G10827,G10828);
  and GNAME8907(G8907,G59426,G59427);
  and GNAME8908(G8908,G59428,G8907);
  nand GNAME8909(G8909,G8787,G59425);
  nand GNAME8910(G8910,G11037,G13858,G13859);
  not GNAME8911(G8911,G59566);
  nor GNAME8912(G8912,G8932,G11042,G8751,G8787);
  and GNAME8913(G8913,G13865,G13866,G9794,G11041);
  nand GNAME8914(G8914,G11043,G8919);
  nor GNAME8915(G8915,G9796,G59426,G11040);
  and GNAME8916(G8916,G8917,G11046);
  nand GNAME8917(G8917,G11038,G9813,G11039);
  not GNAME8918(G8918,G59565);
  or GNAME8919(G8919,G8913,G8912);
  nand GNAME8920(G8920,G11049,G11050);
  nand GNAME8921(G8921,G11054,G11052,G11053);
  not GNAME8922(G8922,G59564);
  and GNAME8923(G8923,G59566,G59565);
  and GNAME8924(G8924,G11061,G11059,G11060);
  nand GNAME8925(G8925,G11063,G11064);
  nand GNAME8926(G8926,G11065,G9772);
  nor GNAME8927(G8927,G59563,G8922);
  not GNAME8928(G8928,G59563);
  nor GNAME8929(G8929,G59426,G8801);
  nand GNAME8930(G8930,G11089,G59561);
  nand GNAME8931(G8931,G11095,G8933);
  and GNAME8932(G8932,G13864,G59427);
  nand GNAME8933(G8933,G11092,G11093);
  nand GNAME8934(G8934,G11117,G11118);
  nand GNAME8935(G8935,G11139,G11140);
  nand GNAME8936(G8936,G11136,G11137);
  nand GNAME8937(G8937,G11142,G9777);
  nand GNAME8938(G8938,G11171,G13901,G13902);
  nand GNAME8939(G8939,G11166,G11168);
  and GNAME8940(G8940,G59427,G59797);
  nand GNAME8941(G8941,G11164,G11159);
  nor GNAME8942(G8942,G13886,G8941);
  nor GNAME8943(G8943,G11096,G13892);
  nor GNAME8944(G8944,G11038,G9795);
  nor GNAME8945(G8945,G13879,G9250);
  nor GNAME8946(G8946,G11066,G11044);
  nand GNAME8947(G8947,G8945,G8946);
  nor GNAME8948(G8948,G8960,G13983);
  and GNAME8949(G8949,G11186,G8948);
  nor GNAME8950(G8950,G59564,G59563);
  nor GNAME8951(G8951,G59565,G59566);
  or GNAME8952(G8952,G8982,G8993);
  or GNAME8953(G8953,G11070,G9038,G9045);
  nor GNAME8954(G8954,G9251,G8953);
  nor GNAME8955(G8955,G8911,G8952);
  and GNAME8956(G8956,G8954,G8955);
  and GNAME8957(G8957,G8950,G8951);
  nor GNAME8958(G8958,G8956,G11191);
  and GNAME8959(G8959,G8910,G1659);
  and GNAME8960(G8960,G8942,G8943);
  and GNAME8961(G8961,G1643,G8944);
  nor GNAME8962(G8962,G11038,G9797);
  and GNAME8963(G8963,G8910,G1648);
  and GNAME8964(G8964,G1642,G8944);
  and GNAME8965(G8965,G8910,G1637);
  and GNAME8966(G8966,G1641,G8944);
  and GNAME8967(G8967,G8910,G1634);
  and GNAME8968(G8968,G1640,G8944);
  and GNAME8969(G8969,G8910,G1633);
  and GNAME8970(G8970,G1639,G8944);
  and GNAME8971(G8971,G8910,G1632);
  and GNAME8972(G8972,G1638,G8944);
  and GNAME8973(G8973,G8910,G1631);
  and GNAME8974(G8974,G1636,G8944);
  and GNAME8975(G8975,G8910,G1630);
  and GNAME8976(G8976,G1635,G8944);
  nor GNAME8977(G8977,G13892,G8931);
  nor GNAME8978(G8978,G11066,G8914);
  nand GNAME8979(G8979,G8945,G8978);
  nor GNAME8980(G8980,G8987,G13983);
  and GNAME8981(G8981,G11268,G8980);
  and GNAME8982(G8982,G8918,G59566);
  nor GNAME8983(G8983,G59566,G8952);
  and GNAME8984(G8984,G8954,G8983);
  and GNAME8985(G8985,G8950,G8982);
  nor GNAME8986(G8986,G8984,G11273);
  and GNAME8987(G8987,G8942,G8977);
  nor GNAME8988(G8988,G9253,G8941);
  nor GNAME8989(G8989,G13873,G13879);
  nand GNAME8990(G8990,G8946,G8989);
  nor GNAME8991(G8991,G8998,G13983);
  and GNAME8992(G8992,G11329,G8991);
  and GNAME8993(G8993,G8911,G59565);
  and GNAME8994(G8994,G8952,G59566);
  and GNAME8995(G8995,G8954,G8994);
  and GNAME8996(G8996,G8950,G8993);
  nor GNAME8997(G8997,G8995,G11334);
  and GNAME8998(G8998,G8943,G8988);
  nand GNAME8999(G8999,G8978,G8989);
  nor GNAME9000(G9000,G9006,G13983);
  and GNAME9001(G9001,G11390,G9000);
  and GNAME9002(G9002,G8952,G8911);
  and GNAME9003(G9003,G8954,G9002);
  and GNAME9004(G9004,G8923,G8950);
  nor GNAME9005(G9005,G9003,G11395);
  and GNAME9006(G9006,G8977,G8988);
  nor GNAME9007(G9007,G11096,G9264);
  nor GNAME9008(G9008,G11044,G8926);
  nand GNAME9009(G9009,G8945,G9008);
  nor GNAME9010(G9010,G9016,G13983);
  and GNAME9011(G9011,G11451,G9010);
  nor GNAME9012(G9012,G13876,G8953);
  and GNAME9013(G9013,G8955,G9012);
  and GNAME9014(G9014,G8927,G8951);
  nor GNAME9015(G9015,G9013,G11456);
  and GNAME9016(G9016,G8942,G9007);
  nor GNAME9017(G9017,G8931,G9264);
  nor GNAME9018(G9018,G8914,G8926);
  nand GNAME9019(G9019,G8945,G9018);
  nor GNAME9020(G9020,G9025,G13983);
  and GNAME9021(G9021,G11512,G9020);
  and GNAME9022(G9022,G8983,G9012);
  and GNAME9023(G9023,G8927,G8982);
  nor GNAME9024(G9024,G9022,G11517);
  and GNAME9025(G9025,G8942,G9017);
  nand GNAME9026(G9026,G8989,G9008);
  nor GNAME9027(G9027,G9032,G13983);
  and GNAME9028(G9028,G11573,G9027);
  and GNAME9029(G9029,G8994,G9012);
  and GNAME9030(G9030,G8927,G8993);
  nor GNAME9031(G9031,G9029,G11578);
  and GNAME9032(G9032,G8988,G9007);
  nand GNAME9033(G9033,G8989,G9018);
  nor GNAME9034(G9034,G9039,G13983);
  and GNAME9035(G9035,G11634,G9034);
  and GNAME9036(G9036,G9002,G9012);
  nor GNAME9037(G9037,G9036,G11639);
  and GNAME9038(G9038,G8923,G8927);
  and GNAME9039(G9039,G8988,G9017);
  nor GNAME9040(G9040,G11165,G13886);
  nor GNAME9041(G9041,G9252,G9250);
  nand GNAME9042(G9042,G8946,G9041);
  nor GNAME9043(G9043,G9050,G13983);
  and GNAME9044(G9044,G11695,G9043);
  and GNAME9045(G9045,G8922,G59563);
  and GNAME9046(G9046,G8953,G13876);
  and GNAME9047(G9047,G8955,G9046);
  and GNAME9048(G9048,G8951,G9045);
  nor GNAME9049(G9049,G9047,G11700);
  and GNAME9050(G9050,G8943,G9040);
  nand GNAME9051(G9051,G8978,G9041);
  nor GNAME9052(G9052,G9057,G13983);
  and GNAME9053(G9053,G11756,G9052);
  and GNAME9054(G9054,G8983,G9046);
  and GNAME9055(G9055,G8982,G9045);
  nor GNAME9056(G9056,G9054,G11761);
  and GNAME9057(G9057,G8977,G9040);
  nor GNAME9058(G9058,G11165,G9253);
  nor GNAME9059(G9059,G13873,G9252);
  nand GNAME9060(G9060,G8946,G9059);
  nor GNAME9061(G9061,G9066,G13983);
  and GNAME9062(G9062,G11817,G9061);
  and GNAME9063(G9063,G8994,G9046);
  and GNAME9064(G9064,G8993,G9045);
  nor GNAME9065(G9065,G9063,G11822);
  and GNAME9066(G9066,G8943,G9058);
  nand GNAME9067(G9067,G8978,G9059);
  nor GNAME9068(G9068,G9073,G13983);
  and GNAME9069(G9069,G11878,G9068);
  and GNAME9070(G9070,G9002,G9046);
  and GNAME9071(G9071,G8923,G9045);
  nor GNAME9072(G9072,G9070,G11883);
  and GNAME9073(G9073,G8977,G9058);
  nand GNAME9074(G9074,G9008,G9041);
  nor GNAME9075(G9075,G9082,G13983);
  and GNAME9076(G9076,G11939,G9075);
  nor GNAME9077(G9077,G8922,G8928);
  and GNAME9078(G9078,G8953,G9251);
  and GNAME9079(G9079,G8955,G9078);
  and GNAME9080(G9080,G8951,G9077);
  nor GNAME9081(G9081,G9079,G11944);
  and GNAME9082(G9082,G9007,G9040);
  nand GNAME9083(G9083,G9018,G9041);
  nor GNAME9084(G9084,G9089,G13983);
  and GNAME9085(G9085,G12000,G9084);
  and GNAME9086(G9086,G8983,G9078);
  and GNAME9087(G9087,G8982,G9077);
  nor GNAME9088(G9088,G9086,G12005);
  and GNAME9089(G9089,G9017,G9040);
  nand GNAME9090(G9090,G9008,G9059);
  nor GNAME9091(G9091,G9096,G13983);
  and GNAME9092(G9092,G12061,G9091);
  and GNAME9093(G9093,G8994,G9078);
  and GNAME9094(G9094,G8993,G9077);
  nor GNAME9095(G9095,G9093,G12066);
  and GNAME9096(G9096,G9007,G9058);
  nand GNAME9097(G9097,G9018,G9059);
  nor GNAME9098(G9098,G9103,G13983);
  and GNAME9099(G9099,G12122,G9098);
  and GNAME9100(G9100,G9002,G9078);
  nor GNAME9101(G9101,G9100,G12127);
  and GNAME9102(G9102,G8923,G9077);
  and GNAME9103(G9103,G9017,G9058);
  and GNAME9104(G9104,G9989,G8809);
  and GNAME9105(G9105,G9793,G9792);
  nor GNAME9106(G9106,G9532,G8747,G22274,G8822);
  nand GNAME9107(G9107,G13907,G13908,G12189,G59426);
  nor GNAME9108(G9108,G59427,G59425);
  not GNAME9109(G9109,G34);
  nand GNAME9110(G9110,G12205,G59390);
  and GNAME9111(G9111,G8817,G8811);
  and GNAME9112(G9112,G8811,G59390);
  nor GNAME9113(G9113,G22042,G21936);
  nor GNAME9114(G9114,G21997,G8851);
  and GNAME9115(G9115,G9113,G9114);
  nor GNAME9116(G9116,G21936,G8849);
  nor GNAME9117(G9117,G21995,G21997);
  and GNAME9118(G9118,G9116,G9117);
  and GNAME9119(G9119,G9114,G9116);
  nor GNAME9120(G9120,G22042,G8847);
  and GNAME9121(G9121,G9117,G9120);
  and GNAME9122(G9122,G9114,G9120);
  nor GNAME9123(G9123,G8847,G8849);
  and GNAME9124(G9124,G9117,G9123);
  and GNAME9125(G9125,G9114,G9123);
  nor GNAME9126(G9126,G21995,G8845);
  and GNAME9127(G9127,G9113,G9126);
  nor GNAME9128(G9128,G8845,G8851);
  and GNAME9129(G9129,G9113,G9128);
  and GNAME9130(G9130,G9116,G9126);
  and GNAME9131(G9131,G9116,G9128);
  and GNAME9132(G9132,G9120,G9126);
  and GNAME9133(G9133,G9120,G9128);
  and GNAME9134(G9134,G9123,G9126);
  and GNAME9135(G9135,G9123,G9128);
  and GNAME9136(G9136,G9113,G9117);
  nand GNAME9137(G9137,G9788,G13930,G13931);
  nor GNAME9138(G9138,G9256,G9137);
  and GNAME9139(G9139,G8759,G9138);
  and GNAME9140(G9140,G8763,G9138);
  and GNAME9141(G9141,G8754,G9138);
  nor GNAME9142(G9142,G13929,G9137);
  and GNAME9143(G9143,G8757,G9142);
  and GNAME9144(G9144,G8759,G9142);
  and GNAME9145(G9145,G8763,G9142);
  and GNAME9146(G9146,G8754,G9142);
  nor GNAME9147(G9147,G12434,G9256);
  and GNAME9148(G9148,G8757,G9147);
  and GNAME9149(G9149,G8759,G9147);
  and GNAME9150(G9150,G8763,G9147);
  and GNAME9151(G9151,G8754,G9147);
  nor GNAME9152(G9152,G12434,G13929);
  and GNAME9153(G9153,G8757,G9152);
  and GNAME9154(G9154,G8759,G9152);
  and GNAME9155(G9155,G8763,G9152);
  and GNAME9156(G9156,G8754,G9152);
  and GNAME9157(G9157,G8757,G9138);
  nor GNAME9158(G9158,G9806,G13898);
  nor GNAME9159(G9159,G11122,G8752);
  and GNAME9160(G9160,G9158,G9159);
  nand GNAME9161(G9161,G11121,G59560);
  nor GNAME9162(G9162,G59561,G9161);
  and GNAME9163(G9163,G9158,G9162);
  nor GNAME9164(G9164,G8752,G9161);
  and GNAME9165(G9165,G9158,G9164);
  nor GNAME9166(G9166,G9806,G9254);
  nor GNAME9167(G9167,G59561,G11122);
  and GNAME9168(G9168,G9166,G9167);
  and GNAME9169(G9169,G9159,G9166);
  and GNAME9170(G9170,G9162,G9166);
  and GNAME9171(G9171,G9164,G9166);
  nor GNAME9172(G9172,G13898,G8939);
  and GNAME9173(G9173,G9167,G9172);
  and GNAME9174(G9174,G9159,G9172);
  and GNAME9175(G9175,G9162,G9172);
  and GNAME9176(G9176,G9164,G9172);
  nor GNAME9177(G9177,G9254,G8939);
  and GNAME9178(G9178,G9167,G9177);
  and GNAME9179(G9179,G9159,G9177);
  and GNAME9180(G9180,G9162,G9177);
  and GNAME9181(G9181,G9164,G9177);
  and GNAME9182(G9182,G9158,G9167);
  nor GNAME9183(G9183,G21598,G9849);
  and GNAME9184(G9184,G8791,G9183);
  nand GNAME9185(G9185,G9832,G8792,G9976);
  nor GNAME9186(G9186,G8796,G9185);
  or GNAME9187(G9187,G8754,G8757);
  nor GNAME9188(G9188,G11172,G9187);
  nor GNAME9189(G9189,G59561,G11143);
  and GNAME9190(G9190,G9188,G9189);
  nor GNAME9191(G9191,G11120,G11172);
  nor GNAME9192(G9192,G11143,G8752);
  and GNAME9193(G9193,G9191,G9192);
  and GNAME9194(G9194,G9189,G9191);
  nor GNAME9195(G9195,G8752,G8937);
  and GNAME9196(G9196,G9188,G9195);
  nor GNAME9197(G9197,G59561,G8937);
  and GNAME9198(G9198,G9188,G9197);
  and GNAME9199(G9199,G9191,G9195);
  and GNAME9200(G9200,G9191,G9197);
  nor GNAME9201(G9201,G8938,G9187);
  and GNAME9202(G9202,G9192,G9201);
  and GNAME9203(G9203,G9189,G9201);
  nor GNAME9204(G9204,G11120,G8938);
  and GNAME9205(G9205,G9192,G9204);
  and GNAME9206(G9206,G9189,G9204);
  and GNAME9207(G9207,G9195,G9201);
  and GNAME9208(G9208,G9197,G9201);
  and GNAME9209(G9209,G9195,G9204);
  and GNAME9210(G9210,G9197,G9204);
  and GNAME9211(G9211,G9188,G9192);
  nor GNAME9212(G9212,G21631,G21670);
  nor GNAME9213(G9213,G21723,G8850);
  and GNAME9214(G9214,G9212,G9213);
  nor GNAME9215(G9215,G21699,G8848);
  and GNAME9216(G9216,G9212,G9215);
  nor GNAME9217(G9217,G8848,G8850);
  and GNAME9218(G9218,G9212,G9217);
  nor GNAME9219(G9219,G21670,G8846);
  nor GNAME9220(G9220,G21699,G21723);
  and GNAME9221(G9221,G9219,G9220);
  and GNAME9222(G9222,G9213,G9219);
  and GNAME9223(G9223,G9215,G9219);
  and GNAME9224(G9224,G9217,G9219);
  nor GNAME9225(G9225,G21631,G8844);
  and GNAME9226(G9226,G9220,G9225);
  and GNAME9227(G9227,G9213,G9225);
  and GNAME9228(G9228,G9215,G9225);
  and GNAME9229(G9229,G9217,G9225);
  nor GNAME9230(G9230,G8844,G8846);
  and GNAME9231(G9231,G9220,G9230);
  and GNAME9232(G9232,G9213,G9230);
  and GNAME9233(G9233,G9215,G9230);
  and GNAME9234(G9234,G9217,G9230);
  and GNAME9235(G9235,G9212,G9220);
  and GNAME9236(G9236,G21598,G8796,G8791);
  and GNAME9237(G9237,G8743,G8792);
  and GNAME9238(G9238,G59428,G8822);
  and GNAME9239(G9239,G13443,G8863);
  and GNAME9240(G9240,G13968,G13969,G13446,G8893);
  and GNAME9241(G9241,G13464,G8872);
  and GNAME9242(G9242,G8863,G13505);
  and GNAME9243(G9243,G9795,G9799);
  and GNAME9244(G9244,G59428,G10319);
  nand GNAME9245(G9245,G9108,G8782,G8746);
  nor GNAME9246(G9246,G9951,G9832,G9849);
  and GNAME9247(G9247,G13815,G9108);
  nor GNAME9248(G9248,G59425,G13802);
  nand GNAME9249(G9249,G13845,G13846);
  nand GNAME9250(G9250,G13871,G13872);
  nand GNAME9251(G9251,G13874,G13875);
  nand GNAME9252(G9252,G13877,G13878);
  nand GNAME9253(G9253,G13884,G13885);
  nand GNAME9254(G9254,G13896,G13897);
  nand GNAME9255(G9255,G13893,G13894);
  nand GNAME9256(G9256,G13927,G13928);
  nand GNAME9257(G9257,G13833,G13834);
  nand GNAME9258(G9258,G13835,G13836);
  nand GNAME9259(G9259,G13837,G13838);
  nand GNAME9260(G9260,G13841,G13842);
  nand GNAME9261(G9261,G13848,G13849);
  nand GNAME9262(G9262,G13880,G13881);
  nand GNAME9263(G9263,G13887,G13888);
  nand GNAME9264(G9264,G13890,G13891);
  nand GNAME9265(G9265,G13899,G13900);
  nand GNAME9266(G9266,G13903,G13904);
  nand GNAME9267(G9267,G13905,G13906);
  nand GNAME9268(G9268,G13911,G13912);
  nand GNAME9269(G9269,G13913,G13914);
  nand GNAME9270(G9270,G13919,G13920);
  nand GNAME9271(G9271,G13921,G13922);
  nand GNAME9272(G9272,G13923,G13924);
  nand GNAME9273(G9273,G13925,G13926);
  nand GNAME9274(G9274,G13932,G13933);
  nand GNAME9275(G9275,G13934,G13935);
  nand GNAME9276(G9276,G13936,G13937);
  nand GNAME9277(G9277,G13938,G13939);
  nand GNAME9278(G9278,G13940,G13941);
  nand GNAME9279(G9279,G13942,G13943);
  nand GNAME9280(G9280,G13944,G13945);
  nand GNAME9281(G9281,G13946,G13947);
  nand GNAME9282(G9282,G13948,G13949);
  nand GNAME9283(G9283,G13950,G13951);
  nand GNAME9284(G9284,G13952,G13953);
  nand GNAME9285(G9285,G13954,G13955);
  nand GNAME9286(G9286,G13956,G13957);
  nand GNAME9287(G9287,G13958,G13959);
  nand GNAME9288(G9288,G13960,G13961);
  nand GNAME9289(G9289,G13962,G13963);
  nand GNAME9290(G9290,G13964,G13965);
  and GNAME9291(G9291,G9850,G9851,G9852,G9853);
  and GNAME9292(G9292,G9854,G9855,G9856,G9857);
  and GNAME9293(G9293,G9858,G9859,G9860,G9861);
  and GNAME9294(G9294,G9862,G9863,G9864,G9865);
  and GNAME9295(G9295,G9918,G9919,G9920,G9921);
  and GNAME9296(G9296,G9922,G9923,G9924,G9925);
  and GNAME9297(G9297,G9926,G9927,G9928,G9929);
  and GNAME9298(G9298,G9930,G9931,G9932,G9933);
  and GNAME9299(G9299,G9935,G9936,G9937,G9938);
  and GNAME9300(G9300,G9939,G9940,G9941,G9942);
  and GNAME9301(G9301,G9943,G9944,G9945,G9946);
  and GNAME9302(G9302,G9947,G9948,G9949,G9950);
  and GNAME9303(G9303,G9901,G9902,G9903,G9904);
  and GNAME9304(G9304,G9905,G9906,G9907,G9908);
  and GNAME9305(G9305,G9909,G9910,G9911,G9912);
  and GNAME9306(G9306,G9913,G9914,G9915,G9916);
  and GNAME9307(G9307,G9884,G9885,G9886,G9887);
  and GNAME9308(G9308,G9888,G9889,G9890,G9891);
  and GNAME9309(G9309,G9892,G9893,G9894,G9895);
  and GNAME9310(G9310,G9896,G9897,G9898,G9899);
  and GNAME9311(G9311,G9833,G9834,G9835,G9836);
  and GNAME9312(G9312,G9837,G9838,G9839,G9840);
  and GNAME9313(G9313,G9841,G9842,G9843,G9844);
  and GNAME9314(G9314,G9845,G9846,G9847,G9848);
  and GNAME9315(G9315,G9816,G9817,G9818,G9819);
  and GNAME9316(G9316,G9820,G9821,G9822,G9823);
  and GNAME9317(G9317,G9824,G9825,G9826,G9827);
  and GNAME9318(G9318,G9828,G9829,G9830,G9831);
  and GNAME9319(G9319,G9867,G9868,G9869,G9870);
  and GNAME9320(G9320,G9871,G9872,G9873,G9874);
  and GNAME9321(G9321,G9875,G9876,G9877,G9878);
  and GNAME9322(G9322,G9879,G9880,G9881,G9882);
  or GNAME9323(G9323,G59398,G59397,G59396,G59395);
  nor GNAME9324(G9324,G9323,G59399,G59400,G59401,G59402);
  or GNAME9325(G9325,G59406,G59405,G59404,G59403);
  nor GNAME9326(G9326,G9325,G59407,G59408,G59409,G59410);
  or GNAME9327(G9327,G59414,G59413,G59412,G59411);
  nor GNAME9328(G9328,G9327,G59415,G59416,G59417,G59418);
  or GNAME9329(G9329,G59422,G59421,G59420,G59419);
  nor GNAME9330(G9330,G9329,G10005,G59423,G59424);
  and GNAME9331(G9331,G10028,G10026,G10025);
  and GNAME9332(G9332,G10034,G10032,G10031);
  and GNAME9333(G9333,G10040,G10038,G10037);
  and GNAME9334(G9334,G10046,G10044,G10043);
  and GNAME9335(G9335,G10052,G10050,G10049);
  and GNAME9336(G9336,G10058,G10056,G10055);
  and GNAME9337(G9337,G10064,G10062,G10061);
  and GNAME9338(G9338,G10070,G10068,G10067);
  and GNAME9339(G9339,G10076,G10074,G10073);
  and GNAME9340(G9340,G10082,G10080,G10079);
  and GNAME9341(G9341,G10088,G10086,G10085);
  and GNAME9342(G9342,G10094,G10092,G10091);
  and GNAME9343(G9343,G10101,G10099,G10095);
  and GNAME9344(G9344,G10107,G10105,G10095);
  and GNAME9345(G9345,G10113,G10111,G10095);
  and GNAME9346(G9346,G10119,G10117,G10095);
  and GNAME9347(G9347,G10125,G10123,G10095);
  and GNAME9348(G9348,G10131,G10129,G10095);
  and GNAME9349(G9349,G10137,G10135,G10095);
  and GNAME9350(G9350,G10143,G10141,G10095);
  and GNAME9351(G9351,G10149,G10147,G10095);
  and GNAME9352(G9352,G10155,G10153,G10095);
  and GNAME9353(G9353,G10161,G10095,G10158);
  and GNAME9354(G9354,G10167,G10095,G10166);
  and GNAME9355(G9355,G10173,G10095,G10172);
  and GNAME9356(G9356,G10179,G10095,G10178);
  and GNAME9357(G9357,G10095,G10184,G10189,G10186);
  and GNAME9358(G9358,G10095,G10190,G10195,G10192);
  and GNAME9359(G9359,G10199,G10200);
  and GNAME9360(G9360,G10205,G10206);
  and GNAME9361(G9361,G10210,G10208,G10213);
  and GNAME9362(G9362,G10216,G10214,G10219);
  and GNAME9363(G9363,G10812,G10809,G10810);
  and GNAME9364(G9364,G9832,G8781,G9951);
  and GNAME9365(G9365,G10838,G10836,G10837);
  and GNAME9366(G9366,G13854,G13855,G13856,G13857);
  and GNAME9367(G9367,G10847,G10845,G10846);
  and GNAME9368(G9368,G10853,G10851,G10852);
  and GNAME9369(G9369,G10859,G10857,G10858);
  and GNAME9370(G9370,G10865,G10863,G10864);
  and GNAME9371(G9371,G10871,G10869,G10870);
  and GNAME9372(G9372,G10877,G10875,G10876);
  and GNAME9373(G9373,G10883,G10881,G10882);
  and GNAME9374(G9374,G10889,G10887,G10888);
  and GNAME9375(G9375,G10895,G10893,G10894);
  and GNAME9376(G9376,G10901,G10899,G10900);
  and GNAME9377(G9377,G10907,G10905,G10906);
  and GNAME9378(G9378,G10913,G10911,G10912);
  and GNAME9379(G9379,G10919,G10917,G10918);
  and GNAME9380(G9380,G10925,G10923,G10924);
  and GNAME9381(G9381,G10931,G10929,G10930);
  and GNAME9382(G9382,G10937,G10935,G10936);
  and GNAME9383(G9383,G10943,G10941,G10942);
  and GNAME9384(G9384,G10949,G10947,G10948);
  and GNAME9385(G9385,G10955,G10953,G10954);
  and GNAME9386(G9386,G10961,G10959,G10960);
  and GNAME9387(G9387,G10967,G10965,G10966);
  and GNAME9388(G9388,G10973,G10971,G10972);
  and GNAME9389(G9389,G10979,G10977,G10978);
  and GNAME9390(G9390,G10985,G10983,G10984);
  and GNAME9391(G9391,G10991,G10989,G10990);
  and GNAME9392(G9392,G10997,G10995,G10996);
  and GNAME9393(G9393,G11003,G11001,G11002);
  and GNAME9394(G9394,G11009,G11007,G11008);
  and GNAME9395(G9395,G11015,G11013,G11018);
  and GNAME9396(G9396,G11021,G11019,G11024);
  and GNAME9397(G9397,G11027,G11025,G11030);
  and GNAME9398(G9398,G11033,G11031,G11036);
  and GNAME9399(G9399,G13869,G13870);
  and GNAME9400(G9400,G13882,G13883);
  and GNAME9401(G9401,G11129,G11127,G11124);
  and GNAME9402(G9402,G11150,G11146,G11149);
  and GNAME9403(G9403,G11178,G11174,G11177);
  and GNAME9404(G9404,G11204,G11202,G11203);
  and GNAME9405(G9405,G11213,G11211,G11212);
  and GNAME9406(G9406,G11222,G11220,G11221);
  and GNAME9407(G9407,G11231,G11229,G11230);
  and GNAME9408(G9408,G11240,G11238,G11239);
  and GNAME9409(G9409,G11249,G11247,G11248);
  and GNAME9410(G9410,G11258,G11256,G11257);
  and GNAME9411(G9411,G11267,G11265,G11266);
  and GNAME9412(G9412,G11286,G11284,G11285);
  and GNAME9413(G9413,G11292,G11290,G11291);
  and GNAME9414(G9414,G11298,G11296,G11297);
  and GNAME9415(G9415,G11304,G11302,G11303);
  and GNAME9416(G9416,G11310,G11308,G11309);
  and GNAME9417(G9417,G11316,G11314,G11315);
  and GNAME9418(G9418,G11322,G11320,G11321);
  and GNAME9419(G9419,G11328,G11326,G11327);
  and GNAME9420(G9420,G11347,G11345,G11346);
  and GNAME9421(G9421,G11353,G11351,G11352);
  and GNAME9422(G9422,G11359,G11357,G11358);
  and GNAME9423(G9423,G11365,G11363,G11364);
  and GNAME9424(G9424,G11371,G11369,G11370);
  and GNAME9425(G9425,G11377,G11375,G11376);
  and GNAME9426(G9426,G11383,G11381,G11382);
  and GNAME9427(G9427,G11389,G11387,G11388);
  and GNAME9428(G9428,G11408,G11406,G11407);
  and GNAME9429(G9429,G11414,G11412,G11413);
  and GNAME9430(G9430,G11420,G11418,G11419);
  and GNAME9431(G9431,G11426,G11424,G11425);
  and GNAME9432(G9432,G11432,G11430,G11431);
  and GNAME9433(G9433,G11438,G11436,G11437);
  and GNAME9434(G9434,G11444,G11442,G11443);
  and GNAME9435(G9435,G11450,G11448,G11449);
  and GNAME9436(G9436,G11469,G11467,G11468);
  and GNAME9437(G9437,G11475,G11473,G11474);
  and GNAME9438(G9438,G11481,G11479,G11480);
  and GNAME9439(G9439,G11487,G11485,G11486);
  and GNAME9440(G9440,G11493,G11491,G11492);
  and GNAME9441(G9441,G11499,G11497,G11498);
  and GNAME9442(G9442,G11505,G11503,G11504);
  and GNAME9443(G9443,G11511,G11509,G11510);
  and GNAME9444(G9444,G11530,G11528,G11529);
  and GNAME9445(G9445,G11536,G11534,G11535);
  and GNAME9446(G9446,G11542,G11540,G11541);
  and GNAME9447(G9447,G11548,G11546,G11547);
  and GNAME9448(G9448,G11554,G11552,G11553);
  and GNAME9449(G9449,G11560,G11558,G11559);
  and GNAME9450(G9450,G11566,G11564,G11565);
  and GNAME9451(G9451,G11572,G11570,G11571);
  and GNAME9452(G9452,G11591,G11589,G11590);
  and GNAME9453(G9453,G11597,G11595,G11596);
  and GNAME9454(G9454,G11603,G11601,G11602);
  and GNAME9455(G9455,G11609,G11607,G11608);
  and GNAME9456(G9456,G11615,G11613,G11614);
  and GNAME9457(G9457,G11621,G11619,G11620);
  and GNAME9458(G9458,G11627,G11625,G11626);
  and GNAME9459(G9459,G11633,G11631,G11632);
  and GNAME9460(G9460,G11652,G11650,G11651);
  and GNAME9461(G9461,G11658,G11656,G11657);
  and GNAME9462(G9462,G11664,G11662,G11663);
  and GNAME9463(G9463,G11670,G11668,G11669);
  and GNAME9464(G9464,G11676,G11674,G11675);
  and GNAME9465(G9465,G11682,G11680,G11681);
  and GNAME9466(G9466,G11688,G11686,G11687);
  and GNAME9467(G9467,G11694,G11692,G11693);
  and GNAME9468(G9468,G11713,G11711,G11712);
  and GNAME9469(G9469,G11719,G11717,G11718);
  and GNAME9470(G9470,G11725,G11723,G11724);
  and GNAME9471(G9471,G11731,G11729,G11730);
  and GNAME9472(G9472,G11737,G11735,G11736);
  and GNAME9473(G9473,G11743,G11741,G11742);
  and GNAME9474(G9474,G11749,G11747,G11748);
  and GNAME9475(G9475,G11755,G11753,G11754);
  and GNAME9476(G9476,G11774,G11772,G11773);
  and GNAME9477(G9477,G11780,G11778,G11779);
  and GNAME9478(G9478,G11786,G11784,G11785);
  and GNAME9479(G9479,G11792,G11790,G11791);
  and GNAME9480(G9480,G11798,G11796,G11797);
  and GNAME9481(G9481,G11804,G11802,G11803);
  and GNAME9482(G9482,G11810,G11808,G11809);
  and GNAME9483(G9483,G11816,G11814,G11815);
  and GNAME9484(G9484,G11835,G11833,G11834);
  and GNAME9485(G9485,G11841,G11839,G11840);
  and GNAME9486(G9486,G11847,G11845,G11846);
  and GNAME9487(G9487,G11853,G11851,G11852);
  and GNAME9488(G9488,G11859,G11857,G11858);
  and GNAME9489(G9489,G11865,G11863,G11864);
  and GNAME9490(G9490,G11871,G11869,G11870);
  and GNAME9491(G9491,G11877,G11875,G11876);
  and GNAME9492(G9492,G11896,G11894,G11895);
  and GNAME9493(G9493,G11902,G11900,G11901);
  and GNAME9494(G9494,G11908,G11906,G11907);
  and GNAME9495(G9495,G11914,G11912,G11913);
  and GNAME9496(G9496,G11920,G11918,G11919);
  and GNAME9497(G9497,G11926,G11924,G11925);
  and GNAME9498(G9498,G11932,G11930,G11931);
  and GNAME9499(G9499,G11938,G11936,G11937);
  and GNAME9500(G9500,G11957,G11955,G11956);
  and GNAME9501(G9501,G11963,G11961,G11962);
  and GNAME9502(G9502,G11969,G11967,G11968);
  and GNAME9503(G9503,G11975,G11973,G11974);
  and GNAME9504(G9504,G11981,G11979,G11980);
  and GNAME9505(G9505,G11987,G11985,G11986);
  and GNAME9506(G9506,G11993,G11991,G11992);
  and GNAME9507(G9507,G11999,G11997,G11998);
  and GNAME9508(G9508,G12018,G12016,G12017);
  and GNAME9509(G9509,G12024,G12022,G12023);
  and GNAME9510(G9510,G12030,G12028,G12029);
  and GNAME9511(G9511,G12036,G12034,G12035);
  and GNAME9512(G9512,G12042,G12040,G12041);
  and GNAME9513(G9513,G12048,G12046,G12047);
  and GNAME9514(G9514,G12054,G12052,G12053);
  and GNAME9515(G9515,G12060,G12058,G12059);
  and GNAME9516(G9516,G12079,G12077,G12078);
  and GNAME9517(G9517,G12085,G12083,G12084);
  and GNAME9518(G9518,G12091,G12089,G12090);
  and GNAME9519(G9519,G12097,G12095,G12096);
  and GNAME9520(G9520,G12103,G12101,G12102);
  and GNAME9521(G9521,G12109,G12107,G12108);
  and GNAME9522(G9522,G12115,G12113,G12114);
  and GNAME9523(G9523,G12121,G12119,G12120);
  and GNAME9524(G9524,G12140,G12138,G12139);
  and GNAME9525(G9525,G12146,G12144,G12145);
  and GNAME9526(G9526,G12152,G12150,G12151);
  and GNAME9527(G9527,G12158,G12156,G12157);
  and GNAME9528(G9528,G12164,G12162,G12163);
  and GNAME9529(G9529,G12170,G12168,G12169);
  and GNAME9530(G9530,G12176,G12174,G12175);
  and GNAME9531(G9531,G12182,G12180,G12181);
  nand GNAME9532(G9532,G22276,G12185,G12186);
  and GNAME9533(G9533,G12306,G12307,G12308,G12309);
  and GNAME9534(G9534,G12310,G12311,G12312,G12313);
  and GNAME9535(G9535,G12314,G12315,G12316,G12317);
  and GNAME9536(G9536,G12318,G12319,G12320,G12321);
  and GNAME9537(G9537,G12322,G12323,G12324,G12325);
  and GNAME9538(G9538,G12326,G12327,G12328,G12329);
  and GNAME9539(G9539,G12330,G12331,G12332,G12333);
  and GNAME9540(G9540,G12334,G12335,G12336,G12337);
  and GNAME9541(G9541,G12338,G12339,G12340,G12341);
  and GNAME9542(G9542,G12342,G12343,G12344,G12345);
  and GNAME9543(G9543,G12346,G12347,G12348,G12349);
  and GNAME9544(G9544,G12350,G12351,G12352,G12353);
  and GNAME9545(G9545,G12354,G12355,G12356,G12357);
  and GNAME9546(G9546,G12358,G12359,G12360,G12361);
  and GNAME9547(G9547,G12362,G12363,G12364,G12365);
  and GNAME9548(G9548,G12366,G12367,G12368,G12369);
  and GNAME9549(G9549,G12370,G12371,G12372,G12373);
  and GNAME9550(G9550,G12374,G12375,G12376,G12377);
  and GNAME9551(G9551,G12378,G12379,G12380,G12381);
  and GNAME9552(G9552,G12382,G12383,G12384,G12385);
  and GNAME9553(G9553,G12386,G12387,G12388,G12389);
  and GNAME9554(G9554,G12390,G12391,G12392,G12393);
  and GNAME9555(G9555,G12394,G12395,G12396,G12397);
  and GNAME9556(G9556,G12398,G12399,G12400,G12401);
  and GNAME9557(G9557,G12402,G12403,G12404,G12405);
  and GNAME9558(G9558,G12406,G12407,G12408,G12409);
  and GNAME9559(G9559,G12410,G12411,G12412,G12413);
  and GNAME9560(G9560,G12414,G12415,G12416,G12417);
  and GNAME9561(G9561,G12418,G12419,G12420,G12421);
  and GNAME9562(G9562,G12422,G12423,G12424,G12425);
  and GNAME9563(G9563,G12426,G12427,G12428,G12429);
  and GNAME9564(G9564,G12430,G12431,G12432,G12433);
  and GNAME9565(G9565,G12435,G12436,G12437,G12438);
  and GNAME9566(G9566,G12439,G12440,G12441,G12442);
  and GNAME9567(G9567,G12443,G12444,G12445,G12446);
  and GNAME9568(G9568,G12447,G12448,G12449,G12450);
  and GNAME9569(G9569,G12451,G12452,G12453,G12454);
  and GNAME9570(G9570,G12455,G12456,G12457,G12458);
  and GNAME9571(G9571,G12459,G12460,G12461,G12462);
  and GNAME9572(G9572,G12463,G12464,G12465,G12466);
  and GNAME9573(G9573,G12467,G12468,G12469,G12470);
  and GNAME9574(G9574,G12471,G12472,G12473,G12474);
  and GNAME9575(G9575,G12475,G12476,G12477,G12478);
  and GNAME9576(G9576,G12479,G12480,G12481,G12482);
  and GNAME9577(G9577,G12483,G12484,G12485,G12486);
  and GNAME9578(G9578,G12487,G12488,G12489,G12490);
  and GNAME9579(G9579,G12491,G12492,G12493,G12494);
  and GNAME9580(G9580,G12495,G12496,G12497,G12498);
  and GNAME9581(G9581,G12499,G12500,G12501,G12502);
  and GNAME9582(G9582,G12503,G12504,G12505,G12506);
  and GNAME9583(G9583,G12507,G12508,G12509,G12510);
  and GNAME9584(G9584,G12511,G12512,G12513,G12514);
  and GNAME9585(G9585,G12515,G12516,G12517,G12518);
  and GNAME9586(G9586,G12519,G12520,G12521,G12522);
  and GNAME9587(G9587,G12523,G12524,G12525,G12526);
  and GNAME9588(G9588,G12527,G12528,G12529,G12530);
  and GNAME9589(G9589,G12531,G12532,G12533,G12534);
  and GNAME9590(G9590,G12535,G12536,G12537,G12538);
  and GNAME9591(G9591,G12539,G12540,G12541,G12542);
  and GNAME9592(G9592,G12543,G12544,G12545,G12546);
  and GNAME9593(G9593,G12547,G12548,G12549,G12550);
  and GNAME9594(G9594,G12551,G12552,G12553,G12554);
  and GNAME9595(G9595,G12555,G12556,G12557,G12558);
  and GNAME9596(G9596,G12559,G12560,G12561,G12562);
  and GNAME9597(G9597,G12563,G12564,G12565,G12566);
  and GNAME9598(G9598,G12567,G12568,G12569,G12570);
  and GNAME9599(G9599,G12571,G12572,G12573,G12574);
  and GNAME9600(G9600,G12575,G12576,G12577,G12578);
  and GNAME9601(G9601,G12580,G12581,G12582,G12583);
  and GNAME9602(G9602,G12584,G12585,G12586,G12587);
  and GNAME9603(G9603,G12588,G12589,G12590,G12591);
  and GNAME9604(G9604,G12592,G12593,G12594,G12595);
  and GNAME9605(G9605,G12597,G12598,G12599,G12600);
  and GNAME9606(G9606,G12601,G12602,G12603,G12604);
  and GNAME9607(G9607,G12605,G12606,G12607,G12608);
  and GNAME9608(G9608,G12609,G12610,G12611,G12612);
  and GNAME9609(G9609,G12614,G12615,G12616,G12617);
  and GNAME9610(G9610,G12618,G12619,G12620,G12621);
  and GNAME9611(G9611,G12622,G12623,G12624,G12625);
  and GNAME9612(G9612,G12626,G12627,G12628,G12629);
  and GNAME9613(G9613,G12631,G12632,G12633,G12634);
  and GNAME9614(G9614,G12635,G12636,G12637,G12638);
  and GNAME9615(G9615,G12639,G12640,G12641,G12642);
  and GNAME9616(G9616,G12643,G12644,G12645,G12646);
  and GNAME9617(G9617,G12648,G12649,G12650,G12651);
  and GNAME9618(G9618,G12652,G12653,G12654,G12655);
  and GNAME9619(G9619,G12656,G12657,G12658,G12659);
  and GNAME9620(G9620,G12660,G12661,G12662,G12663);
  and GNAME9621(G9621,G12665,G12666,G12667,G12668);
  and GNAME9622(G9622,G12669,G12670,G12671,G12672);
  and GNAME9623(G9623,G12673,G12674,G12675,G12676);
  and GNAME9624(G9624,G12677,G12678,G12679,G12680);
  and GNAME9625(G9625,G12682,G12683,G12684,G12685);
  and GNAME9626(G9626,G12686,G12687,G12688,G12689);
  and GNAME9627(G9627,G12690,G12691,G12692,G12693);
  and GNAME9628(G9628,G12694,G12695,G12696,G12697);
  and GNAME9629(G9629,G12699,G12700,G12701,G12702);
  and GNAME9630(G9630,G12703,G12704,G12705,G12706);
  and GNAME9631(G9631,G12707,G12708,G12709,G12710);
  and GNAME9632(G9632,G12711,G12712,G12713,G12714);
  and GNAME9633(G9633,G12716,G12717,G12718,G12719);
  and GNAME9634(G9634,G12720,G12721,G12722,G12723);
  and GNAME9635(G9635,G12724,G12725,G12726,G12727);
  and GNAME9636(G9636,G12728,G12729,G12730,G12731);
  and GNAME9637(G9637,G12733,G12734,G12735,G12736);
  and GNAME9638(G9638,G12737,G12738,G12739,G12740);
  and GNAME9639(G9639,G12741,G12742,G12743,G12744);
  and GNAME9640(G9640,G12745,G12746,G12747,G12748);
  and GNAME9641(G9641,G12750,G12751,G12752,G12753);
  and GNAME9642(G9642,G12754,G12755,G12756,G12757);
  and GNAME9643(G9643,G12758,G12759,G12760,G12761);
  and GNAME9644(G9644,G12762,G12763,G12764,G12765);
  and GNAME9645(G9645,G12767,G12768,G12769,G12770);
  and GNAME9646(G9646,G12771,G12772,G12773,G12774);
  and GNAME9647(G9647,G12775,G12776,G12777,G12778);
  and GNAME9648(G9648,G12779,G12780,G12781,G12782);
  and GNAME9649(G9649,G12784,G12785,G12786,G12787);
  and GNAME9650(G9650,G12788,G12789,G12790,G12791);
  and GNAME9651(G9651,G12792,G12793,G12794,G12795);
  and GNAME9652(G9652,G12796,G12797,G12798,G12799);
  and GNAME9653(G9653,G12801,G12802,G12803,G12804);
  and GNAME9654(G9654,G12805,G12806,G12807,G12808);
  and GNAME9655(G9655,G12809,G12810,G12811,G12812);
  and GNAME9656(G9656,G12813,G12814,G12815,G12816);
  and GNAME9657(G9657,G12818,G12819,G12820,G12821);
  and GNAME9658(G9658,G12822,G12823,G12824,G12825);
  and GNAME9659(G9659,G12826,G12827,G12828,G12829);
  and GNAME9660(G9660,G12830,G12831,G12832,G12833);
  and GNAME9661(G9661,G9883,G12994,G12995);
  and GNAME9662(G9662,G13030,G13031,G13032,G13033);
  and GNAME9663(G9663,G13034,G13035,G13036,G13037);
  and GNAME9664(G9664,G13038,G13039,G13040,G13041);
  and GNAME9665(G9665,G13042,G13043,G13044,G13045);
  and GNAME9666(G9666,G13013,G13014,G13015,G13016);
  and GNAME9667(G9667,G13017,G13018,G13019,G13020);
  and GNAME9668(G9668,G13021,G13022,G13023,G13024);
  and GNAME9669(G9669,G13025,G13026,G13027,G13028);
  and GNAME9670(G9670,G12996,G12997,G12998,G12999);
  and GNAME9671(G9671,G13000,G13001,G13002,G13003);
  and GNAME9672(G9672,G13004,G13005,G13006,G13007);
  and GNAME9673(G9673,G13008,G13009,G13010,G13011);
  and GNAME9674(G9674,G13085,G13086,G13087,G13088);
  and GNAME9675(G9675,G13089,G13090,G13091,G13092);
  and GNAME9676(G9676,G13093,G13094,G13095,G13096);
  and GNAME9677(G9677,G13097,G13098,G13099,G13100);
  and GNAME9678(G9678,G13068,G13069,G13070,G13071);
  and GNAME9679(G9679,G13072,G13073,G13074,G13075);
  and GNAME9680(G9680,G13076,G13077,G13078,G13079);
  and GNAME9681(G9681,G13080,G13081,G13082,G13083);
  and GNAME9682(G9682,G13051,G13052,G13053,G13054);
  and GNAME9683(G9683,G13055,G13056,G13057,G13058);
  and GNAME9684(G9684,G13059,G13060,G13061,G13062);
  and GNAME9685(G9685,G13063,G13064,G13065,G13066);
  and GNAME9686(G9686,G13140,G13141,G13142,G13143);
  and GNAME9687(G9687,G13144,G13145,G13146,G13147);
  and GNAME9688(G9688,G13148,G13149,G13150,G13151);
  and GNAME9689(G9689,G13152,G13153,G13154,G13155);
  and GNAME9690(G9690,G13123,G13124,G13125,G13126);
  and GNAME9691(G9691,G13127,G13128,G13129,G13130);
  and GNAME9692(G9692,G13131,G13132,G13133,G13134);
  and GNAME9693(G9693,G13135,G13136,G13137,G13138);
  and GNAME9694(G9694,G13106,G13107,G13108,G13109);
  and GNAME9695(G9695,G13110,G13111,G13112,G13113);
  and GNAME9696(G9696,G13114,G13115,G13116,G13117);
  and GNAME9697(G9697,G13118,G13119,G13120,G13121);
  and GNAME9698(G9698,G13195,G13196,G13197,G13198);
  and GNAME9699(G9699,G13199,G13200,G13201,G13202);
  and GNAME9700(G9700,G13203,G13204,G13205,G13206);
  and GNAME9701(G9701,G13207,G13208,G13209,G13210);
  and GNAME9702(G9702,G13178,G13179,G13180,G13181);
  and GNAME9703(G9703,G13182,G13183,G13184,G13185);
  and GNAME9704(G9704,G13186,G13187,G13188,G13189);
  and GNAME9705(G9705,G13190,G13191,G13192,G13193);
  and GNAME9706(G9706,G13161,G13162,G13163,G13164);
  and GNAME9707(G9707,G13165,G13166,G13167,G13168);
  and GNAME9708(G9708,G13169,G13170,G13171,G13172);
  and GNAME9709(G9709,G13173,G13174,G13175,G13176);
  and GNAME9710(G9710,G13251,G13252,G13253,G13254);
  and GNAME9711(G9711,G13255,G13256,G13257,G13258);
  and GNAME9712(G9712,G13259,G13260,G13261,G13262);
  and GNAME9713(G9713,G13263,G13264,G13265,G13266);
  and GNAME9714(G9714,G13234,G13235,G13236,G13237);
  and GNAME9715(G9715,G13238,G13239,G13240,G13241);
  and GNAME9716(G9716,G13242,G13243,G13244,G13245);
  and GNAME9717(G9717,G13246,G13247,G13248,G13249);
  and GNAME9718(G9718,G13217,G13218,G13219,G13220);
  and GNAME9719(G9719,G13221,G13222,G13223,G13224);
  and GNAME9720(G9720,G13225,G13226,G13227,G13228);
  and GNAME9721(G9721,G13229,G13230,G13231,G13232);
  and GNAME9722(G9722,G13307,G13308,G13309,G13310);
  and GNAME9723(G9723,G13311,G13312,G13313,G13314);
  and GNAME9724(G9724,G13315,G13316,G13317,G13318);
  and GNAME9725(G9725,G13319,G13320,G13321,G13322);
  and GNAME9726(G9726,G13290,G13291,G13292,G13293);
  and GNAME9727(G9727,G13294,G13295,G13296,G13297);
  and GNAME9728(G9728,G13298,G13299,G13300,G13301);
  and GNAME9729(G9729,G13302,G13303,G13304,G13305);
  and GNAME9730(G9730,G13273,G13274,G13275,G13276);
  and GNAME9731(G9731,G13277,G13278,G13279,G13280);
  and GNAME9732(G9732,G13281,G13282,G13283,G13284);
  and GNAME9733(G9733,G13285,G13286,G13287,G13288);
  and GNAME9734(G9734,G13328,G13326,G13327);
  and GNAME9735(G9735,G13363,G13364,G13365,G13366);
  and GNAME9736(G9736,G13367,G13368,G13369,G13370);
  and GNAME9737(G9737,G13371,G13372,G13373,G13374);
  and GNAME9738(G9738,G13375,G13376,G13377,G13378);
  and GNAME9739(G9739,G13346,G13347,G13348,G13349);
  and GNAME9740(G9740,G13350,G13351,G13352,G13353);
  and GNAME9741(G9741,G13354,G13355,G13356,G13357);
  and GNAME9742(G9742,G13358,G13359,G13360,G13361);
  and GNAME9743(G9743,G13329,G13330,G13331,G13332);
  and GNAME9744(G9744,G13333,G13334,G13335,G13336);
  and GNAME9745(G9745,G13337,G13338,G13339,G13340);
  and GNAME9746(G9746,G13341,G13342,G13343,G13344);
  and GNAME9747(G9747,G13384,G13382,G13383);
  and GNAME9748(G9748,G13419,G13420,G13421,G13422);
  and GNAME9749(G9749,G13423,G13424,G13425,G13426);
  and GNAME9750(G9750,G13427,G13428,G13429,G13430);
  and GNAME9751(G9751,G13431,G13432,G13433,G13434);
  and GNAME9752(G9752,G13402,G13403,G13404,G13405);
  and GNAME9753(G9753,G13406,G13407,G13408,G13409);
  and GNAME9754(G9754,G13410,G13411,G13412,G13413);
  and GNAME9755(G9755,G13414,G13415,G13416,G13417);
  and GNAME9756(G9756,G13385,G13386,G13387,G13388);
  and GNAME9757(G9757,G13389,G13390,G13391,G13392);
  and GNAME9758(G9758,G13393,G13394,G13395,G13396);
  and GNAME9759(G9759,G13397,G13398,G13399,G13400);
  and GNAME9760(G9760,G13440,G13438,G13439);
  and GNAME9761(G9761,G13444,G13445);
  and GNAME9762(G9762,G9815,G8852,G13447,G13966);
  and GNAME9763(G9763,G13460,G13458,G13459);
  and GNAME9764(G9764,G13618,G13616,G13617);
  and GNAME9765(G9765,G13669,G13670,G13674,G13671,G13667);
  and GNAME9766(G9766,G13728,G13729,G13733,G13730,G13726);
  and GNAME9767(G9767,G13787,G13788,G13792,G13789,G13785);
  and GNAME9768(G9768,G13796,G13797,G13801,G13798,G13794);
  or GNAME9769(G9769,G8810,G8803);
  and GNAME9770(G9770,G13980,G9972,G9974);
  not GNAME9771(G9771,G35);
  or GNAME9772(G9772,G8924,G8925);
  and GNAME9773(G9773,G11073,G11071,G11072);
  nand GNAME9774(G9774,G11085,G9813,G8909);
  nand GNAME9775(G9775,G11087,G59426);
  and GNAME9776(G9776,G8759,G9866);
  nand GNAME9777(G9777,G8759,G13895);
  nand GNAME9778(G9778,G8888,G11083,G11084);
  not GNAME9779(G9779,G8856);
  not GNAME9780(G9780,G9243);
  not GNAME9781(G9781,G8743);
  not GNAME9782(G9782,G8745);
  not GNAME9783(G9783,G8784);
  not GNAME9784(G9784,G8811);
  not GNAME9785(G9785,G9111);
  not GNAME9786(G9786,G9112);
  not GNAME9787(G9787,G8759);
  not GNAME9788(G9788,G8769);
  not GNAME9789(G9789,G8824);
  not GNAME9790(G9790,G8827);
  not GNAME9791(G9791,G8826);
  not GNAME9792(G9792,G8828);
  not GNAME9793(G9793,G8825);
  not GNAME9794(G9794,G8907);
  not GNAME9795(G9795,G8940);
  not GNAME9796(G9796,G8833);
  not GNAME9797(G9797,G8802);
  not GNAME9798(G9798,G8790);
  not GNAME9799(G9799,G8813);
  nand GNAME9800(G9800,G8910,G8833);
  not GNAME9801(G9801,G8919);
  not GNAME9802(G9802,G8820);
  not GNAME9803(G9803,G8887);
  not GNAME9804(G9804,G8800);
  not GNAME9805(G9805,G8853);
  not GNAME9806(G9806,G8939);
  nand GNAME9807(G9807,G9238,G8796,G21598);
  or GNAME9808(G9808,G59393,G59394,G59758,G13985);
  nand GNAME9809(G9809,G8897,G9976,G59428);
  nand GNAME9810(G9810,G1588,G8839);
  nand GNAME9811(G9811,G8833,G8751,G8787);
  nand GNAME9812(G9812,G59425,G59428,G8802);
  nand GNAME9813(G9813,G59795,G8908);
  nand GNAME9814(G9814,G8817,G8812);
  not GNAME9815(G9815,G8894);
  nand GNAME9816(G9816,G59543,G8755);
  nand GNAME9817(G9817,G59535,G8758);
  nand GNAME9818(G9818,G59527,G8760);
  nand GNAME9819(G9819,G59519,G8764);
  nand GNAME9820(G9820,G59511,G8765);
  nand GNAME9821(G9821,G59503,G8766);
  nand GNAME9822(G9822,G59495,G8767);
  nand GNAME9823(G9823,G59487,G8770);
  nand GNAME9824(G9824,G59479,G8771);
  nand GNAME9825(G9825,G59471,G8772);
  nand GNAME9826(G9826,G59463,G8773);
  nand GNAME9827(G9827,G59455,G8775);
  nand GNAME9828(G9828,G59447,G8776);
  nand GNAME9829(G9829,G59439,G8777);
  nand GNAME9830(G9830,G59431,G8778);
  nand GNAME9831(G9831,G8779,G59551);
  not GNAME9832(G9832,G8780);
  nand GNAME9833(G9833,G8779,G59555);
  nand GNAME9834(G9834,G8755,G59547);
  nand GNAME9835(G9835,G8758,G59539);
  nand GNAME9836(G9836,G8760,G59531);
  nand GNAME9837(G9837,G8764,G59523);
  nand GNAME9838(G9838,G8765,G59515);
  nand GNAME9839(G9839,G8766,G59507);
  nand GNAME9840(G9840,G8767,G59499);
  nand GNAME9841(G9841,G8770,G59491);
  nand GNAME9842(G9842,G8771,G59483);
  nand GNAME9843(G9843,G8772,G59475);
  nand GNAME9844(G9844,G8773,G59467);
  nand GNAME9845(G9845,G8775,G59459);
  nand GNAME9846(G9846,G8776,G59451);
  nand GNAME9847(G9847,G8777,G59443);
  nand GNAME9848(G9848,G8778,G59435);
  not GNAME9849(G9849,G8796);
  nand GNAME9850(G9850,G8779,G59556);
  nand GNAME9851(G9851,G8755,G59548);
  nand GNAME9852(G9852,G8758,G59540);
  nand GNAME9853(G9853,G8760,G59532);
  nand GNAME9854(G9854,G8764,G59524);
  nand GNAME9855(G9855,G8765,G59516);
  nand GNAME9856(G9856,G8766,G59508);
  nand GNAME9857(G9857,G8767,G59500);
  nand GNAME9858(G9858,G8770,G59492);
  nand GNAME9859(G9859,G8771,G59484);
  nand GNAME9860(G9860,G8772,G59476);
  nand GNAME9861(G9861,G8773,G59468);
  nand GNAME9862(G9862,G8775,G59460);
  nand GNAME9863(G9863,G8776,G59452);
  nand GNAME9864(G9864,G8777,G59444);
  nand GNAME9865(G9865,G8778,G59436);
  not GNAME9866(G9866,G8792);
  nand GNAME9867(G9867,G8779,G59554);
  nand GNAME9868(G9868,G8755,G59546);
  nand GNAME9869(G9869,G8758,G59538);
  nand GNAME9870(G9870,G8760,G59530);
  nand GNAME9871(G9871,G8764,G59522);
  nand GNAME9872(G9872,G8765,G59514);
  nand GNAME9873(G9873,G8766,G59506);
  nand GNAME9874(G9874,G8767,G59498);
  nand GNAME9875(G9875,G8770,G59490);
  nand GNAME9876(G9876,G8771,G59482);
  nand GNAME9877(G9877,G8772,G59474);
  nand GNAME9878(G9878,G8773,G59466);
  nand GNAME9879(G9879,G8775,G59458);
  nand GNAME9880(G9880,G8776,G59450);
  nand GNAME9881(G9881,G8777,G59442);
  nand GNAME9882(G9882,G8778,G59434);
  not GNAME9883(G9883,G8781);
  nand GNAME9884(G9884,G8755,G59544);
  nand GNAME9885(G9885,G8758,G59536);
  nand GNAME9886(G9886,G8760,G59528);
  nand GNAME9887(G9887,G8764,G59520);
  nand GNAME9888(G9888,G8765,G59512);
  nand GNAME9889(G9889,G8766,G59504);
  nand GNAME9890(G9890,G8767,G59496);
  nand GNAME9891(G9891,G8770,G59488);
  nand GNAME9892(G9892,G8771,G59480);
  nand GNAME9893(G9893,G8772,G59472);
  nand GNAME9894(G9894,G8773,G59464);
  nand GNAME9895(G9895,G8775,G59456);
  nand GNAME9896(G9896,G8776,G59448);
  nand GNAME9897(G9897,G8777,G59440);
  nand GNAME9898(G9898,G8778,G59432);
  nand GNAME9899(G9899,G8779,G59552);
  not GNAME9900(G9900,G8783);
  nand GNAME9901(G9901,G8755,G59542);
  nand GNAME9902(G9902,G8758,G59534);
  nand GNAME9903(G9903,G8760,G59526);
  nand GNAME9904(G9904,G8764,G59518);
  nand GNAME9905(G9905,G8765,G59510);
  nand GNAME9906(G9906,G8766,G59502);
  nand GNAME9907(G9907,G8767,G59494);
  nand GNAME9908(G9908,G8770,G59486);
  nand GNAME9909(G9909,G8771,G59478);
  nand GNAME9910(G9910,G8772,G59470);
  nand GNAME9911(G9911,G8773,G59462);
  nand GNAME9912(G9912,G8775,G59454);
  nand GNAME9913(G9913,G8776,G59446);
  nand GNAME9914(G9914,G8777,G59438);
  nand GNAME9915(G9915,G8778,G59430);
  nand GNAME9916(G9916,G8779,G59550);
  not GNAME9917(G9917,G8782);
  nand GNAME9918(G9918,G8755,G59541);
  nand GNAME9919(G9919,G8758,G59533);
  nand GNAME9920(G9920,G8760,G59525);
  nand GNAME9921(G9921,G8764,G59517);
  nand GNAME9922(G9922,G8765,G59509);
  nand GNAME9923(G9923,G8766,G59501);
  nand GNAME9924(G9924,G8767,G59493);
  nand GNAME9925(G9925,G8770,G59485);
  nand GNAME9926(G9926,G8771,G59477);
  nand GNAME9927(G9927,G8772,G59469);
  nand GNAME9928(G9928,G8773,G59461);
  nand GNAME9929(G9929,G8775,G59453);
  nand GNAME9930(G9930,G8776,G59445);
  nand GNAME9931(G9931,G8777,G59437);
  nand GNAME9932(G9932,G8778,G59429);
  nand GNAME9933(G9933,G8779,G59549);
  not GNAME9934(G9934,G8852);
  nand GNAME9935(G9935,G8755,G59545);
  nand GNAME9936(G9936,G8758,G59537);
  nand GNAME9937(G9937,G8760,G59529);
  nand GNAME9938(G9938,G8764,G59521);
  nand GNAME9939(G9939,G8765,G59513);
  nand GNAME9940(G9940,G8766,G59505);
  nand GNAME9941(G9941,G8767,G59497);
  nand GNAME9942(G9942,G8770,G59489);
  nand GNAME9943(G9943,G8771,G59481);
  nand GNAME9944(G9944,G8772,G59473);
  nand GNAME9945(G9945,G8773,G59465);
  nand GNAME9946(G9946,G8775,G59457);
  nand GNAME9947(G9947,G8776,G59449);
  nand GNAME9948(G9948,G8777,G59441);
  nand GNAME9949(G9949,G8778,G59433);
  nand GNAME9950(G9950,G8779,G59553);
  not GNAME9951(G9951,G8746);
  not GNAME9952(G9952,G8786);
  not GNAME9953(G9953,G8788);
  nand GNAME9954(G9954,G8795,G59426,G13986);
  not GNAME9955(G9955,G8799);
  nand GNAME9956(G9956,G9954,G8877);
  nand GNAME9957(G9957,G9956,G21598);
  nand GNAME9958(G9958,G59426,G9866);
  or GNAME9959(G9959,G8751,G8743,G8785);
  nor GNAME9960(G9960,G8805,G8806);
  not GNAME9961(G9961,G8807);
  nand GNAME9962(G9962,G59392,G59802);
  nand GNAME9963(G9963,G8793,G9951,G9866);
  nand GNAME9964(G9964,G9963,G8781);
  nand GNAME9965(G9965,G8789,G8796);
  nand GNAME9966(G9966,G8784,G9965,G9832);
  nand GNAME9967(G9967,G8801,G13846);
  nand GNAME9968(G9968,G9966,G9883);
  nand GNAME9969(G9969,G8800,G8809);
  nand GNAME9970(G9970,G9969,G59801);
  nand GNAME9971(G9971,G59428,G8810);
  or GNAME9972(G9972,G1588,G8815);
  nand GNAME9973(G9973,G59426,G59428);
  nand GNAME9974(G9974,G9973,G8816);
  nand GNAME9975(G9975,G8804,G59390);
  nand GNAME9976(G9976,G9975,G8805);
  not GNAME9977(G9977,G8818);
  nand GNAME9978(G9978,G8818,G9866);
  nand GNAME9979(G9979,G8796,G9978);
  nand GNAME9980(G9980,G9977,G59797);
  nand GNAME9981(G9981,G9979,G9980);
  nand GNAME9982(G9982,G9981,G59426);
  nand GNAME9983(G9983,G9866,G8820);
  nand GNAME9984(G9984,G9982,G9983);
  nand GNAME9985(G9985,G8749,G9984);
  nand GNAME9986(G9986,G9985,G59428);
  and GNAME9987(G9987,G9797,G9986);
  nand GNAME9988(G9988,G8818,G13847);
  nand GNAME9989(G9989,G8749,G9988);
  or GNAME9990(G9990,G9104,G9804);
  not GNAME9991(G9991,G8864);
  nand GNAME9992(G9992,G9991,G9779);
  nand GNAME9993(G9993,G9992,G8790);
  nand GNAME9994(G9994,G9993,G9954,G8877);
  nand GNAME9995(G9995,G8822,G59426,G8795);
  nand GNAME9996(G9996,G8788,G8790);
  nand GNAME9997(G9997,G9995,G9996);
  nand GNAME9998(G9998,G8789,G9997);
  nand GNAME9999(G9999,G8801,G9994);
  and GNAME10000(G10000,G9998,G9999);
  or GNAME10001(G10001,G9104,G10000);
  nand GNAME10002(G10002,G9990,G59796);
  nand GNAME10003(G10003,G59426,G22263,G8795,G8822);
  nand GNAME10004(G10004,G9990,G59795);
  and GNAME10005(G10005,G59394,G59393);
  nand GNAME10006(G10006,G13985,G59792);
  and GNAME10007(G10007,G59393,G59758);
  or GNAME10008(G10008,G10007,G8831);
  or GNAME10009(G10009,G8830,G8832);
  nand GNAME10010(G10010,G13985,G59791);
  nand GNAME10011(G10011,G13985,G59790);
  not GNAME10012(G10012,G8842);
  not GNAME10013(G10013,G8835);
  nand GNAME10014(G10014,G8836,G8827,G8835);
  nand GNAME10015(G10015,G21700,G8842,G59427);
  nand GNAME10016(G10016,G10013,G8827,G8836,G9282);
  or GNAME10017(G10017,G8814,G21700,G10012);
  nand GNAME10018(G10018,G10016,G10017);
  nand GNAME10019(G10019,G9977,G8835);
  nand GNAME10020(G10020,G8827,G8838,G10013);
  nand GNAME10021(G10021,G10019,G8797);
  nand GNAME10022(G10022,G10020,G10021);
  nand GNAME10023(G10023,G8837,G59757);
  nand GNAME10024(G10024,G10018,G21700);
  nand GNAME10025(G10025,G59630,G8840);
  nand GNAME10026(G10026,G8843,G21998);
  nand GNAME10027(G10027,G22411,G8841);
  nand GNAME10028(G10028,G10012,G59789);
  nand GNAME10029(G10029,G8837,G59756);
  nand GNAME10030(G10030,G10018,G21632);
  nand GNAME10031(G10031,G8840,G59629);
  nand GNAME10032(G10032,G8843,G21937);
  nand GNAME10033(G10033,G8841,G22412);
  nand GNAME10034(G10034,G10012,G59788);
  nand GNAME10035(G10035,G8837,G59755);
  nand GNAME10036(G10036,G10018,G21686);
  nand GNAME10037(G10037,G8840,G59628);
  nand GNAME10038(G10038,G8843,G21985);
  nand GNAME10039(G10039,G8841,G22450);
  nand GNAME10040(G10040,G10012,G59787);
  nand GNAME10041(G10041,G8837,G59754);
  nand GNAME10042(G10042,G10018,G21687);
  nand GNAME10043(G10043,G8840,G59627);
  nand GNAME10044(G10044,G8843,G21986);
  nand GNAME10045(G10045,G8841,G22451);
  nand GNAME10046(G10046,G10012,G59786);
  nand GNAME10047(G10047,G8837,G59753);
  nand GNAME10048(G10048,G10018,G21688);
  nand GNAME10049(G10049,G8840,G59626);
  nand GNAME10050(G10050,G8843,G21987);
  nand GNAME10051(G10051,G8841,G22452);
  nand GNAME10052(G10052,G10012,G59785);
  nand GNAME10053(G10053,G8837,G59752);
  nand GNAME10054(G10054,G10018,G21689);
  nand GNAME10055(G10055,G8840,G59625);
  nand GNAME10056(G10056,G8843,G21988);
  nand GNAME10057(G10057,G8841,G22453);
  nand GNAME10058(G10058,G10012,G59784);
  nand GNAME10059(G10059,G8837,G59751);
  nand GNAME10060(G10060,G10018,G21690);
  nand GNAME10061(G10061,G8840,G59624);
  nand GNAME10062(G10062,G8843,G21989);
  nand GNAME10063(G10063,G8841,G22454);
  nand GNAME10064(G10064,G10012,G59783);
  nand GNAME10065(G10065,G8837,G59750);
  nand GNAME10066(G10066,G10018,G21691);
  nand GNAME10067(G10067,G8840,G59623);
  nand GNAME10068(G10068,G8843,G22027);
  nand GNAME10069(G10069,G8841,G22455);
  nand GNAME10070(G10070,G10012,G59782);
  nand GNAME10071(G10071,G8837,G59749);
  nand GNAME10072(G10072,G10018,G21692);
  nand GNAME10073(G10073,G8840,G59622);
  nand GNAME10074(G10074,G8843,G22030);
  nand GNAME10075(G10075,G8841,G22456);
  nand GNAME10076(G10076,G10012,G59781);
  nand GNAME10077(G10077,G8837,G59748);
  nand GNAME10078(G10078,G10018,G21693);
  nand GNAME10079(G10079,G8840,G59621);
  nand GNAME10080(G10080,G8843,G22033);
  nand GNAME10081(G10081,G8841,G22457);
  nand GNAME10082(G10082,G10012,G59780);
  nand GNAME10083(G10083,G8837,G59747);
  nand GNAME10084(G10084,G10018,G21694);
  nand GNAME10085(G10085,G8840,G59620);
  nand GNAME10086(G10086,G8843,G22036);
  nand GNAME10087(G10087,G8841,G22458);
  nand GNAME10088(G10088,G10012,G59779);
  nand GNAME10089(G10089,G8837,G59746);
  nand GNAME10090(G10090,G10018,G21695);
  nand GNAME10091(G10091,G8840,G59619);
  nand GNAME10092(G10092,G8843,G22039);
  nand GNAME10093(G10093,G8841,G22459);
  nand GNAME10094(G10094,G10012,G59778);
  nand GNAME10095(G10095,G8842,G8787,G8814);
  nand GNAME10096(G10096,G8837,G59745);
  nand GNAME10097(G10097,G10018,G21696);
  nand GNAME10098(G10098,G8840,G59618);
  nand GNAME10099(G10099,G8843,G22045);
  nand GNAME10100(G10100,G8841,G22463);
  nand GNAME10101(G10101,G10012,G59777);
  nand GNAME10102(G10102,G8837,G59744);
  nand GNAME10103(G10103,G10018,G21697);
  nand GNAME10104(G10104,G8840,G59617);
  nand GNAME10105(G10105,G8843,G22048);
  nand GNAME10106(G10106,G8841,G22464);
  nand GNAME10107(G10107,G10012,G59776);
  nand GNAME10108(G10108,G8837,G59743);
  nand GNAME10109(G10109,G10018,G21698);
  nand GNAME10110(G10110,G8840,G59616);
  nand GNAME10111(G10111,G8843,G22051);
  nand GNAME10112(G10112,G8841,G22465);
  nand GNAME10113(G10113,G10012,G59775);
  nand GNAME10114(G10114,G8837,G59742);
  nand GNAME10115(G10115,G10018,G21726);
  nand GNAME10116(G10116,G8840,G59615);
  nand GNAME10117(G10117,G8843,G21990);
  nand GNAME10118(G10118,G8841,G22466);
  nand GNAME10119(G10119,G10012,G59774);
  nand GNAME10120(G10120,G8837,G59741);
  nand GNAME10121(G10121,G10018,G21729);
  nand GNAME10122(G10122,G8840,G59614);
  nand GNAME10123(G10123,G8843,G21991);
  nand GNAME10124(G10124,G8841,G22467);
  nand GNAME10125(G10125,G10012,G59773);
  nand GNAME10126(G10126,G8837,G59740);
  nand GNAME10127(G10127,G10018,G21701);
  nand GNAME10128(G10128,G8840,G59613);
  nand GNAME10129(G10129,G8843,G21935);
  nand GNAME10130(G10130,G8841,G22413);
  nand GNAME10131(G10131,G10012,G59772);
  nand GNAME10132(G10132,G8837,G59739);
  nand GNAME10133(G10133,G10018,G21733);
  nand GNAME10134(G10134,G8840,G59612);
  nand GNAME10135(G10135,G8843,G21992);
  nand GNAME10136(G10136,G8841,G22468);
  nand GNAME10137(G10137,G10012,G59771);
  nand GNAME10138(G10138,G8837,G59738);
  nand GNAME10139(G10139,G10018,G21736);
  nand GNAME10140(G10140,G8840,G59611);
  nand GNAME10141(G10141,G8843,G21993);
  nand GNAME10142(G10142,G8841,G22469);
  nand GNAME10143(G10143,G10012,G59770);
  nand GNAME10144(G10144,G8837,G59737);
  nand GNAME10145(G10145,G10018,G21702);
  nand GNAME10146(G10146,G8840,G59610);
  nand GNAME10147(G10147,G8843,G21994);
  nand GNAME10148(G10148,G8841,G22349);
  nand GNAME10149(G10149,G10012,G59769);
  nand GNAME10150(G10150,G8837,G59736);
  nand GNAME10151(G10151,G10018,G21630);
  nand GNAME10152(G10152,G8840,G59609);
  nand GNAME10153(G10153,G8843,G21934);
  nand GNAME10154(G10154,G8841,G22348);
  nand GNAME10155(G10155,G10012,G59768);
  nand GNAME10156(G10156,G8837,G59735);
  nand GNAME10157(G10157,G10018,G21709);
  nand GNAME10158(G10158,G8840,G59608);
  nand GNAME10159(G10159,G8843,G21971);
  nand GNAME10160(G10160,G8841,G22440);
  nand GNAME10161(G10161,G10012,G59767);
  nand GNAME10162(G10162,G8837,G59734);
  nand GNAME10163(G10163,G10018,G21666);
  nand GNAME10164(G10164,G8840,G59607);
  nand GNAME10165(G10165,G8843,G22006);
  nand GNAME10166(G10166,G8841,G22441);
  nand GNAME10167(G10167,G10012,G59766);
  nand GNAME10168(G10168,G8837,G59733);
  nand GNAME10169(G10169,G10018,G21667);
  nand GNAME10170(G10170,G8840,G59606);
  nand GNAME10171(G10171,G8843,G21996);
  nand GNAME10172(G10172,G8841,G22409);
  nand GNAME10173(G10173,G10012,G59765);
  nand GNAME10174(G10174,G8837,G59732);
  nand GNAME10175(G10175,G10018,G21633);
  nand GNAME10176(G10176,G8840,G59605);
  nand GNAME10177(G10177,G8843,G21938);
  nand GNAME10178(G10178,G8841,G22351);
  nand GNAME10179(G10179,G10012,G59764);
  and GNAME10180(G10180,G8836,G8796,G8782);
  or GNAME10181(G10181,G10180,G8843);
  and GNAME10182(G10182,G8820,G8782,G8842);
  or GNAME10183(G10183,G10182,G8841);
  nand GNAME10184(G10184,G8837,G59731);
  nand GNAME10185(G10185,G10018,G21668);
  nand GNAME10186(G10186,G10183,G22445);
  nand GNAME10187(G10187,G8840,G59604);
  nand GNAME10188(G10188,G10181,G22010);
  nand GNAME10189(G10189,G10012,G59763);
  nand GNAME10190(G10190,G8837,G59730);
  nand GNAME10191(G10191,G10018,G21669);
  nand GNAME10192(G10192,G10183,G22448);
  nand GNAME10193(G10193,G8840,G59603);
  nand GNAME10194(G10194,G10181,G22013);
  nand GNAME10195(G10195,G10012,G59762);
  nand GNAME10196(G10196,G8837,G59729);
  nand GNAME10197(G10197,G10018,G21670);
  nand GNAME10198(G10198,G10183,G22410);
  nand GNAME10199(G10199,G8840,G59602);
  nand GNAME10200(G10200,G10012,G59761);
  nand GNAME10201(G10201,G10181,G21997);
  nand GNAME10202(G10202,G8837,G59728);
  nand GNAME10203(G10203,G10018,G21631);
  nand GNAME10204(G10204,G10183,G22350);
  nand GNAME10205(G10205,G8840,G59601);
  nand GNAME10206(G10206,G10012,G59760);
  nand GNAME10207(G10207,G10181,G21936);
  nand GNAME10208(G10208,G8837,G59727);
  nand GNAME10209(G10209,G10018,G21723);
  nand GNAME10210(G10210,G10183,G22462);
  nand GNAME10211(G10211,G8840,G59600);
  nand GNAME10212(G10212,G10181,G22042);
  nand GNAME10213(G10213,G59759,G10012);
  nand GNAME10214(G10214,G8837,G59726);
  nand GNAME10215(G10215,G10018,G21699);
  nand GNAME10216(G10216,G10183,G22408);
  nand GNAME10217(G10217,G8840,G59599);
  nand GNAME10218(G10218,G10181,G21995);
  nand GNAME10219(G10219,G59758,G10012);
  not GNAME10220(G10220,G8855);
  nand GNAME10221(G10221,G59428,G10220);
  nand GNAME10222(G10222,G21598,G8856);
  nand GNAME10223(G10223,G10221,G10222);
  nand GNAME10224(G10224,G8857,G59757);
  nand GNAME10225(G10225,G21700,G8858);
  nand GNAME10226(G10226,G8857,G59756);
  nand GNAME10227(G10227,G21937,G8859);
  nand GNAME10228(G10228,G21632,G8858);
  nand GNAME10229(G10229,G8857,G59755);
  nand GNAME10230(G10230,G21985,G8859);
  nand GNAME10231(G10231,G21686,G8858);
  nand GNAME10232(G10232,G8857,G59754);
  nand GNAME10233(G10233,G21986,G8859);
  nand GNAME10234(G10234,G21687,G8858);
  nand GNAME10235(G10235,G8857,G59753);
  nand GNAME10236(G10236,G21987,G8859);
  nand GNAME10237(G10237,G21688,G8858);
  nand GNAME10238(G10238,G8857,G59752);
  nand GNAME10239(G10239,G21988,G8859);
  nand GNAME10240(G10240,G21689,G8858);
  nand GNAME10241(G10241,G8857,G59751);
  nand GNAME10242(G10242,G21989,G8859);
  nand GNAME10243(G10243,G21690,G8858);
  nand GNAME10244(G10244,G8857,G59750);
  nand GNAME10245(G10245,G22027,G8859);
  nand GNAME10246(G10246,G21691,G8858);
  nand GNAME10247(G10247,G8857,G59749);
  nand GNAME10248(G10248,G22030,G8859);
  nand GNAME10249(G10249,G21692,G8858);
  nand GNAME10250(G10250,G8857,G59748);
  nand GNAME10251(G10251,G22033,G8859);
  nand GNAME10252(G10252,G21693,G8858);
  nand GNAME10253(G10253,G8857,G59747);
  nand GNAME10254(G10254,G22036,G8859);
  nand GNAME10255(G10255,G21694,G8858);
  nand GNAME10256(G10256,G8857,G59746);
  nand GNAME10257(G10257,G22039,G8859);
  nand GNAME10258(G10258,G21695,G8858);
  nand GNAME10259(G10259,G8857,G59745);
  nand GNAME10260(G10260,G22045,G8859);
  nand GNAME10261(G10261,G21696,G8858);
  nand GNAME10262(G10262,G8857,G59744);
  nand GNAME10263(G10263,G22048,G8859);
  nand GNAME10264(G10264,G21697,G8858);
  nand GNAME10265(G10265,G8857,G59743);
  nand GNAME10266(G10266,G22051,G8859);
  nand GNAME10267(G10267,G21698,G8858);
  nand GNAME10268(G10268,G8857,G59742);
  nand GNAME10269(G10269,G21990,G8859);
  nand GNAME10270(G10270,G21726,G8858);
  nand GNAME10271(G10271,G8857,G59741);
  nand GNAME10272(G10272,G21991,G8859);
  nand GNAME10273(G10273,G21729,G8858);
  nand GNAME10274(G10274,G8857,G59740);
  nand GNAME10275(G10275,G21935,G8859);
  nand GNAME10276(G10276,G21701,G8858);
  nand GNAME10277(G10277,G8857,G59739);
  nand GNAME10278(G10278,G21992,G8859);
  nand GNAME10279(G10279,G21733,G8858);
  nand GNAME10280(G10280,G8857,G59738);
  nand GNAME10281(G10281,G21993,G8859);
  nand GNAME10282(G10282,G21736,G8858);
  nand GNAME10283(G10283,G8857,G59737);
  nand GNAME10284(G10284,G21994,G8859);
  nand GNAME10285(G10285,G21702,G8858);
  nand GNAME10286(G10286,G8857,G59736);
  nand GNAME10287(G10287,G21934,G8859);
  nand GNAME10288(G10288,G21630,G8858);
  nand GNAME10289(G10289,G8857,G59735);
  nand GNAME10290(G10290,G21971,G8859);
  nand GNAME10291(G10291,G21709,G8858);
  nand GNAME10292(G10292,G8857,G59734);
  nand GNAME10293(G10293,G22006,G8859);
  nand GNAME10294(G10294,G21666,G8858);
  nand GNAME10295(G10295,G8857,G59733);
  nand GNAME10296(G10296,G21996,G8859);
  nand GNAME10297(G10297,G21667,G8858);
  nand GNAME10298(G10298,G8857,G59732);
  nand GNAME10299(G10299,G21938,G8859);
  nand GNAME10300(G10300,G21633,G8858);
  nand GNAME10301(G10301,G8857,G59731);
  nand GNAME10302(G10302,G22010,G8859);
  nand GNAME10303(G10303,G21668,G8858);
  nand GNAME10304(G10304,G8857,G59730);
  nand GNAME10305(G10305,G22013,G8859);
  nand GNAME10306(G10306,G21669,G8858);
  nand GNAME10307(G10307,G8857,G59729);
  nand GNAME10308(G10308,G21670,G8858);
  nand GNAME10309(G10309,G21997,G8859);
  nand GNAME10310(G10310,G8857,G59728);
  nand GNAME10311(G10311,G21631,G8858);
  nand GNAME10312(G10312,G21936,G8859);
  nand GNAME10313(G10313,G8857,G59727);
  nand GNAME10314(G10314,G22042,G8859);
  nand GNAME10315(G10315,G21723,G8858);
  nand GNAME10316(G10316,G8857,G59726);
  nand GNAME10317(G10317,G21699,G8858);
  nand GNAME10318(G10318,G21995,G8859);
  not GNAME10319(G10319,G8861);
  not GNAME10320(G10320,G9244);
  not GNAME10321(G10321,G8862);
  or GNAME10322(G10322,G8801,G8863);
  nand GNAME10323(G10323,G8788,G22263);
  nand GNAME10324(G10324,G10322,G10323);
  nand GNAME10325(G10325,G8749,G10324);
  nand GNAME10326(G10326,G21598,G8864);
  nand GNAME10327(G10327,G10326,G10320,G10325);
  nand GNAME10328(G10328,G8865,G59725);
  nand GNAME10329(G10329,G21700,G8866);
  nand GNAME10330(G10330,G8867,G1635);
  nand GNAME10331(G10331,G1654,G8868);
  nand GNAME10332(G10332,G8865,G59724);
  nand GNAME10333(G10333,G21632,G8866);
  nand GNAME10334(G10334,G22412,G8869);
  nand GNAME10335(G10335,G8867,G1636);
  nand GNAME10336(G10336,G8868,G1655);
  nand GNAME10337(G10337,G8865,G59723);
  nand GNAME10338(G10338,G21686,G8866);
  nand GNAME10339(G10339,G22450,G8869);
  nand GNAME10340(G10340,G8867,G1638);
  nand GNAME10341(G10341,G8868,G1656);
  nand GNAME10342(G10342,G8865,G59722);
  nand GNAME10343(G10343,G21687,G8866);
  nand GNAME10344(G10344,G22451,G8869);
  nand GNAME10345(G10345,G8867,G1639);
  nand GNAME10346(G10346,G8868,G1657);
  nand GNAME10347(G10347,G8865,G59721);
  nand GNAME10348(G10348,G21688,G8866);
  nand GNAME10349(G10349,G22452,G8869);
  nand GNAME10350(G10350,G8867,G1640);
  nand GNAME10351(G10351,G8868,G1658);
  nand GNAME10352(G10352,G8865,G59720);
  nand GNAME10353(G10353,G21689,G8866);
  nand GNAME10354(G10354,G22453,G8869);
  nand GNAME10355(G10355,G8867,G1641);
  nand GNAME10356(G10356,G8868,G1628);
  nand GNAME10357(G10357,G8865,G59719);
  nand GNAME10358(G10358,G21690,G8866);
  nand GNAME10359(G10359,G22454,G8869);
  nand GNAME10360(G10360,G8867,G1642);
  nand GNAME10361(G10361,G8868,G1629);
  nand GNAME10362(G10362,G8865,G59718);
  nand GNAME10363(G10363,G21691,G8866);
  nand GNAME10364(G10364,G22455,G8869);
  nand GNAME10365(G10365,G8867,G1643);
  nand GNAME10366(G10366,G8865,G59717);
  nand GNAME10367(G10367,G21692,G8866);
  nand GNAME10368(G10368,G22456,G8869);
  nand GNAME10369(G10369,G8867,G1644);
  nand GNAME10370(G10370,G8868,G1630);
  nand GNAME10371(G10371,G8865,G59716);
  nand GNAME10372(G10372,G21693,G8866);
  nand GNAME10373(G10373,G22457,G8869);
  nand GNAME10374(G10374,G8867,G1645);
  nand GNAME10375(G10375,G8868,G1631);
  nand GNAME10376(G10376,G8865,G59715);
  nand GNAME10377(G10377,G21694,G8866);
  nand GNAME10378(G10378,G22458,G8869);
  nand GNAME10379(G10379,G8867,G1646);
  nand GNAME10380(G10380,G8868,G1632);
  nand GNAME10381(G10381,G8865,G59714);
  nand GNAME10382(G10382,G21695,G8866);
  nand GNAME10383(G10383,G22459,G8869);
  nand GNAME10384(G10384,G8867,G1647);
  nand GNAME10385(G10385,G8868,G1633);
  nand GNAME10386(G10386,G8865,G59713);
  nand GNAME10387(G10387,G21696,G8866);
  nand GNAME10388(G10388,G22463,G8869);
  nand GNAME10389(G10389,G8867,G1649);
  nand GNAME10390(G10390,G8868,G1634);
  nand GNAME10391(G10391,G8865,G59712);
  nand GNAME10392(G10392,G21697,G8866);
  nand GNAME10393(G10393,G22464,G8869);
  nand GNAME10394(G10394,G8867,G1650);
  nand GNAME10395(G10395,G8868,G1637);
  nand GNAME10396(G10396,G8865,G59711);
  nand GNAME10397(G10397,G21698,G8866);
  nand GNAME10398(G10398,G22465,G8869);
  nand GNAME10399(G10399,G8867,G1651);
  nand GNAME10400(G10400,G8868,G1648);
  nand GNAME10401(G10401,G8865,G59710);
  nand GNAME10402(G10402,G21726,G8866);
  nand GNAME10403(G10403,G22466,G8869);
  nand GNAME10404(G10404,G8867,G1652);
  nand GNAME10405(G10405,G8868,G1659);
  nand GNAME10406(G10406,G1653,G8870);
  nand GNAME10407(G10407,G8865,G59709);
  nand GNAME10408(G10408,G21729,G8866);
  nand GNAME10409(G10409,G22467,G8869);
  nand GNAME10410(G10410,G1654,G8870);
  nand GNAME10411(G10411,G8865,G59708);
  nand GNAME10412(G10412,G21701,G8866);
  nand GNAME10413(G10413,G22413,G8869);
  nand GNAME10414(G10414,G1655,G8870);
  nand GNAME10415(G10415,G8865,G59707);
  nand GNAME10416(G10416,G21733,G8866);
  nand GNAME10417(G10417,G22468,G8869);
  nand GNAME10418(G10418,G1656,G8870);
  nand GNAME10419(G10419,G8865,G59706);
  nand GNAME10420(G10420,G21736,G8866);
  nand GNAME10421(G10421,G22469,G8869);
  nand GNAME10422(G10422,G1657,G8870);
  nand GNAME10423(G10423,G8865,G59705);
  nand GNAME10424(G10424,G21702,G8866);
  nand GNAME10425(G10425,G22349,G8869);
  nand GNAME10426(G10426,G1658,G8870);
  nand GNAME10427(G10427,G8865,G59704);
  nand GNAME10428(G10428,G21630,G8866);
  nand GNAME10429(G10429,G22348,G8869);
  nand GNAME10430(G10430,G1628,G8870);
  nand GNAME10431(G10431,G8865,G59703);
  nand GNAME10432(G10432,G21709,G8866);
  nand GNAME10433(G10433,G22440,G8869);
  nand GNAME10434(G10434,G1629,G8870);
  nand GNAME10435(G10435,G8865,G59702);
  nand GNAME10436(G10436,G21666,G8866);
  nand GNAME10437(G10437,G22441,G8869);
  nand GNAME10438(G10438,G8865,G59701);
  nand GNAME10439(G10439,G21667,G8866);
  nand GNAME10440(G10440,G22409,G8869);
  nand GNAME10441(G10441,G1630,G8870);
  nand GNAME10442(G10442,G8865,G59700);
  nand GNAME10443(G10443,G21633,G8866);
  nand GNAME10444(G10444,G22351,G8869);
  nand GNAME10445(G10445,G1631,G8870);
  nand GNAME10446(G10446,G8865,G59699);
  nand GNAME10447(G10447,G21668,G8866);
  nand GNAME10448(G10448,G22445,G8869);
  nand GNAME10449(G10449,G1632,G8870);
  nand GNAME10450(G10450,G8865,G59698);
  nand GNAME10451(G10451,G21669,G8866);
  nand GNAME10452(G10452,G22448,G8869);
  nand GNAME10453(G10453,G1633,G8870);
  nand GNAME10454(G10454,G8865,G59697);
  nand GNAME10455(G10455,G22410,G8869);
  nand GNAME10456(G10456,G21670,G8866);
  nand GNAME10457(G10457,G1634,G8870);
  nand GNAME10458(G10458,G8865,G59696);
  nand GNAME10459(G10459,G22350,G8869);
  nand GNAME10460(G10460,G21631,G8866);
  nand GNAME10461(G10461,G1637,G8870);
  nand GNAME10462(G10462,G8865,G59695);
  nand GNAME10463(G10463,G22462,G8869);
  nand GNAME10464(G10464,G21723,G8866);
  nand GNAME10465(G10465,G1648,G8870);
  nand GNAME10466(G10466,G8865,G59694);
  nand GNAME10467(G10467,G22408,G8869);
  nand GNAME10468(G10468,G21699,G8866);
  nand GNAME10469(G10469,G1659,G8870);
  not GNAME10470(G10470,G8871);
  nand GNAME10471(G10471,G8871,G59428,G9977);
  or GNAME10472(G10472,G59392,G8872);
  nand GNAME10473(G10473,G10471,G10472);
  nand GNAME10474(G10474,G21598,G10473,G8790);
  nand GNAME10475(G10475,G8873,G59692);
  nand GNAME10476(G10476,G59647,G8874);
  nand GNAME10477(G10477,G59724,G8876);
  nand GNAME10478(G10478,G8873,G59691);
  nand GNAME10479(G10479,G8874,G59648);
  nand GNAME10480(G10480,G59723,G8876);
  nand GNAME10481(G10481,G8873,G59690);
  nand GNAME10482(G10482,G8874,G59649);
  nand GNAME10483(G10483,G59722,G8876);
  nand GNAME10484(G10484,G8873,G59689);
  nand GNAME10485(G10485,G8874,G59650);
  nand GNAME10486(G10486,G59721,G8876);
  nand GNAME10487(G10487,G8873,G59688);
  nand GNAME10488(G10488,G8874,G59651);
  nand GNAME10489(G10489,G59720,G8876);
  nand GNAME10490(G10490,G8873,G59687);
  nand GNAME10491(G10491,G8874,G59652);
  nand GNAME10492(G10492,G59719,G8876);
  nand GNAME10493(G10493,G8873,G59686);
  nand GNAME10494(G10494,G8874,G59653);
  nand GNAME10495(G10495,G59718,G8876);
  nand GNAME10496(G10496,G8873,G59685);
  nand GNAME10497(G10497,G8874,G59654);
  nand GNAME10498(G10498,G59717,G8876);
  nand GNAME10499(G10499,G8873,G59684);
  nand GNAME10500(G10500,G8874,G59655);
  nand GNAME10501(G10501,G59716,G8876);
  nand GNAME10502(G10502,G8873,G59683);
  nand GNAME10503(G10503,G8874,G59656);
  nand GNAME10504(G10504,G59715,G8876);
  nand GNAME10505(G10505,G8873,G59682);
  nand GNAME10506(G10506,G8874,G59657);
  nand GNAME10507(G10507,G59714,G8876);
  nand GNAME10508(G10508,G8873,G59681);
  nand GNAME10509(G10509,G8874,G59658);
  nand GNAME10510(G10510,G59713,G8876);
  nand GNAME10511(G10511,G8873,G59680);
  nand GNAME10512(G10512,G8874,G59659);
  nand GNAME10513(G10513,G59712,G8876);
  nand GNAME10514(G10514,G8873,G59679);
  nand GNAME10515(G10515,G8874,G59660);
  nand GNAME10516(G10516,G59711,G8876);
  nand GNAME10517(G10517,G8873,G59678);
  nand GNAME10518(G10518,G8874,G59661);
  nand GNAME10519(G10519,G59710,G8876);
  nand GNAME10520(G10520,G8873,G59677);
  nand GNAME10521(G10521,G8874,G59631);
  nand GNAME10522(G10522,G59709,G8875);
  nand GNAME10523(G10523,G8873,G59676);
  nand GNAME10524(G10524,G8874,G59632);
  nand GNAME10525(G10525,G59708,G8875);
  nand GNAME10526(G10526,G8873,G59675);
  nand GNAME10527(G10527,G8874,G59633);
  nand GNAME10528(G10528,G59707,G8875);
  nand GNAME10529(G10529,G8873,G59674);
  nand GNAME10530(G10530,G8874,G59634);
  nand GNAME10531(G10531,G59706,G8875);
  nand GNAME10532(G10532,G8873,G59673);
  nand GNAME10533(G10533,G8874,G59635);
  nand GNAME10534(G10534,G59705,G8875);
  nand GNAME10535(G10535,G8873,G59672);
  nand GNAME10536(G10536,G8874,G59636);
  nand GNAME10537(G10537,G59704,G8875);
  nand GNAME10538(G10538,G8873,G59671);
  nand GNAME10539(G10539,G8874,G59637);
  nand GNAME10540(G10540,G59703,G8875);
  nand GNAME10541(G10541,G8873,G59670);
  nand GNAME10542(G10542,G8874,G59638);
  nand GNAME10543(G10543,G59702,G8875);
  nand GNAME10544(G10544,G8873,G59669);
  nand GNAME10545(G10545,G8874,G59639);
  nand GNAME10546(G10546,G59701,G8875);
  nand GNAME10547(G10547,G8873,G59668);
  nand GNAME10548(G10548,G8874,G59640);
  nand GNAME10549(G10549,G59700,G8875);
  nand GNAME10550(G10550,G8873,G59667);
  nand GNAME10551(G10551,G8874,G59641);
  nand GNAME10552(G10552,G59699,G8875);
  nand GNAME10553(G10553,G8873,G59666);
  nand GNAME10554(G10554,G8874,G59642);
  nand GNAME10555(G10555,G59698,G8875);
  nand GNAME10556(G10556,G8873,G59665);
  nand GNAME10557(G10557,G8874,G59643);
  nand GNAME10558(G10558,G59697,G8875);
  nand GNAME10559(G10559,G8873,G59664);
  nand GNAME10560(G10560,G8874,G59644);
  nand GNAME10561(G10561,G59696,G8875);
  nand GNAME10562(G10562,G8873,G59663);
  nand GNAME10563(G10563,G8874,G59645);
  nand GNAME10564(G10564,G59695,G8875);
  nand GNAME10565(G10565,G8873,G59662);
  nand GNAME10566(G10566,G8874,G59646);
  nand GNAME10567(G10567,G59694,G8875);
  or GNAME10568(G10568,G8801,G8877);
  or GNAME10569(G10569,G1588,G8878);
  nand GNAME10570(G10570,G59661,G8879);
  nand GNAME10571(G10571,G59710,G8880);
  nand GNAME10572(G10572,G59660,G8879);
  nand GNAME10573(G10573,G59711,G8880);
  nand GNAME10574(G10574,G59659,G8879);
  nand GNAME10575(G10575,G59712,G8880);
  nand GNAME10576(G10576,G59658,G8879);
  nand GNAME10577(G10577,G59713,G8880);
  nand GNAME10578(G10578,G59657,G8879);
  nand GNAME10579(G10579,G59714,G8880);
  nand GNAME10580(G10580,G59656,G8879);
  nand GNAME10581(G10581,G59715,G8880);
  nand GNAME10582(G10582,G59655,G8879);
  nand GNAME10583(G10583,G59716,G8880);
  nand GNAME10584(G10584,G59654,G8879);
  nand GNAME10585(G10585,G59717,G8880);
  nand GNAME10586(G10586,G59653,G8879);
  nand GNAME10587(G10587,G59718,G8880);
  nand GNAME10588(G10588,G59652,G8879);
  nand GNAME10589(G10589,G59719,G8880);
  nand GNAME10590(G10590,G59651,G8879);
  nand GNAME10591(G10591,G59720,G8880);
  nand GNAME10592(G10592,G59650,G8879);
  nand GNAME10593(G10593,G59721,G8880);
  nand GNAME10594(G10594,G59649,G8879);
  nand GNAME10595(G10595,G59722,G8880);
  nand GNAME10596(G10596,G59648,G8879);
  nand GNAME10597(G10597,G59723,G8880);
  nand GNAME10598(G10598,G59647,G8879);
  nand GNAME10599(G10599,G59724,G8880);
  nand GNAME10600(G10600,G59646,G8879);
  nand GNAME10601(G10601,G59694,G8880);
  nand GNAME10602(G10602,G1659,G8881);
  nand GNAME10603(G10603,G59645,G8879);
  nand GNAME10604(G10604,G59695,G8880);
  nand GNAME10605(G10605,G1648,G8881);
  nand GNAME10606(G10606,G59644,G8879);
  nand GNAME10607(G10607,G59696,G8880);
  nand GNAME10608(G10608,G1637,G8881);
  nand GNAME10609(G10609,G59643,G8879);
  nand GNAME10610(G10610,G59697,G8880);
  nand GNAME10611(G10611,G1634,G8881);
  nand GNAME10612(G10612,G59642,G8879);
  nand GNAME10613(G10613,G59698,G8880);
  nand GNAME10614(G10614,G1633,G8881);
  nand GNAME10615(G10615,G59641,G8879);
  nand GNAME10616(G10616,G59699,G8880);
  nand GNAME10617(G10617,G1632,G8881);
  nand GNAME10618(G10618,G59640,G8879);
  nand GNAME10619(G10619,G59700,G8880);
  nand GNAME10620(G10620,G1631,G8881);
  nand GNAME10621(G10621,G59639,G8879);
  nand GNAME10622(G10622,G59701,G8880);
  nand GNAME10623(G10623,G1630,G8881);
  nand GNAME10624(G10624,G1629,G8881);
  nand GNAME10625(G10625,G59638,G8879);
  nand GNAME10626(G10626,G59702,G8880);
  nand GNAME10627(G10627,G1628,G8881);
  nand GNAME10628(G10628,G59637,G8879);
  nand GNAME10629(G10629,G59703,G8880);
  nand GNAME10630(G10630,G1658,G8881);
  nand GNAME10631(G10631,G59636,G8879);
  nand GNAME10632(G10632,G59704,G8880);
  nand GNAME10633(G10633,G1657,G8881);
  nand GNAME10634(G10634,G59635,G8879);
  nand GNAME10635(G10635,G59705,G8880);
  nand GNAME10636(G10636,G1656,G8881);
  nand GNAME10637(G10637,G59634,G8879);
  nand GNAME10638(G10638,G59706,G8880);
  nand GNAME10639(G10639,G1655,G8881);
  nand GNAME10640(G10640,G59633,G8879);
  nand GNAME10641(G10641,G59707,G8880);
  nand GNAME10642(G10642,G1654,G8881);
  nand GNAME10643(G10643,G59632,G8879);
  nand GNAME10644(G10644,G59708,G8880);
  nand GNAME10645(G10645,G59631,G8879);
  nand GNAME10646(G10646,G1653,G8881);
  nand GNAME10647(G10647,G59709,G8880);
  nand GNAME10648(G10648,G8787,G8816);
  nand GNAME10649(G10649,G59630,G8882);
  nand GNAME10650(G10650,G21998,G8883);
  nand GNAME10651(G10651,G21700,G8884);
  nand GNAME10652(G10652,G22411,G8885);
  nand GNAME10653(G10653,G59789,G8886);
  nand GNAME10654(G10654,G59629,G8882);
  nand GNAME10655(G10655,G21937,G8883);
  nand GNAME10656(G10656,G21632,G8884);
  nand GNAME10657(G10657,G22412,G8885);
  nand GNAME10658(G10658,G59788,G8886);
  nand GNAME10659(G10659,G59628,G8882);
  nand GNAME10660(G10660,G21985,G8883);
  nand GNAME10661(G10661,G21686,G8884);
  nand GNAME10662(G10662,G22450,G8885);
  nand GNAME10663(G10663,G59787,G8886);
  nand GNAME10664(G10664,G59627,G8882);
  nand GNAME10665(G10665,G21986,G8883);
  nand GNAME10666(G10666,G21687,G8884);
  nand GNAME10667(G10667,G22451,G8885);
  nand GNAME10668(G10668,G59786,G8886);
  nand GNAME10669(G10669,G59626,G8882);
  nand GNAME10670(G10670,G21987,G8883);
  nand GNAME10671(G10671,G21688,G8884);
  nand GNAME10672(G10672,G22452,G8885);
  nand GNAME10673(G10673,G59785,G8886);
  nand GNAME10674(G10674,G59625,G8882);
  nand GNAME10675(G10675,G21988,G8883);
  nand GNAME10676(G10676,G21689,G8884);
  nand GNAME10677(G10677,G22453,G8885);
  nand GNAME10678(G10678,G59784,G8886);
  nand GNAME10679(G10679,G59624,G8882);
  nand GNAME10680(G10680,G21989,G8883);
  nand GNAME10681(G10681,G21690,G8884);
  nand GNAME10682(G10682,G22454,G8885);
  nand GNAME10683(G10683,G59783,G8886);
  nand GNAME10684(G10684,G59623,G8882);
  nand GNAME10685(G10685,G22027,G8883);
  nand GNAME10686(G10686,G21691,G8884);
  nand GNAME10687(G10687,G22455,G8885);
  nand GNAME10688(G10688,G59782,G8886);
  nand GNAME10689(G10689,G59622,G8882);
  nand GNAME10690(G10690,G22030,G8883);
  nand GNAME10691(G10691,G21692,G8884);
  nand GNAME10692(G10692,G22456,G8885);
  nand GNAME10693(G10693,G59781,G8886);
  nand GNAME10694(G10694,G59621,G8882);
  nand GNAME10695(G10695,G22033,G8883);
  nand GNAME10696(G10696,G21693,G8884);
  nand GNAME10697(G10697,G22457,G8885);
  nand GNAME10698(G10698,G59780,G8886);
  nand GNAME10699(G10699,G59620,G8882);
  nand GNAME10700(G10700,G22036,G8883);
  nand GNAME10701(G10701,G21694,G8884);
  nand GNAME10702(G10702,G22458,G8885);
  nand GNAME10703(G10703,G59779,G8886);
  nand GNAME10704(G10704,G59619,G8882);
  nand GNAME10705(G10705,G22039,G8883);
  nand GNAME10706(G10706,G21695,G8884);
  nand GNAME10707(G10707,G22459,G8885);
  nand GNAME10708(G10708,G59778,G8886);
  nand GNAME10709(G10709,G59618,G8882);
  nand GNAME10710(G10710,G22045,G8883);
  nand GNAME10711(G10711,G21696,G8884);
  nand GNAME10712(G10712,G22463,G8885);
  nand GNAME10713(G10713,G59777,G8886);
  nand GNAME10714(G10714,G59617,G8882);
  nand GNAME10715(G10715,G22048,G8883);
  nand GNAME10716(G10716,G21697,G8884);
  nand GNAME10717(G10717,G22464,G8885);
  nand GNAME10718(G10718,G59776,G8886);
  nand GNAME10719(G10719,G59616,G8882);
  nand GNAME10720(G10720,G22051,G8883);
  nand GNAME10721(G10721,G21698,G8884);
  nand GNAME10722(G10722,G22465,G8885);
  nand GNAME10723(G10723,G59775,G8886);
  nand GNAME10724(G10724,G59615,G8882);
  nand GNAME10725(G10725,G21990,G8883);
  nand GNAME10726(G10726,G21726,G8884);
  nand GNAME10727(G10727,G22466,G8885);
  nand GNAME10728(G10728,G59774,G8886);
  nand GNAME10729(G10729,G59614,G8882);
  nand GNAME10730(G10730,G21991,G8883);
  nand GNAME10731(G10731,G21729,G8884);
  nand GNAME10732(G10732,G22467,G8885);
  nand GNAME10733(G10733,G59773,G8886);
  nand GNAME10734(G10734,G59613,G8882);
  nand GNAME10735(G10735,G21935,G8883);
  nand GNAME10736(G10736,G21701,G8884);
  nand GNAME10737(G10737,G22413,G8885);
  nand GNAME10738(G10738,G59772,G8886);
  nand GNAME10739(G10739,G59612,G8882);
  nand GNAME10740(G10740,G21992,G8883);
  nand GNAME10741(G10741,G21733,G8884);
  nand GNAME10742(G10742,G22468,G8885);
  nand GNAME10743(G10743,G59771,G8886);
  nand GNAME10744(G10744,G59611,G8882);
  nand GNAME10745(G10745,G21993,G8883);
  nand GNAME10746(G10746,G21736,G8884);
  nand GNAME10747(G10747,G22469,G8885);
  nand GNAME10748(G10748,G59770,G8886);
  nand GNAME10749(G10749,G59610,G8882);
  nand GNAME10750(G10750,G21994,G8883);
  nand GNAME10751(G10751,G21702,G8884);
  nand GNAME10752(G10752,G22349,G8885);
  nand GNAME10753(G10753,G59769,G8886);
  nand GNAME10754(G10754,G59609,G8882);
  nand GNAME10755(G10755,G21934,G8883);
  nand GNAME10756(G10756,G21630,G8884);
  nand GNAME10757(G10757,G22348,G8885);
  nand GNAME10758(G10758,G59768,G8886);
  nand GNAME10759(G10759,G59608,G8882);
  nand GNAME10760(G10760,G21971,G8883);
  nand GNAME10761(G10761,G21709,G8884);
  nand GNAME10762(G10762,G22440,G8885);
  nand GNAME10763(G10763,G59767,G8886);
  nand GNAME10764(G10764,G59607,G8882);
  nand GNAME10765(G10765,G22006,G8883);
  nand GNAME10766(G10766,G21666,G8884);
  nand GNAME10767(G10767,G22441,G8885);
  nand GNAME10768(G10768,G59766,G8886);
  nand GNAME10769(G10769,G59606,G8882);
  nand GNAME10770(G10770,G21996,G8883);
  nand GNAME10771(G10771,G21667,G8884);
  nand GNAME10772(G10772,G22409,G8885);
  nand GNAME10773(G10773,G59765,G8886);
  nand GNAME10774(G10774,G59605,G8882);
  nand GNAME10775(G10775,G21938,G8883);
  nand GNAME10776(G10776,G21633,G8884);
  nand GNAME10777(G10777,G22351,G8885);
  nand GNAME10778(G10778,G59764,G8886);
  nand GNAME10779(G10779,G59604,G8882);
  nand GNAME10780(G10780,G22010,G8883);
  nand GNAME10781(G10781,G21668,G8884);
  nand GNAME10782(G10782,G22445,G8885);
  nand GNAME10783(G10783,G59763,G8886);
  nand GNAME10784(G10784,G59603,G8882);
  nand GNAME10785(G10785,G22013,G8883);
  nand GNAME10786(G10786,G21669,G8884);
  nand GNAME10787(G10787,G22448,G8885);
  nand GNAME10788(G10788,G59762,G8886);
  nand GNAME10789(G10789,G59602,G8882);
  nand GNAME10790(G10790,G22410,G8885);
  nand GNAME10791(G10791,G59761,G8886);
  nand GNAME10792(G10792,G21670,G8884);
  nand GNAME10793(G10793,G21997,G8883);
  nand GNAME10794(G10794,G59601,G8882);
  nand GNAME10795(G10795,G22350,G8885);
  nand GNAME10796(G10796,G59760,G8886);
  nand GNAME10797(G10797,G21631,G8884);
  nand GNAME10798(G10798,G21936,G8883);
  nand GNAME10799(G10799,G59600,G8882);
  nand GNAME10800(G10800,G22462,G8885);
  nand GNAME10801(G10801,G22042,G8883);
  nand GNAME10802(G10802,G21723,G8884);
  nand GNAME10803(G10803,G59759,G8886);
  nand GNAME10804(G10804,G59599,G8882);
  nand GNAME10805(G10805,G22408,G8885);
  nand GNAME10806(G10806,G21699,G8884);
  nand GNAME10807(G10807,G59758,G8886);
  nand GNAME10808(G10808,G21995,G8883);
  nand GNAME10809(G10809,G8780,G8784);
  nand GNAME10810(G10810,G9849,G8826);
  nand GNAME10811(G10811,G8783,G9849);
  nand GNAME10812(G10812,G10811,G8887);
  nand GNAME10813(G10813,G8783,G8782);
  nand GNAME10814(G10814,G9783,G9832);
  nand GNAME10815(G10815,G9900,G8749,G8796);
  nand GNAME10816(G10816,G10815,G9917);
  nand GNAME10817(G10817,G9832,G9977);
  nand GNAME10818(G10818,G10817,G9883);
  nand GNAME10819(G10819,G10818,G9849);
  nand GNAME10820(G10820,G8781,G9977);
  nand GNAME10821(G10821,G10819,G10820);
  nand GNAME10822(G10822,G8749,G10821);
  nand GNAME10823(G10823,G10822,G9900);
  nand GNAME10824(G10824,G22263,G10816,G9883);
  nand GNAME10825(G10825,G10823,G21598);
  nand GNAME10826(G10826,G8888,G10824,G10825);
  nand GNAME10827(G10827,G10826,G8800);
  nand GNAME10828(G10828,G8787,G8810);
  or GNAME10829(G10829,G8828,G8822,G8786,G10319);
  nand GNAME10830(G10830,G8891,G8783,G8797);
  or GNAME10831(G10831,G9900,G8750);
  nand GNAME10832(G10832,G10321,G10830,G10831,G8902);
  nand GNAME10833(G10833,G9249,G9934);
  nand GNAME10834(G10834,G8781,G8746);
  nand GNAME10835(G10835,G9900,G9781,G9951);
  nand GNAME10836(G10836,G10835,G9934);
  nand GNAME10837(G10837,G8781,G8823);
  nand GNAME10838(G10838,G9805,G8860);
  or GNAME10839(G10839,G8750,G8783);
  nand GNAME10840(G10840,G13970,G8853);
  nand GNAME10841(G10841,G10840,G9789);
  nand GNAME10842(G10842,G8792,G8896);
  nand GNAME10843(G10843,G9934,G8897);
  nand GNAME10844(G10844,G8899,G8900);
  nand GNAME10845(G10845,G22931,G8890);
  nand GNAME10846(G10846,G21998,G8901);
  nand GNAME10847(G10847,G21700,G8903);
  nand GNAME10848(G10848,G22411,G8904);
  nand GNAME10849(G10849,G59789,G8905);
  nand GNAME10850(G10850,G8906,G59598);
  nand GNAME10851(G10851,G8906,G59597);
  nand GNAME10852(G10852,G8890,G22932);
  nand GNAME10853(G10853,G21937,G8901);
  nand GNAME10854(G10854,G21632,G8903);
  nand GNAME10855(G10855,G22412,G8904);
  nand GNAME10856(G10856,G59788,G8905);
  nand GNAME10857(G10857,G8906,G59596);
  nand GNAME10858(G10858,G8890,G22883);
  nand GNAME10859(G10859,G21985,G8901);
  nand GNAME10860(G10860,G21686,G8903);
  nand GNAME10861(G10861,G22450,G8904);
  nand GNAME10862(G10862,G59787,G8905);
  nand GNAME10863(G10863,G8906,G59595);
  nand GNAME10864(G10864,G8890,G22882);
  nand GNAME10865(G10865,G21986,G8901);
  nand GNAME10866(G10866,G21687,G8903);
  nand GNAME10867(G10867,G22451,G8904);
  nand GNAME10868(G10868,G59786,G8905);
  nand GNAME10869(G10869,G8906,G59594);
  nand GNAME10870(G10870,G8890,G22934);
  nand GNAME10871(G10871,G21987,G8901);
  nand GNAME10872(G10872,G21688,G8903);
  nand GNAME10873(G10873,G22452,G8904);
  nand GNAME10874(G10874,G59785,G8905);
  nand GNAME10875(G10875,G8906,G59593);
  nand GNAME10876(G10876,G8890,G22881);
  nand GNAME10877(G10877,G21988,G8901);
  nand GNAME10878(G10878,G21689,G8903);
  nand GNAME10879(G10879,G22453,G8904);
  nand GNAME10880(G10880,G59784,G8905);
  nand GNAME10881(G10881,G8906,G59592);
  nand GNAME10882(G10882,G8890,G22880);
  nand GNAME10883(G10883,G21989,G8901);
  nand GNAME10884(G10884,G21690,G8903);
  nand GNAME10885(G10885,G22454,G8904);
  nand GNAME10886(G10886,G59783,G8905);
  nand GNAME10887(G10887,G8906,G59591);
  nand GNAME10888(G10888,G8890,G22958);
  nand GNAME10889(G10889,G22027,G8901);
  nand GNAME10890(G10890,G21691,G8903);
  nand GNAME10891(G10891,G22455,G8904);
  nand GNAME10892(G10892,G59782,G8905);
  nand GNAME10893(G10893,G8906,G59590);
  nand GNAME10894(G10894,G8890,G22959);
  nand GNAME10895(G10895,G22030,G8901);
  nand GNAME10896(G10896,G21692,G8903);
  nand GNAME10897(G10897,G22456,G8904);
  nand GNAME10898(G10898,G59781,G8905);
  nand GNAME10899(G10899,G8890,G22960);
  nand GNAME10900(G10900,G22033,G8901);
  nand GNAME10901(G10901,G21693,G8903);
  nand GNAME10902(G10902,G22457,G8904);
  nand GNAME10903(G10903,G59780,G8905);
  nand GNAME10904(G10904,G8906,G59589);
  nand GNAME10905(G10905,G8890,G22961);
  nand GNAME10906(G10906,G22036,G8901);
  nand GNAME10907(G10907,G21694,G8903);
  nand GNAME10908(G10908,G22458,G8904);
  nand GNAME10909(G10909,G59779,G8905);
  nand GNAME10910(G10910,G8906,G59588);
  nand GNAME10911(G10911,G8890,G22962);
  nand GNAME10912(G10912,G22039,G8901);
  nand GNAME10913(G10913,G21695,G8903);
  nand GNAME10914(G10914,G22459,G8904);
  nand GNAME10915(G10915,G59778,G8905);
  nand GNAME10916(G10916,G8906,G59587);
  nand GNAME10917(G10917,G8890,G22964);
  nand GNAME10918(G10918,G22045,G8901);
  nand GNAME10919(G10919,G21696,G8903);
  nand GNAME10920(G10920,G22463,G8904);
  nand GNAME10921(G10921,G59777,G8905);
  nand GNAME10922(G10922,G8906,G59586);
  nand GNAME10923(G10923,G8890,G22965);
  nand GNAME10924(G10924,G22048,G8901);
  nand GNAME10925(G10925,G21697,G8903);
  nand GNAME10926(G10926,G22464,G8904);
  nand GNAME10927(G10927,G59776,G8905);
  nand GNAME10928(G10928,G8906,G59585);
  nand GNAME10929(G10929,G8890,G22966);
  nand GNAME10930(G10930,G22051,G8901);
  nand GNAME10931(G10931,G21698,G8903);
  nand GNAME10932(G10932,G22465,G8904);
  nand GNAME10933(G10933,G59775,G8905);
  nand GNAME10934(G10934,G8906,G59584);
  nand GNAME10935(G10935,G8890,G22936);
  nand GNAME10936(G10936,G21990,G8901);
  nand GNAME10937(G10937,G21726,G8903);
  nand GNAME10938(G10938,G22466,G8904);
  nand GNAME10939(G10939,G59774,G8905);
  nand GNAME10940(G10940,G8906,G59583);
  nand GNAME10941(G10941,G8890,G22937);
  nand GNAME10942(G10942,G21991,G8901);
  nand GNAME10943(G10943,G21729,G8903);
  nand GNAME10944(G10944,G22467,G8904);
  nand GNAME10945(G10945,G59773,G8905);
  nand GNAME10946(G10946,G8906,G59582);
  nand GNAME10947(G10947,G8890,G22938);
  nand GNAME10948(G10948,G21935,G8901);
  nand GNAME10949(G10949,G21701,G8903);
  nand GNAME10950(G10950,G22413,G8904);
  nand GNAME10951(G10951,G59772,G8905);
  nand GNAME10952(G10952,G8906,G59581);
  nand GNAME10953(G10953,G8890,G22939);
  nand GNAME10954(G10954,G21992,G8901);
  nand GNAME10955(G10955,G21733,G8903);
  nand GNAME10956(G10956,G22468,G8904);
  nand GNAME10957(G10957,G59771,G8905);
  nand GNAME10958(G10958,G8906,G59580);
  nand GNAME10959(G10959,G8890,G22940);
  nand GNAME10960(G10960,G21993,G8901);
  nand GNAME10961(G10961,G21736,G8903);
  nand GNAME10962(G10962,G22469,G8904);
  nand GNAME10963(G10963,G59770,G8905);
  nand GNAME10964(G10964,G8906,G59579);
  nand GNAME10965(G10965,G8890,G22941);
  nand GNAME10966(G10966,G21994,G8901);
  nand GNAME10967(G10967,G21702,G8903);
  nand GNAME10968(G10968,G22349,G8904);
  nand GNAME10969(G10969,G59769,G8905);
  nand GNAME10970(G10970,G8906,G59578);
  nand GNAME10971(G10971,G8890,G22942);
  nand GNAME10972(G10972,G21934,G8901);
  nand GNAME10973(G10973,G21630,G8903);
  nand GNAME10974(G10974,G22348,G8904);
  nand GNAME10975(G10975,G59768,G8905);
  nand GNAME10976(G10976,G8906,G59577);
  nand GNAME10977(G10977,G8890,G22924);
  nand GNAME10978(G10978,G21971,G8901);
  nand GNAME10979(G10979,G21709,G8903);
  nand GNAME10980(G10980,G22440,G8904);
  nand GNAME10981(G10981,G59767,G8905);
  nand GNAME10982(G10982,G8906,G59576);
  nand GNAME10983(G10983,G8890,G22925);
  nand GNAME10984(G10984,G22006,G8901);
  nand GNAME10985(G10985,G21666,G8903);
  nand GNAME10986(G10986,G22441,G8904);
  nand GNAME10987(G10987,G59766,G8905);
  nand GNAME10988(G10988,G8906,G59575);
  nand GNAME10989(G10989,G8890,G22926);
  nand GNAME10990(G10990,G21996,G8901);
  nand GNAME10991(G10991,G21667,G8903);
  nand GNAME10992(G10992,G22409,G8904);
  nand GNAME10993(G10993,G59765,G8905);
  nand GNAME10994(G10994,G8906,G59574);
  nand GNAME10995(G10995,G8890,G22927);
  nand GNAME10996(G10996,G21938,G8901);
  nand GNAME10997(G10997,G21633,G8903);
  nand GNAME10998(G10998,G22351,G8904);
  nand GNAME10999(G10999,G59764,G8905);
  nand GNAME11000(G11000,G8906,G59573);
  nand GNAME11001(G11001,G8890,G22928);
  nand GNAME11002(G11002,G22010,G8901);
  nand GNAME11003(G11003,G21668,G8903);
  nand GNAME11004(G11004,G22445,G8904);
  nand GNAME11005(G11005,G59763,G8905);
  nand GNAME11006(G11006,G8906,G59572);
  nand GNAME11007(G11007,G8890,G22929);
  nand GNAME11008(G11008,G22013,G8901);
  nand GNAME11009(G11009,G21669,G8903);
  nand GNAME11010(G11010,G22448,G8904);
  nand GNAME11011(G11011,G59762,G8905);
  nand GNAME11012(G11012,G8906,G59571);
  nand GNAME11013(G11013,G8890,G22930);
  nand GNAME11014(G11014,G22410,G8904);
  nand GNAME11015(G11015,G59761,G8905);
  nand GNAME11016(G11016,G21670,G8903);
  nand GNAME11017(G11017,G21997,G8901);
  nand GNAME11018(G11018,G8906,G59570);
  nand GNAME11019(G11019,G8890,G22933);
  nand GNAME11020(G11020,G22350,G8904);
  nand GNAME11021(G11021,G59760,G8905);
  nand GNAME11022(G11022,G21631,G8903);
  nand GNAME11023(G11023,G21936,G8901);
  nand GNAME11024(G11024,G8906,G59569);
  nand GNAME11025(G11025,G8890,G22935);
  nand GNAME11026(G11026,G22462,G8904);
  nand GNAME11027(G11027,G22042,G8901);
  nand GNAME11028(G11028,G59759,G8905);
  nand GNAME11029(G11029,G21723,G8903);
  nand GNAME11030(G11030,G8906,G59568);
  nand GNAME11031(G11031,G8890,G22943);
  nand GNAME11032(G11032,G22408,G8904);
  nand GNAME11033(G11033,G59758,G8905);
  nand GNAME11034(G11034,G21995,G8901);
  nand GNAME11035(G11035,G21699,G8903);
  nand GNAME11036(G11036,G8906,G59567);
  or GNAME11037(G11037,G8801,G8909);
  not GNAME11038(G11038,G8910);
  or GNAME11039(G11039,G21598,G13984);
  not GNAME11040(G11040,G8917);
  nand GNAME11041(G11041,G59561,G8795);
  nor GNAME11042(G11042,G8785,G59427);
  nand GNAME11043(G11043,G8912,G8913);
  not GNAME11044(G11044,G8914);
  nand GNAME11045(G11045,G8751,G9796);
  nand GNAME11046(G11046,G11045,G9799);
  nand GNAME11047(G11047,G11044,G8915);
  nand GNAME11048(G11048,G21699,G8916);
  nand GNAME11049(G11049,G8907,G13867,G13868);
  nand GNAME11050(G11050,G8745,G8795);
  not GNAME11051(G11051,G8920);
  nand GNAME11052(G11052,G8751,G8952);
  nand GNAME11053(G11053,G59560,G8795);
  nand GNAME11054(G11054,G8813,G59565);
  not GNAME11055(G11055,G8921);
  nand GNAME11056(G11056,G9250,G8915);
  nand GNAME11057(G11057,G21723,G8916);
  nand GNAME11058(G11058,G11040,G59565);
  nand GNAME11059(G11059,G8751,G9251);
  nand GNAME11060(G11060,G59559,G8795);
  nand GNAME11061(G11061,G8813,G59564);
  nand GNAME11062(G11062,G8921,G9801);
  nand GNAME11063(G11063,G11062,G11051);
  nand GNAME11064(G11064,G8919,G11055);
  nand GNAME11065(G11065,G8925,G8924);
  not GNAME11066(G11066,G8926);
  nand GNAME11067(G11067,G8915,G11066);
  nand GNAME11068(G11068,G21631,G8916);
  nand GNAME11069(G11069,G11040,G59564);
  nor GNAME11070(G11070,G8923,G8928);
  nand GNAME11071(G11071,G8751,G8953);
  nand GNAME11072(G11072,G59558,G8795);
  nand GNAME11073(G11073,G8813,G59563);
  nand GNAME11074(G11074,G8915,G13879);
  nand GNAME11075(G11075,G21670,G8916);
  nand GNAME11076(G11076,G11040,G59563);
  nand GNAME11077(G11077,G10470,G8799);
  nand GNAME11078(G11078,G11077,G9977);
  nand GNAME11079(G11079,G11078,G10321);
  nand GNAME11080(G11080,G11079,G21598);
  nand GNAME11081(G11081,G8786,G22263);
  nand GNAME11082(G11082,G11080,G11081);
  nand GNAME11083(G11083,G8749,G11082);
  or GNAME11084(G11084,G9105,G8801);
  nand GNAME11085(G11085,G9778,G8800);
  nand GNAME11086(G11086,G9976,G8894);
  nand GNAME11087(G11087,G11086,G13455);
  nand GNAME11088(G11088,G8792,G59426);
  nand GNAME11089(G11089,G11088,G9775,G9802);
  not GNAME11090(G11090,G8930);
  nand GNAME11091(G11091,G8792,G11090);
  nand GNAME11092(G11092,G11091,G59426);
  nand GNAME11093(G11093,G8914,G8930);
  not GNAME11094(G11094,G8933);
  nand GNAME11095(G11095,G9866,G8930,G59426);
  not GNAME11096(G11096,G8931);
  nand GNAME11097(G11097,G8797,G8891);
  nand GNAME11098(G11098,G11097,G8750);
  nand GNAME11099(G11099,G8783,G11098);
  nand GNAME11100(G11100,G9866,G8896);
  nand GNAME11101(G11101,G8861,G10321,G11099,G11100);
  nand GNAME11102(G11102,G8796,G8821);
  nand GNAME11103(G11103,G11102,G8900);
  nand GNAME11104(G11104,G9952,G8898);
  nand GNAME11105(G11105,G8855,G10470);
  or GNAME11106(G11106,G59561,G9105);
  nand GNAME11107(G11107,G11105,G11096);
  nand GNAME11108(G11108,G11104,G11044);
  nand GNAME11109(G11109,G11103,G21699);
  nand GNAME11110(G11110,G11101,G21995);
  nand GNAME11111(G11111,G11109,G11110,G11108,G11106,G11107);
  nand GNAME11112(G11112,G8914,G13864);
  nand GNAME11113(G11113,G21995,G8929);
  nand GNAME11114(G11114,G11112,G59427);
  nand GNAME11115(G11115,G11111,G8790);
  nand GNAME11116(G11116,G11115,G11113,G11114);
  nand GNAME11117(G11117,G11089,G59560);
  nand GNAME11118(G11118,G8751,G9250);
  not GNAME11119(G11119,G8934);
  not GNAME11120(G11120,G9187);
  nand GNAME11121(G11121,G59561,G9866);
  not GNAME11122(G11122,G9161);
  or GNAME11123(G11123,G8754,G11122);
  nand GNAME11124(G11124,G11123,G8825);
  nand GNAME11125(G11125,G11105,G13886);
  nand GNAME11126(G11126,G11104,G9250);
  nand GNAME11127(G11127,G11103,G21723);
  nand GNAME11128(G11128,G11101,G22042);
  nand GNAME11129(G11129,G9187,G8828);
  nand GNAME11130(G11130,G9401,G11126,G11128,G11125);
  nand GNAME11131(G11131,G9250,G8932);
  nand GNAME11132(G11132,G22042,G8929);
  nand GNAME11133(G11133,G11130,G8790);
  nand GNAME11134(G11134,G11133,G11131,G11132);
  nand GNAME11135(G11135,G8934,G11094);
  nand GNAME11136(G11136,G9775,G11135);
  nand GNAME11137(G11137,G8933,G11119);
  not GNAME11138(G11138,G8936);
  nand GNAME11139(G11139,G11089,G59559);
  nand GNAME11140(G11140,G8751,G11066);
  not GNAME11141(G11141,G8935);
  nand GNAME11142(G11142,G9787,G9255);
  not GNAME11143(G11143,G8937);
  not GNAME11144(G11144,G9776);
  nand GNAME11145(G11145,G11105,G13892);
  nand GNAME11146(G11146,G11104,G11066);
  nand GNAME11147(G11147,G11103,G21631);
  nand GNAME11148(G11148,G11101,G21936);
  nand GNAME11149(G11149,G8825,G13898);
  nand GNAME11150(G11150,G8828,G11143);
  nand GNAME11151(G11151,G9402,G11147,G11145,G11148);
  nand GNAME11152(G11152,G11066,G8932);
  nand GNAME11153(G11153,G21936,G8929);
  nand GNAME11154(G11154,G11151,G8790);
  nand GNAME11155(G11155,G11154,G11152,G11153);
  nand GNAME11156(G11156,G11089,G59558);
  nand GNAME11157(G11157,G11156,G11162);
  nand GNAME11158(G11158,G11163,G11138);
  nand GNAME11159(G11159,G11160,G11157,G11158);
  nand GNAME11160(G11160,G8935,G8820);
  nand GNAME11161(G11161,G8936,G11160);
  nand GNAME11162(G11162,G8751,G13879);
  nand GNAME11163(G11163,G9802,G11141);
  nand GNAME11164(G11164,G11156,G11161,G11162,G11163);
  not GNAME11165(G11165,G8941);
  nand GNAME11166(G11166,G11144,G8753);
  nand GNAME11167(G11167,G8761,G11144);
  nand GNAME11168(G11168,G11167,G59558);
  and GNAME11169(G11169,G8768,G9866);
  or GNAME11170(G11170,G11169,G8753);
  nand GNAME11171(G11171,G8792,G8774);
  not GNAME11172(G11172,G8938);
  nand GNAME11173(G11173,G11105,G8941);
  nand GNAME11174(G11174,G11104,G13879);
  nand GNAME11175(G11175,G11103,G21670);
  nand GNAME11176(G11176,G11101,G21997);
  nand GNAME11177(G11177,G8828,G11172);
  nand GNAME11178(G11178,G8825,G9806);
  nand GNAME11179(G11179,G9403,G11175,G11173,G11176);
  nand GNAME11180(G11180,G21997,G8929);
  nand GNAME11181(G11181,G11179,G8790);
  nand GNAME11182(G11182,G11180,G11181);
  nand GNAME11183(G11183,G8792,G8962);
  nand GNAME11184(G11184,G59426,G8959);
  nand GNAME11185(G11185,G11183,G11184);
  not GNAME11186(G11186,G8947);
  nand GNAME11187(G11187,G8833,G8956);
  nand GNAME11188(G11188,G59426,G11186);
  nand GNAME11189(G11189,G11187,G11188);
  nand GNAME11190(G11190,G8947,G8948);
  and GNAME11191(G11191,G11190,G9800);
  nand GNAME11192(G11192,G8956,G8947,G8948);
  nand GNAME11193(G11193,G8957,G8958);
  nand GNAME11194(G11194,G11192,G11193);
  and GNAME11195(G11195,G8947,G59426);
  nor GNAME11196(G11196,G11195,G8802,G8958);
  or GNAME11197(G11197,G8957,G11196);
  nand GNAME11198(G11198,G11197,G8910);
  nand GNAME11199(G11199,G1652,G8949);
  nand GNAME11200(G11200,G11198,G59556);
  nand GNAME11201(G11201,G11194,G1659);
  nand GNAME11202(G11202,G11189,G8959);
  nand GNAME11203(G11203,G8960,G8961);
  nand GNAME11204(G11204,G11185,G8957);
  nand GNAME11205(G11205,G8796,G8962);
  nand GNAME11206(G11206,G59426,G8963);
  nand GNAME11207(G11207,G11205,G11206);
  nand GNAME11208(G11208,G1651,G8949);
  nand GNAME11209(G11209,G11198,G59555);
  nand GNAME11210(G11210,G11194,G1648);
  nand GNAME11211(G11211,G11189,G8963);
  nand GNAME11212(G11212,G8960,G8964);
  nand GNAME11213(G11213,G11207,G8957);
  nand GNAME11214(G11214,G8781,G8962);
  nand GNAME11215(G11215,G59426,G8965);
  nand GNAME11216(G11216,G11214,G11215);
  nand GNAME11217(G11217,G1650,G8949);
  nand GNAME11218(G11218,G11198,G59554);
  nand GNAME11219(G11219,G11194,G1637);
  nand GNAME11220(G11220,G11189,G8965);
  nand GNAME11221(G11221,G8960,G8966);
  nand GNAME11222(G11222,G11216,G8957);
  nand GNAME11223(G11223,G8746,G8962);
  nand GNAME11224(G11224,G59426,G8967);
  nand GNAME11225(G11225,G11223,G11224);
  nand GNAME11226(G11226,G1649,G8949);
  nand GNAME11227(G11227,G11198,G59553);
  nand GNAME11228(G11228,G11194,G1634);
  nand GNAME11229(G11229,G11189,G8967);
  nand GNAME11230(G11230,G8960,G8968);
  nand GNAME11231(G11231,G11225,G8957);
  nand GNAME11232(G11232,G8783,G8962);
  nand GNAME11233(G11233,G59426,G8969);
  nand GNAME11234(G11234,G11232,G11233);
  nand GNAME11235(G11235,G1647,G8949);
  nand GNAME11236(G11236,G11198,G59552);
  nand GNAME11237(G11237,G11194,G1633);
  nand GNAME11238(G11238,G11189,G8969);
  nand GNAME11239(G11239,G8960,G8970);
  nand GNAME11240(G11240,G11234,G8957);
  nand GNAME11241(G11241,G8780,G8962);
  nand GNAME11242(G11242,G59426,G8971);
  nand GNAME11243(G11243,G11241,G11242);
  nand GNAME11244(G11244,G1646,G8949);
  nand GNAME11245(G11245,G11198,G59551);
  nand GNAME11246(G11246,G11194,G1632);
  nand GNAME11247(G11247,G11189,G8971);
  nand GNAME11248(G11248,G8960,G8972);
  nand GNAME11249(G11249,G11243,G8957);
  nand GNAME11250(G11250,G8782,G8962);
  nand GNAME11251(G11251,G59426,G8973);
  nand GNAME11252(G11252,G11250,G11251);
  nand GNAME11253(G11253,G1645,G8949);
  nand GNAME11254(G11254,G11198,G59550);
  nand GNAME11255(G11255,G11194,G1631);
  nand GNAME11256(G11256,G11189,G8973);
  nand GNAME11257(G11257,G8960,G8974);
  nand GNAME11258(G11258,G11252,G8957);
  nand GNAME11259(G11259,G8852,G8962);
  nand GNAME11260(G11260,G59426,G8975);
  nand GNAME11261(G11261,G11259,G11260);
  nand GNAME11262(G11262,G1644,G8949);
  nand GNAME11263(G11263,G11198,G59549);
  nand GNAME11264(G11264,G11194,G1630);
  nand GNAME11265(G11265,G11189,G8975);
  nand GNAME11266(G11266,G8960,G8976);
  nand GNAME11267(G11267,G11261,G8957);
  not GNAME11268(G11268,G8979);
  nand GNAME11269(G11269,G8833,G8984);
  nand GNAME11270(G11270,G59426,G11268);
  nand GNAME11271(G11271,G11269,G11270);
  nand GNAME11272(G11272,G8979,G8980);
  and GNAME11273(G11273,G11272,G9800);
  nand GNAME11274(G11274,G8984,G8979,G8980);
  nand GNAME11275(G11275,G8985,G8986);
  nand GNAME11276(G11276,G11274,G11275);
  and GNAME11277(G11277,G8979,G59426);
  nor GNAME11278(G11278,G11277,G8802,G8986);
  or GNAME11279(G11279,G8985,G11278);
  nand GNAME11280(G11280,G11279,G8910);
  nand GNAME11281(G11281,G1652,G8981);
  nand GNAME11282(G11282,G11280,G59548);
  nand GNAME11283(G11283,G11276,G1659);
  nand GNAME11284(G11284,G11271,G8959);
  nand GNAME11285(G11285,G8961,G8987);
  nand GNAME11286(G11286,G11185,G8985);
  nand GNAME11287(G11287,G1651,G8981);
  nand GNAME11288(G11288,G11280,G59547);
  nand GNAME11289(G11289,G11276,G1648);
  nand GNAME11290(G11290,G11271,G8963);
  nand GNAME11291(G11291,G8964,G8987);
  nand GNAME11292(G11292,G11207,G8985);
  nand GNAME11293(G11293,G1650,G8981);
  nand GNAME11294(G11294,G11280,G59546);
  nand GNAME11295(G11295,G11276,G1637);
  nand GNAME11296(G11296,G11271,G8965);
  nand GNAME11297(G11297,G8966,G8987);
  nand GNAME11298(G11298,G11216,G8985);
  nand GNAME11299(G11299,G1649,G8981);
  nand GNAME11300(G11300,G11280,G59545);
  nand GNAME11301(G11301,G11276,G1634);
  nand GNAME11302(G11302,G11271,G8967);
  nand GNAME11303(G11303,G8968,G8987);
  nand GNAME11304(G11304,G11225,G8985);
  nand GNAME11305(G11305,G1647,G8981);
  nand GNAME11306(G11306,G11280,G59544);
  nand GNAME11307(G11307,G11276,G1633);
  nand GNAME11308(G11308,G11271,G8969);
  nand GNAME11309(G11309,G8970,G8987);
  nand GNAME11310(G11310,G11234,G8985);
  nand GNAME11311(G11311,G1646,G8981);
  nand GNAME11312(G11312,G11280,G59543);
  nand GNAME11313(G11313,G11276,G1632);
  nand GNAME11314(G11314,G11271,G8971);
  nand GNAME11315(G11315,G8972,G8987);
  nand GNAME11316(G11316,G11243,G8985);
  nand GNAME11317(G11317,G1645,G8981);
  nand GNAME11318(G11318,G11280,G59542);
  nand GNAME11319(G11319,G11276,G1631);
  nand GNAME11320(G11320,G11271,G8973);
  nand GNAME11321(G11321,G8974,G8987);
  nand GNAME11322(G11322,G11252,G8985);
  nand GNAME11323(G11323,G1644,G8981);
  nand GNAME11324(G11324,G11280,G59541);
  nand GNAME11325(G11325,G11276,G1630);
  nand GNAME11326(G11326,G11271,G8975);
  nand GNAME11327(G11327,G8976,G8987);
  nand GNAME11328(G11328,G11261,G8985);
  not GNAME11329(G11329,G8990);
  nand GNAME11330(G11330,G8833,G8995);
  nand GNAME11331(G11331,G59426,G11329);
  nand GNAME11332(G11332,G11330,G11331);
  nand GNAME11333(G11333,G8990,G8991);
  and GNAME11334(G11334,G11333,G9800);
  nand GNAME11335(G11335,G8995,G8990,G8991);
  nand GNAME11336(G11336,G8996,G8997);
  nand GNAME11337(G11337,G11335,G11336);
  and GNAME11338(G11338,G8990,G59426);
  nor GNAME11339(G11339,G11338,G8802,G8997);
  or GNAME11340(G11340,G8996,G11339);
  nand GNAME11341(G11341,G11340,G8910);
  nand GNAME11342(G11342,G1652,G8992);
  nand GNAME11343(G11343,G11341,G59540);
  nand GNAME11344(G11344,G11337,G1659);
  nand GNAME11345(G11345,G11332,G8959);
  nand GNAME11346(G11346,G8961,G8998);
  nand GNAME11347(G11347,G11185,G8996);
  nand GNAME11348(G11348,G1651,G8992);
  nand GNAME11349(G11349,G11341,G59539);
  nand GNAME11350(G11350,G11337,G1648);
  nand GNAME11351(G11351,G11332,G8963);
  nand GNAME11352(G11352,G8964,G8998);
  nand GNAME11353(G11353,G11207,G8996);
  nand GNAME11354(G11354,G1650,G8992);
  nand GNAME11355(G11355,G11341,G59538);
  nand GNAME11356(G11356,G11337,G1637);
  nand GNAME11357(G11357,G11332,G8965);
  nand GNAME11358(G11358,G8966,G8998);
  nand GNAME11359(G11359,G11216,G8996);
  nand GNAME11360(G11360,G1649,G8992);
  nand GNAME11361(G11361,G11341,G59537);
  nand GNAME11362(G11362,G11337,G1634);
  nand GNAME11363(G11363,G11332,G8967);
  nand GNAME11364(G11364,G8968,G8998);
  nand GNAME11365(G11365,G11225,G8996);
  nand GNAME11366(G11366,G1647,G8992);
  nand GNAME11367(G11367,G11341,G59536);
  nand GNAME11368(G11368,G11337,G1633);
  nand GNAME11369(G11369,G11332,G8969);
  nand GNAME11370(G11370,G8970,G8998);
  nand GNAME11371(G11371,G11234,G8996);
  nand GNAME11372(G11372,G1646,G8992);
  nand GNAME11373(G11373,G11341,G59535);
  nand GNAME11374(G11374,G11337,G1632);
  nand GNAME11375(G11375,G11332,G8971);
  nand GNAME11376(G11376,G8972,G8998);
  nand GNAME11377(G11377,G11243,G8996);
  nand GNAME11378(G11378,G1645,G8992);
  nand GNAME11379(G11379,G11341,G59534);
  nand GNAME11380(G11380,G11337,G1631);
  nand GNAME11381(G11381,G11332,G8973);
  nand GNAME11382(G11382,G8974,G8998);
  nand GNAME11383(G11383,G11252,G8996);
  nand GNAME11384(G11384,G1644,G8992);
  nand GNAME11385(G11385,G11341,G59533);
  nand GNAME11386(G11386,G11337,G1630);
  nand GNAME11387(G11387,G11332,G8975);
  nand GNAME11388(G11388,G8976,G8998);
  nand GNAME11389(G11389,G11261,G8996);
  not GNAME11390(G11390,G8999);
  nand GNAME11391(G11391,G8833,G9003);
  nand GNAME11392(G11392,G59426,G11390);
  nand GNAME11393(G11393,G11391,G11392);
  nand GNAME11394(G11394,G8999,G9000);
  and GNAME11395(G11395,G11394,G9800);
  nand GNAME11396(G11396,G9000,G9003);
  nand GNAME11397(G11397,G9004,G9005);
  nand GNAME11398(G11398,G11396,G11397);
  and GNAME11399(G11399,G8999,G59426);
  nor GNAME11400(G11400,G11399,G8802,G9005);
  or GNAME11401(G11401,G9004,G11400);
  nand GNAME11402(G11402,G11401,G8910);
  nand GNAME11403(G11403,G1652,G9001);
  nand GNAME11404(G11404,G11402,G59532);
  nand GNAME11405(G11405,G11398,G1659);
  nand GNAME11406(G11406,G11393,G8959);
  nand GNAME11407(G11407,G8961,G9006);
  nand GNAME11408(G11408,G11185,G9004);
  nand GNAME11409(G11409,G1651,G9001);
  nand GNAME11410(G11410,G11402,G59531);
  nand GNAME11411(G11411,G11398,G1648);
  nand GNAME11412(G11412,G11393,G8963);
  nand GNAME11413(G11413,G8964,G9006);
  nand GNAME11414(G11414,G11207,G9004);
  nand GNAME11415(G11415,G1650,G9001);
  nand GNAME11416(G11416,G11402,G59530);
  nand GNAME11417(G11417,G11398,G1637);
  nand GNAME11418(G11418,G11393,G8965);
  nand GNAME11419(G11419,G8966,G9006);
  nand GNAME11420(G11420,G11216,G9004);
  nand GNAME11421(G11421,G1649,G9001);
  nand GNAME11422(G11422,G11402,G59529);
  nand GNAME11423(G11423,G11398,G1634);
  nand GNAME11424(G11424,G11393,G8967);
  nand GNAME11425(G11425,G8968,G9006);
  nand GNAME11426(G11426,G11225,G9004);
  nand GNAME11427(G11427,G1647,G9001);
  nand GNAME11428(G11428,G11402,G59528);
  nand GNAME11429(G11429,G11398,G1633);
  nand GNAME11430(G11430,G11393,G8969);
  nand GNAME11431(G11431,G8970,G9006);
  nand GNAME11432(G11432,G11234,G9004);
  nand GNAME11433(G11433,G1646,G9001);
  nand GNAME11434(G11434,G11402,G59527);
  nand GNAME11435(G11435,G11398,G1632);
  nand GNAME11436(G11436,G11393,G8971);
  nand GNAME11437(G11437,G8972,G9006);
  nand GNAME11438(G11438,G11243,G9004);
  nand GNAME11439(G11439,G1645,G9001);
  nand GNAME11440(G11440,G11402,G59526);
  nand GNAME11441(G11441,G11398,G1631);
  nand GNAME11442(G11442,G11393,G8973);
  nand GNAME11443(G11443,G8974,G9006);
  nand GNAME11444(G11444,G11252,G9004);
  nand GNAME11445(G11445,G1644,G9001);
  nand GNAME11446(G11446,G11402,G59525);
  nand GNAME11447(G11447,G11398,G1630);
  nand GNAME11448(G11448,G11393,G8975);
  nand GNAME11449(G11449,G8976,G9006);
  nand GNAME11450(G11450,G11261,G9004);
  not GNAME11451(G11451,G9009);
  nand GNAME11452(G11452,G8833,G9013);
  nand GNAME11453(G11453,G59426,G11451);
  nand GNAME11454(G11454,G11452,G11453);
  nand GNAME11455(G11455,G9009,G9010);
  and GNAME11456(G11456,G11455,G9800);
  nand GNAME11457(G11457,G9013,G9009,G9010);
  nand GNAME11458(G11458,G9014,G9015);
  nand GNAME11459(G11459,G11457,G11458);
  and GNAME11460(G11460,G9009,G59426);
  nor GNAME11461(G11461,G11460,G8802,G9015);
  or GNAME11462(G11462,G9014,G11461);
  nand GNAME11463(G11463,G11462,G8910);
  nand GNAME11464(G11464,G1652,G9011);
  nand GNAME11465(G11465,G11463,G59524);
  nand GNAME11466(G11466,G11459,G1659);
  nand GNAME11467(G11467,G11454,G8959);
  nand GNAME11468(G11468,G8961,G9016);
  nand GNAME11469(G11469,G11185,G9014);
  nand GNAME11470(G11470,G1651,G9011);
  nand GNAME11471(G11471,G11463,G59523);
  nand GNAME11472(G11472,G11459,G1648);
  nand GNAME11473(G11473,G11454,G8963);
  nand GNAME11474(G11474,G8964,G9016);
  nand GNAME11475(G11475,G11207,G9014);
  nand GNAME11476(G11476,G1650,G9011);
  nand GNAME11477(G11477,G11463,G59522);
  nand GNAME11478(G11478,G11459,G1637);
  nand GNAME11479(G11479,G11454,G8965);
  nand GNAME11480(G11480,G8966,G9016);
  nand GNAME11481(G11481,G11216,G9014);
  nand GNAME11482(G11482,G1649,G9011);
  nand GNAME11483(G11483,G11463,G59521);
  nand GNAME11484(G11484,G11459,G1634);
  nand GNAME11485(G11485,G11454,G8967);
  nand GNAME11486(G11486,G8968,G9016);
  nand GNAME11487(G11487,G11225,G9014);
  nand GNAME11488(G11488,G1647,G9011);
  nand GNAME11489(G11489,G11463,G59520);
  nand GNAME11490(G11490,G11459,G1633);
  nand GNAME11491(G11491,G11454,G8969);
  nand GNAME11492(G11492,G8970,G9016);
  nand GNAME11493(G11493,G11234,G9014);
  nand GNAME11494(G11494,G1646,G9011);
  nand GNAME11495(G11495,G11463,G59519);
  nand GNAME11496(G11496,G11459,G1632);
  nand GNAME11497(G11497,G11454,G8971);
  nand GNAME11498(G11498,G8972,G9016);
  nand GNAME11499(G11499,G11243,G9014);
  nand GNAME11500(G11500,G1645,G9011);
  nand GNAME11501(G11501,G11463,G59518);
  nand GNAME11502(G11502,G11459,G1631);
  nand GNAME11503(G11503,G11454,G8973);
  nand GNAME11504(G11504,G8974,G9016);
  nand GNAME11505(G11505,G11252,G9014);
  nand GNAME11506(G11506,G1644,G9011);
  nand GNAME11507(G11507,G11463,G59517);
  nand GNAME11508(G11508,G11459,G1630);
  nand GNAME11509(G11509,G11454,G8975);
  nand GNAME11510(G11510,G8976,G9016);
  nand GNAME11511(G11511,G11261,G9014);
  not GNAME11512(G11512,G9019);
  nand GNAME11513(G11513,G8833,G9022);
  nand GNAME11514(G11514,G59426,G11512);
  nand GNAME11515(G11515,G11513,G11514);
  nand GNAME11516(G11516,G9019,G9020);
  and GNAME11517(G11517,G11516,G9800);
  nand GNAME11518(G11518,G9020,G9022);
  nand GNAME11519(G11519,G9023,G9024);
  nand GNAME11520(G11520,G11518,G11519);
  and GNAME11521(G11521,G9019,G59426);
  nor GNAME11522(G11522,G11521,G8802,G9024);
  or GNAME11523(G11523,G9023,G11522);
  nand GNAME11524(G11524,G11523,G8910);
  nand GNAME11525(G11525,G1652,G9021);
  nand GNAME11526(G11526,G11524,G59516);
  nand GNAME11527(G11527,G11520,G1659);
  nand GNAME11528(G11528,G11515,G8959);
  nand GNAME11529(G11529,G8961,G9025);
  nand GNAME11530(G11530,G11185,G9023);
  nand GNAME11531(G11531,G1651,G9021);
  nand GNAME11532(G11532,G11524,G59515);
  nand GNAME11533(G11533,G11520,G1648);
  nand GNAME11534(G11534,G11515,G8963);
  nand GNAME11535(G11535,G8964,G9025);
  nand GNAME11536(G11536,G11207,G9023);
  nand GNAME11537(G11537,G1650,G9021);
  nand GNAME11538(G11538,G11524,G59514);
  nand GNAME11539(G11539,G11520,G1637);
  nand GNAME11540(G11540,G11515,G8965);
  nand GNAME11541(G11541,G8966,G9025);
  nand GNAME11542(G11542,G11216,G9023);
  nand GNAME11543(G11543,G1649,G9021);
  nand GNAME11544(G11544,G11524,G59513);
  nand GNAME11545(G11545,G11520,G1634);
  nand GNAME11546(G11546,G11515,G8967);
  nand GNAME11547(G11547,G8968,G9025);
  nand GNAME11548(G11548,G11225,G9023);
  nand GNAME11549(G11549,G1647,G9021);
  nand GNAME11550(G11550,G11524,G59512);
  nand GNAME11551(G11551,G11520,G1633);
  nand GNAME11552(G11552,G11515,G8969);
  nand GNAME11553(G11553,G8970,G9025);
  nand GNAME11554(G11554,G11234,G9023);
  nand GNAME11555(G11555,G1646,G9021);
  nand GNAME11556(G11556,G11524,G59511);
  nand GNAME11557(G11557,G11520,G1632);
  nand GNAME11558(G11558,G11515,G8971);
  nand GNAME11559(G11559,G8972,G9025);
  nand GNAME11560(G11560,G11243,G9023);
  nand GNAME11561(G11561,G1645,G9021);
  nand GNAME11562(G11562,G11524,G59510);
  nand GNAME11563(G11563,G11520,G1631);
  nand GNAME11564(G11564,G11515,G8973);
  nand GNAME11565(G11565,G8974,G9025);
  nand GNAME11566(G11566,G11252,G9023);
  nand GNAME11567(G11567,G1644,G9021);
  nand GNAME11568(G11568,G11524,G59509);
  nand GNAME11569(G11569,G11520,G1630);
  nand GNAME11570(G11570,G11515,G8975);
  nand GNAME11571(G11571,G8976,G9025);
  nand GNAME11572(G11572,G11261,G9023);
  not GNAME11573(G11573,G9026);
  nand GNAME11574(G11574,G8833,G9029);
  nand GNAME11575(G11575,G59426,G11573);
  nand GNAME11576(G11576,G11574,G11575);
  nand GNAME11577(G11577,G9026,G9027);
  and GNAME11578(G11578,G11577,G9800);
  nand GNAME11579(G11579,G9029,G9026,G9027);
  nand GNAME11580(G11580,G9030,G9031);
  nand GNAME11581(G11581,G11579,G11580);
  and GNAME11582(G11582,G9026,G59426);
  nor GNAME11583(G11583,G11582,G8802,G9031);
  or GNAME11584(G11584,G9030,G11583);
  nand GNAME11585(G11585,G11584,G8910);
  nand GNAME11586(G11586,G1652,G9028);
  nand GNAME11587(G11587,G11585,G59508);
  nand GNAME11588(G11588,G11581,G1659);
  nand GNAME11589(G11589,G11576,G8959);
  nand GNAME11590(G11590,G8961,G9032);
  nand GNAME11591(G11591,G11185,G9030);
  nand GNAME11592(G11592,G1651,G9028);
  nand GNAME11593(G11593,G11585,G59507);
  nand GNAME11594(G11594,G11581,G1648);
  nand GNAME11595(G11595,G11576,G8963);
  nand GNAME11596(G11596,G8964,G9032);
  nand GNAME11597(G11597,G11207,G9030);
  nand GNAME11598(G11598,G1650,G9028);
  nand GNAME11599(G11599,G11585,G59506);
  nand GNAME11600(G11600,G11581,G1637);
  nand GNAME11601(G11601,G11576,G8965);
  nand GNAME11602(G11602,G8966,G9032);
  nand GNAME11603(G11603,G11216,G9030);
  nand GNAME11604(G11604,G1649,G9028);
  nand GNAME11605(G11605,G11585,G59505);
  nand GNAME11606(G11606,G11581,G1634);
  nand GNAME11607(G11607,G11576,G8967);
  nand GNAME11608(G11608,G8968,G9032);
  nand GNAME11609(G11609,G11225,G9030);
  nand GNAME11610(G11610,G1647,G9028);
  nand GNAME11611(G11611,G11585,G59504);
  nand GNAME11612(G11612,G11581,G1633);
  nand GNAME11613(G11613,G11576,G8969);
  nand GNAME11614(G11614,G8970,G9032);
  nand GNAME11615(G11615,G11234,G9030);
  nand GNAME11616(G11616,G1646,G9028);
  nand GNAME11617(G11617,G11585,G59503);
  nand GNAME11618(G11618,G11581,G1632);
  nand GNAME11619(G11619,G11576,G8971);
  nand GNAME11620(G11620,G8972,G9032);
  nand GNAME11621(G11621,G11243,G9030);
  nand GNAME11622(G11622,G1645,G9028);
  nand GNAME11623(G11623,G11585,G59502);
  nand GNAME11624(G11624,G11581,G1631);
  nand GNAME11625(G11625,G11576,G8973);
  nand GNAME11626(G11626,G8974,G9032);
  nand GNAME11627(G11627,G11252,G9030);
  nand GNAME11628(G11628,G1644,G9028);
  nand GNAME11629(G11629,G11585,G59501);
  nand GNAME11630(G11630,G11581,G1630);
  nand GNAME11631(G11631,G11576,G8975);
  nand GNAME11632(G11632,G8976,G9032);
  nand GNAME11633(G11633,G11261,G9030);
  not GNAME11634(G11634,G9033);
  nand GNAME11635(G11635,G8833,G9036);
  nand GNAME11636(G11636,G59426,G11634);
  nand GNAME11637(G11637,G11635,G11636);
  nand GNAME11638(G11638,G9033,G9034);
  and GNAME11639(G11639,G11638,G9800);
  nand GNAME11640(G11640,G9034,G9036);
  nand GNAME11641(G11641,G9037,G9038);
  nand GNAME11642(G11642,G11640,G11641);
  and GNAME11643(G11643,G9033,G59426);
  nor GNAME11644(G11644,G11643,G8802,G9037);
  or GNAME11645(G11645,G9038,G11644);
  nand GNAME11646(G11646,G11645,G8910);
  nand GNAME11647(G11647,G1652,G9035);
  nand GNAME11648(G11648,G11646,G59500);
  nand GNAME11649(G11649,G11642,G1659);
  nand GNAME11650(G11650,G11637,G8959);
  nand GNAME11651(G11651,G8961,G9039);
  nand GNAME11652(G11652,G11185,G9038);
  nand GNAME11653(G11653,G1651,G9035);
  nand GNAME11654(G11654,G11646,G59499);
  nand GNAME11655(G11655,G11642,G1648);
  nand GNAME11656(G11656,G11637,G8963);
  nand GNAME11657(G11657,G8964,G9039);
  nand GNAME11658(G11658,G11207,G9038);
  nand GNAME11659(G11659,G1650,G9035);
  nand GNAME11660(G11660,G11646,G59498);
  nand GNAME11661(G11661,G11642,G1637);
  nand GNAME11662(G11662,G11637,G8965);
  nand GNAME11663(G11663,G8966,G9039);
  nand GNAME11664(G11664,G11216,G9038);
  nand GNAME11665(G11665,G1649,G9035);
  nand GNAME11666(G11666,G11646,G59497);
  nand GNAME11667(G11667,G11642,G1634);
  nand GNAME11668(G11668,G11637,G8967);
  nand GNAME11669(G11669,G8968,G9039);
  nand GNAME11670(G11670,G11225,G9038);
  nand GNAME11671(G11671,G1647,G9035);
  nand GNAME11672(G11672,G11646,G59496);
  nand GNAME11673(G11673,G11642,G1633);
  nand GNAME11674(G11674,G11637,G8969);
  nand GNAME11675(G11675,G8970,G9039);
  nand GNAME11676(G11676,G11234,G9038);
  nand GNAME11677(G11677,G1646,G9035);
  nand GNAME11678(G11678,G11646,G59495);
  nand GNAME11679(G11679,G11642,G1632);
  nand GNAME11680(G11680,G11637,G8971);
  nand GNAME11681(G11681,G8972,G9039);
  nand GNAME11682(G11682,G11243,G9038);
  nand GNAME11683(G11683,G1645,G9035);
  nand GNAME11684(G11684,G11646,G59494);
  nand GNAME11685(G11685,G11642,G1631);
  nand GNAME11686(G11686,G11637,G8973);
  nand GNAME11687(G11687,G8974,G9039);
  nand GNAME11688(G11688,G11252,G9038);
  nand GNAME11689(G11689,G1644,G9035);
  nand GNAME11690(G11690,G11646,G59493);
  nand GNAME11691(G11691,G11642,G1630);
  nand GNAME11692(G11692,G11637,G8975);
  nand GNAME11693(G11693,G8976,G9039);
  nand GNAME11694(G11694,G11261,G9038);
  not GNAME11695(G11695,G9042);
  nand GNAME11696(G11696,G59426,G11695);
  nand GNAME11697(G11697,G8833,G9047);
  nand GNAME11698(G11698,G11696,G11697);
  nand GNAME11699(G11699,G9042,G9043);
  and GNAME11700(G11700,G11699,G9800);
  nand GNAME11701(G11701,G9047,G9042,G9043);
  nand GNAME11702(G11702,G9048,G9049);
  nand GNAME11703(G11703,G11701,G11702);
  and GNAME11704(G11704,G9042,G59426);
  nor GNAME11705(G11705,G11704,G8802,G9049);
  or GNAME11706(G11706,G9048,G11705);
  nand GNAME11707(G11707,G11706,G8910);
  nand GNAME11708(G11708,G1652,G9044);
  nand GNAME11709(G11709,G11707,G59492);
  nand GNAME11710(G11710,G11703,G1659);
  nand GNAME11711(G11711,G11698,G8959);
  nand GNAME11712(G11712,G8961,G9050);
  nand GNAME11713(G11713,G11185,G9048);
  nand GNAME11714(G11714,G1651,G9044);
  nand GNAME11715(G11715,G11707,G59491);
  nand GNAME11716(G11716,G11703,G1648);
  nand GNAME11717(G11717,G11698,G8963);
  nand GNAME11718(G11718,G8964,G9050);
  nand GNAME11719(G11719,G11207,G9048);
  nand GNAME11720(G11720,G1650,G9044);
  nand GNAME11721(G11721,G11707,G59490);
  nand GNAME11722(G11722,G11703,G1637);
  nand GNAME11723(G11723,G11698,G8965);
  nand GNAME11724(G11724,G8966,G9050);
  nand GNAME11725(G11725,G11216,G9048);
  nand GNAME11726(G11726,G1649,G9044);
  nand GNAME11727(G11727,G11707,G59489);
  nand GNAME11728(G11728,G11703,G1634);
  nand GNAME11729(G11729,G11698,G8967);
  nand GNAME11730(G11730,G8968,G9050);
  nand GNAME11731(G11731,G11225,G9048);
  nand GNAME11732(G11732,G1647,G9044);
  nand GNAME11733(G11733,G11707,G59488);
  nand GNAME11734(G11734,G11703,G1633);
  nand GNAME11735(G11735,G11698,G8969);
  nand GNAME11736(G11736,G8970,G9050);
  nand GNAME11737(G11737,G11234,G9048);
  nand GNAME11738(G11738,G1646,G9044);
  nand GNAME11739(G11739,G11707,G59487);
  nand GNAME11740(G11740,G11703,G1632);
  nand GNAME11741(G11741,G11698,G8971);
  nand GNAME11742(G11742,G8972,G9050);
  nand GNAME11743(G11743,G11243,G9048);
  nand GNAME11744(G11744,G1645,G9044);
  nand GNAME11745(G11745,G11707,G59486);
  nand GNAME11746(G11746,G11703,G1631);
  nand GNAME11747(G11747,G11698,G8973);
  nand GNAME11748(G11748,G8974,G9050);
  nand GNAME11749(G11749,G11252,G9048);
  nand GNAME11750(G11750,G1644,G9044);
  nand GNAME11751(G11751,G11707,G59485);
  nand GNAME11752(G11752,G11703,G1630);
  nand GNAME11753(G11753,G11698,G8975);
  nand GNAME11754(G11754,G8976,G9050);
  nand GNAME11755(G11755,G11261,G9048);
  not GNAME11756(G11756,G9051);
  nand GNAME11757(G11757,G59426,G11756);
  nand GNAME11758(G11758,G8833,G9054);
  nand GNAME11759(G11759,G11757,G11758);
  nand GNAME11760(G11760,G9051,G9052);
  and GNAME11761(G11761,G11760,G9800);
  nand GNAME11762(G11762,G9054,G9051,G9052);
  nand GNAME11763(G11763,G9055,G9056);
  nand GNAME11764(G11764,G11762,G11763);
  and GNAME11765(G11765,G9051,G59426);
  nor GNAME11766(G11766,G11765,G8802,G9056);
  or GNAME11767(G11767,G9055,G11766);
  nand GNAME11768(G11768,G11767,G8910);
  nand GNAME11769(G11769,G1652,G9053);
  nand GNAME11770(G11770,G11768,G59484);
  nand GNAME11771(G11771,G11764,G1659);
  nand GNAME11772(G11772,G11759,G8959);
  nand GNAME11773(G11773,G8961,G9057);
  nand GNAME11774(G11774,G11185,G9055);
  nand GNAME11775(G11775,G1651,G9053);
  nand GNAME11776(G11776,G11768,G59483);
  nand GNAME11777(G11777,G11764,G1648);
  nand GNAME11778(G11778,G11759,G8963);
  nand GNAME11779(G11779,G8964,G9057);
  nand GNAME11780(G11780,G11207,G9055);
  nand GNAME11781(G11781,G1650,G9053);
  nand GNAME11782(G11782,G11768,G59482);
  nand GNAME11783(G11783,G11764,G1637);
  nand GNAME11784(G11784,G11759,G8965);
  nand GNAME11785(G11785,G8966,G9057);
  nand GNAME11786(G11786,G11216,G9055);
  nand GNAME11787(G11787,G1649,G9053);
  nand GNAME11788(G11788,G11768,G59481);
  nand GNAME11789(G11789,G11764,G1634);
  nand GNAME11790(G11790,G11759,G8967);
  nand GNAME11791(G11791,G8968,G9057);
  nand GNAME11792(G11792,G11225,G9055);
  nand GNAME11793(G11793,G1647,G9053);
  nand GNAME11794(G11794,G11768,G59480);
  nand GNAME11795(G11795,G11764,G1633);
  nand GNAME11796(G11796,G11759,G8969);
  nand GNAME11797(G11797,G8970,G9057);
  nand GNAME11798(G11798,G11234,G9055);
  nand GNAME11799(G11799,G1646,G9053);
  nand GNAME11800(G11800,G11768,G59479);
  nand GNAME11801(G11801,G11764,G1632);
  nand GNAME11802(G11802,G11759,G8971);
  nand GNAME11803(G11803,G8972,G9057);
  nand GNAME11804(G11804,G11243,G9055);
  nand GNAME11805(G11805,G1645,G9053);
  nand GNAME11806(G11806,G11768,G59478);
  nand GNAME11807(G11807,G11764,G1631);
  nand GNAME11808(G11808,G11759,G8973);
  nand GNAME11809(G11809,G8974,G9057);
  nand GNAME11810(G11810,G11252,G9055);
  nand GNAME11811(G11811,G1644,G9053);
  nand GNAME11812(G11812,G11768,G59477);
  nand GNAME11813(G11813,G11764,G1630);
  nand GNAME11814(G11814,G11759,G8975);
  nand GNAME11815(G11815,G8976,G9057);
  nand GNAME11816(G11816,G11261,G9055);
  not GNAME11817(G11817,G9060);
  nand GNAME11818(G11818,G59426,G11817);
  nand GNAME11819(G11819,G8833,G9063);
  nand GNAME11820(G11820,G11818,G11819);
  nand GNAME11821(G11821,G9060,G9061);
  and GNAME11822(G11822,G11821,G9800);
  nand GNAME11823(G11823,G9063,G9060,G9061);
  nand GNAME11824(G11824,G9064,G9065);
  nand GNAME11825(G11825,G11823,G11824);
  and GNAME11826(G11826,G9060,G59426);
  nor GNAME11827(G11827,G11826,G8802,G9065);
  or GNAME11828(G11828,G9064,G11827);
  nand GNAME11829(G11829,G11828,G8910);
  nand GNAME11830(G11830,G1652,G9062);
  nand GNAME11831(G11831,G11829,G59476);
  nand GNAME11832(G11832,G11825,G1659);
  nand GNAME11833(G11833,G11820,G8959);
  nand GNAME11834(G11834,G8961,G9066);
  nand GNAME11835(G11835,G11185,G9064);
  nand GNAME11836(G11836,G1651,G9062);
  nand GNAME11837(G11837,G11829,G59475);
  nand GNAME11838(G11838,G11825,G1648);
  nand GNAME11839(G11839,G11820,G8963);
  nand GNAME11840(G11840,G8964,G9066);
  nand GNAME11841(G11841,G11207,G9064);
  nand GNAME11842(G11842,G1650,G9062);
  nand GNAME11843(G11843,G11829,G59474);
  nand GNAME11844(G11844,G11825,G1637);
  nand GNAME11845(G11845,G11820,G8965);
  nand GNAME11846(G11846,G8966,G9066);
  nand GNAME11847(G11847,G11216,G9064);
  nand GNAME11848(G11848,G1649,G9062);
  nand GNAME11849(G11849,G11829,G59473);
  nand GNAME11850(G11850,G11825,G1634);
  nand GNAME11851(G11851,G11820,G8967);
  nand GNAME11852(G11852,G8968,G9066);
  nand GNAME11853(G11853,G11225,G9064);
  nand GNAME11854(G11854,G1647,G9062);
  nand GNAME11855(G11855,G11829,G59472);
  nand GNAME11856(G11856,G11825,G1633);
  nand GNAME11857(G11857,G11820,G8969);
  nand GNAME11858(G11858,G8970,G9066);
  nand GNAME11859(G11859,G11234,G9064);
  nand GNAME11860(G11860,G1646,G9062);
  nand GNAME11861(G11861,G11829,G59471);
  nand GNAME11862(G11862,G11825,G1632);
  nand GNAME11863(G11863,G11820,G8971);
  nand GNAME11864(G11864,G8972,G9066);
  nand GNAME11865(G11865,G11243,G9064);
  nand GNAME11866(G11866,G1645,G9062);
  nand GNAME11867(G11867,G11829,G59470);
  nand GNAME11868(G11868,G11825,G1631);
  nand GNAME11869(G11869,G11820,G8973);
  nand GNAME11870(G11870,G8974,G9066);
  nand GNAME11871(G11871,G11252,G9064);
  nand GNAME11872(G11872,G1644,G9062);
  nand GNAME11873(G11873,G11829,G59469);
  nand GNAME11874(G11874,G11825,G1630);
  nand GNAME11875(G11875,G11820,G8975);
  nand GNAME11876(G11876,G8976,G9066);
  nand GNAME11877(G11877,G11261,G9064);
  not GNAME11878(G11878,G9067);
  nand GNAME11879(G11879,G59426,G11878);
  nand GNAME11880(G11880,G8833,G9070);
  nand GNAME11881(G11881,G11879,G11880);
  nand GNAME11882(G11882,G9067,G9068);
  and GNAME11883(G11883,G11882,G9800);
  nand GNAME11884(G11884,G9068,G9070);
  nand GNAME11885(G11885,G9071,G9072);
  nand GNAME11886(G11886,G11884,G11885);
  and GNAME11887(G11887,G9067,G59426);
  nor GNAME11888(G11888,G11887,G8802,G9072);
  or GNAME11889(G11889,G9071,G11888);
  nand GNAME11890(G11890,G11889,G8910);
  nand GNAME11891(G11891,G1652,G9069);
  nand GNAME11892(G11892,G11890,G59468);
  nand GNAME11893(G11893,G11886,G1659);
  nand GNAME11894(G11894,G11881,G8959);
  nand GNAME11895(G11895,G8961,G9073);
  nand GNAME11896(G11896,G11185,G9071);
  nand GNAME11897(G11897,G1651,G9069);
  nand GNAME11898(G11898,G11890,G59467);
  nand GNAME11899(G11899,G11886,G1648);
  nand GNAME11900(G11900,G11881,G8963);
  nand GNAME11901(G11901,G8964,G9073);
  nand GNAME11902(G11902,G11207,G9071);
  nand GNAME11903(G11903,G1650,G9069);
  nand GNAME11904(G11904,G11890,G59466);
  nand GNAME11905(G11905,G11886,G1637);
  nand GNAME11906(G11906,G11881,G8965);
  nand GNAME11907(G11907,G8966,G9073);
  nand GNAME11908(G11908,G11216,G9071);
  nand GNAME11909(G11909,G1649,G9069);
  nand GNAME11910(G11910,G11890,G59465);
  nand GNAME11911(G11911,G11886,G1634);
  nand GNAME11912(G11912,G11881,G8967);
  nand GNAME11913(G11913,G8968,G9073);
  nand GNAME11914(G11914,G11225,G9071);
  nand GNAME11915(G11915,G1647,G9069);
  nand GNAME11916(G11916,G11890,G59464);
  nand GNAME11917(G11917,G11886,G1633);
  nand GNAME11918(G11918,G11881,G8969);
  nand GNAME11919(G11919,G8970,G9073);
  nand GNAME11920(G11920,G11234,G9071);
  nand GNAME11921(G11921,G1646,G9069);
  nand GNAME11922(G11922,G11890,G59463);
  nand GNAME11923(G11923,G11886,G1632);
  nand GNAME11924(G11924,G11881,G8971);
  nand GNAME11925(G11925,G8972,G9073);
  nand GNAME11926(G11926,G11243,G9071);
  nand GNAME11927(G11927,G1645,G9069);
  nand GNAME11928(G11928,G11890,G59462);
  nand GNAME11929(G11929,G11886,G1631);
  nand GNAME11930(G11930,G11881,G8973);
  nand GNAME11931(G11931,G8974,G9073);
  nand GNAME11932(G11932,G11252,G9071);
  nand GNAME11933(G11933,G1644,G9069);
  nand GNAME11934(G11934,G11890,G59461);
  nand GNAME11935(G11935,G11886,G1630);
  nand GNAME11936(G11936,G11881,G8975);
  nand GNAME11937(G11937,G8976,G9073);
  nand GNAME11938(G11938,G11261,G9071);
  not GNAME11939(G11939,G9074);
  nand GNAME11940(G11940,G59426,G11939);
  nand GNAME11941(G11941,G8833,G9079);
  nand GNAME11942(G11942,G11940,G11941);
  nand GNAME11943(G11943,G9074,G9075);
  and GNAME11944(G11944,G11943,G9800);
  nand GNAME11945(G11945,G9079,G9074,G9075);
  nand GNAME11946(G11946,G9080,G9081);
  nand GNAME11947(G11947,G11945,G11946);
  and GNAME11948(G11948,G9074,G59426);
  nor GNAME11949(G11949,G11948,G8802,G9081);
  or GNAME11950(G11950,G9080,G11949);
  nand GNAME11951(G11951,G11950,G8910);
  nand GNAME11952(G11952,G1652,G9076);
  nand GNAME11953(G11953,G11951,G59460);
  nand GNAME11954(G11954,G11947,G1659);
  nand GNAME11955(G11955,G11942,G8959);
  nand GNAME11956(G11956,G8961,G9082);
  nand GNAME11957(G11957,G11185,G9080);
  nand GNAME11958(G11958,G1651,G9076);
  nand GNAME11959(G11959,G11951,G59459);
  nand GNAME11960(G11960,G11947,G1648);
  nand GNAME11961(G11961,G11942,G8963);
  nand GNAME11962(G11962,G8964,G9082);
  nand GNAME11963(G11963,G11207,G9080);
  nand GNAME11964(G11964,G1650,G9076);
  nand GNAME11965(G11965,G11951,G59458);
  nand GNAME11966(G11966,G11947,G1637);
  nand GNAME11967(G11967,G11942,G8965);
  nand GNAME11968(G11968,G8966,G9082);
  nand GNAME11969(G11969,G11216,G9080);
  nand GNAME11970(G11970,G1649,G9076);
  nand GNAME11971(G11971,G11951,G59457);
  nand GNAME11972(G11972,G11947,G1634);
  nand GNAME11973(G11973,G11942,G8967);
  nand GNAME11974(G11974,G8968,G9082);
  nand GNAME11975(G11975,G11225,G9080);
  nand GNAME11976(G11976,G1647,G9076);
  nand GNAME11977(G11977,G11951,G59456);
  nand GNAME11978(G11978,G11947,G1633);
  nand GNAME11979(G11979,G11942,G8969);
  nand GNAME11980(G11980,G8970,G9082);
  nand GNAME11981(G11981,G11234,G9080);
  nand GNAME11982(G11982,G1646,G9076);
  nand GNAME11983(G11983,G11951,G59455);
  nand GNAME11984(G11984,G11947,G1632);
  nand GNAME11985(G11985,G11942,G8971);
  nand GNAME11986(G11986,G8972,G9082);
  nand GNAME11987(G11987,G11243,G9080);
  nand GNAME11988(G11988,G1645,G9076);
  nand GNAME11989(G11989,G11951,G59454);
  nand GNAME11990(G11990,G11947,G1631);
  nand GNAME11991(G11991,G11942,G8973);
  nand GNAME11992(G11992,G8974,G9082);
  nand GNAME11993(G11993,G11252,G9080);
  nand GNAME11994(G11994,G1644,G9076);
  nand GNAME11995(G11995,G11951,G59453);
  nand GNAME11996(G11996,G11947,G1630);
  nand GNAME11997(G11997,G11942,G8975);
  nand GNAME11998(G11998,G8976,G9082);
  nand GNAME11999(G11999,G11261,G9080);
  not GNAME12000(G12000,G9083);
  nand GNAME12001(G12001,G59426,G12000);
  nand GNAME12002(G12002,G8833,G9086);
  nand GNAME12003(G12003,G12001,G12002);
  nand GNAME12004(G12004,G9083,G9084);
  and GNAME12005(G12005,G12004,G9800);
  nand GNAME12006(G12006,G9086,G9083,G9084);
  nand GNAME12007(G12007,G9087,G9088);
  nand GNAME12008(G12008,G12006,G12007);
  and GNAME12009(G12009,G9083,G59426);
  nor GNAME12010(G12010,G12009,G8802,G9088);
  or GNAME12011(G12011,G9087,G12010);
  nand GNAME12012(G12012,G12011,G8910);
  nand GNAME12013(G12013,G1652,G9085);
  nand GNAME12014(G12014,G12012,G59452);
  nand GNAME12015(G12015,G12008,G1659);
  nand GNAME12016(G12016,G12003,G8959);
  nand GNAME12017(G12017,G8961,G9089);
  nand GNAME12018(G12018,G11185,G9087);
  nand GNAME12019(G12019,G1651,G9085);
  nand GNAME12020(G12020,G12012,G59451);
  nand GNAME12021(G12021,G12008,G1648);
  nand GNAME12022(G12022,G12003,G8963);
  nand GNAME12023(G12023,G8964,G9089);
  nand GNAME12024(G12024,G11207,G9087);
  nand GNAME12025(G12025,G1650,G9085);
  nand GNAME12026(G12026,G12012,G59450);
  nand GNAME12027(G12027,G12008,G1637);
  nand GNAME12028(G12028,G12003,G8965);
  nand GNAME12029(G12029,G8966,G9089);
  nand GNAME12030(G12030,G11216,G9087);
  nand GNAME12031(G12031,G1649,G9085);
  nand GNAME12032(G12032,G12012,G59449);
  nand GNAME12033(G12033,G12008,G1634);
  nand GNAME12034(G12034,G12003,G8967);
  nand GNAME12035(G12035,G8968,G9089);
  nand GNAME12036(G12036,G11225,G9087);
  nand GNAME12037(G12037,G1647,G9085);
  nand GNAME12038(G12038,G12012,G59448);
  nand GNAME12039(G12039,G12008,G1633);
  nand GNAME12040(G12040,G12003,G8969);
  nand GNAME12041(G12041,G8970,G9089);
  nand GNAME12042(G12042,G11234,G9087);
  nand GNAME12043(G12043,G1646,G9085);
  nand GNAME12044(G12044,G12012,G59447);
  nand GNAME12045(G12045,G12008,G1632);
  nand GNAME12046(G12046,G12003,G8971);
  nand GNAME12047(G12047,G8972,G9089);
  nand GNAME12048(G12048,G11243,G9087);
  nand GNAME12049(G12049,G1645,G9085);
  nand GNAME12050(G12050,G12012,G59446);
  nand GNAME12051(G12051,G12008,G1631);
  nand GNAME12052(G12052,G12003,G8973);
  nand GNAME12053(G12053,G8974,G9089);
  nand GNAME12054(G12054,G11252,G9087);
  nand GNAME12055(G12055,G1644,G9085);
  nand GNAME12056(G12056,G12012,G59445);
  nand GNAME12057(G12057,G12008,G1630);
  nand GNAME12058(G12058,G12003,G8975);
  nand GNAME12059(G12059,G8976,G9089);
  nand GNAME12060(G12060,G11261,G9087);
  not GNAME12061(G12061,G9090);
  nand GNAME12062(G12062,G59426,G12061);
  nand GNAME12063(G12063,G8833,G9093);
  nand GNAME12064(G12064,G12062,G12063);
  nand GNAME12065(G12065,G9090,G9091);
  and GNAME12066(G12066,G12065,G9800);
  nand GNAME12067(G12067,G9093,G9090,G9091);
  nand GNAME12068(G12068,G9094,G9095);
  nand GNAME12069(G12069,G12067,G12068);
  and GNAME12070(G12070,G9090,G59426);
  nor GNAME12071(G12071,G12070,G8802,G9095);
  or GNAME12072(G12072,G9094,G12071);
  nand GNAME12073(G12073,G12072,G8910);
  nand GNAME12074(G12074,G1652,G9092);
  nand GNAME12075(G12075,G12073,G59444);
  nand GNAME12076(G12076,G12069,G1659);
  nand GNAME12077(G12077,G12064,G8959);
  nand GNAME12078(G12078,G8961,G9096);
  nand GNAME12079(G12079,G11185,G9094);
  nand GNAME12080(G12080,G1651,G9092);
  nand GNAME12081(G12081,G12073,G59443);
  nand GNAME12082(G12082,G12069,G1648);
  nand GNAME12083(G12083,G12064,G8963);
  nand GNAME12084(G12084,G8964,G9096);
  nand GNAME12085(G12085,G11207,G9094);
  nand GNAME12086(G12086,G1650,G9092);
  nand GNAME12087(G12087,G12073,G59442);
  nand GNAME12088(G12088,G12069,G1637);
  nand GNAME12089(G12089,G12064,G8965);
  nand GNAME12090(G12090,G8966,G9096);
  nand GNAME12091(G12091,G11216,G9094);
  nand GNAME12092(G12092,G1649,G9092);
  nand GNAME12093(G12093,G12073,G59441);
  nand GNAME12094(G12094,G12069,G1634);
  nand GNAME12095(G12095,G12064,G8967);
  nand GNAME12096(G12096,G8968,G9096);
  nand GNAME12097(G12097,G11225,G9094);
  nand GNAME12098(G12098,G1647,G9092);
  nand GNAME12099(G12099,G12073,G59440);
  nand GNAME12100(G12100,G12069,G1633);
  nand GNAME12101(G12101,G12064,G8969);
  nand GNAME12102(G12102,G8970,G9096);
  nand GNAME12103(G12103,G11234,G9094);
  nand GNAME12104(G12104,G1646,G9092);
  nand GNAME12105(G12105,G12073,G59439);
  nand GNAME12106(G12106,G12069,G1632);
  nand GNAME12107(G12107,G12064,G8971);
  nand GNAME12108(G12108,G8972,G9096);
  nand GNAME12109(G12109,G11243,G9094);
  nand GNAME12110(G12110,G1645,G9092);
  nand GNAME12111(G12111,G12073,G59438);
  nand GNAME12112(G12112,G12069,G1631);
  nand GNAME12113(G12113,G12064,G8973);
  nand GNAME12114(G12114,G8974,G9096);
  nand GNAME12115(G12115,G11252,G9094);
  nand GNAME12116(G12116,G1644,G9092);
  nand GNAME12117(G12117,G12073,G59437);
  nand GNAME12118(G12118,G12069,G1630);
  nand GNAME12119(G12119,G12064,G8975);
  nand GNAME12120(G12120,G8976,G9096);
  nand GNAME12121(G12121,G11261,G9094);
  not GNAME12122(G12122,G9097);
  nand GNAME12123(G12123,G59426,G12122);
  nand GNAME12124(G12124,G8833,G9100);
  nand GNAME12125(G12125,G12123,G12124);
  nand GNAME12126(G12126,G9097,G9098);
  and GNAME12127(G12127,G12126,G9800);
  nand GNAME12128(G12128,G9098,G9100);
  nand GNAME12129(G12129,G9101,G9102);
  nand GNAME12130(G12130,G12128,G12129);
  and GNAME12131(G12131,G9097,G59426);
  nor GNAME12132(G12132,G12131,G8802,G9101);
  or GNAME12133(G12133,G9102,G12132);
  nand GNAME12134(G12134,G12133,G8910);
  nand GNAME12135(G12135,G1652,G9099);
  nand GNAME12136(G12136,G12134,G59436);
  nand GNAME12137(G12137,G12130,G1659);
  nand GNAME12138(G12138,G12125,G8959);
  nand GNAME12139(G12139,G11185,G9102);
  nand GNAME12140(G12140,G8961,G9103);
  nand GNAME12141(G12141,G1651,G9099);
  nand GNAME12142(G12142,G12134,G59435);
  nand GNAME12143(G12143,G12130,G1648);
  nand GNAME12144(G12144,G12125,G8963);
  nand GNAME12145(G12145,G11207,G9102);
  nand GNAME12146(G12146,G8964,G9103);
  nand GNAME12147(G12147,G1650,G9099);
  nand GNAME12148(G12148,G12134,G59434);
  nand GNAME12149(G12149,G12130,G1637);
  nand GNAME12150(G12150,G12125,G8965);
  nand GNAME12151(G12151,G11216,G9102);
  nand GNAME12152(G12152,G8966,G9103);
  nand GNAME12153(G12153,G1649,G9099);
  nand GNAME12154(G12154,G12134,G59433);
  nand GNAME12155(G12155,G12130,G1634);
  nand GNAME12156(G12156,G12125,G8967);
  nand GNAME12157(G12157,G11225,G9102);
  nand GNAME12158(G12158,G8968,G9103);
  nand GNAME12159(G12159,G1647,G9099);
  nand GNAME12160(G12160,G12134,G59432);
  nand GNAME12161(G12161,G12130,G1633);
  nand GNAME12162(G12162,G12125,G8969);
  nand GNAME12163(G12163,G11234,G9102);
  nand GNAME12164(G12164,G8970,G9103);
  nand GNAME12165(G12165,G1646,G9099);
  nand GNAME12166(G12166,G12134,G59431);
  nand GNAME12167(G12167,G12130,G1632);
  nand GNAME12168(G12168,G12125,G8971);
  nand GNAME12169(G12169,G11243,G9102);
  nand GNAME12170(G12170,G8972,G9103);
  nand GNAME12171(G12171,G1645,G9099);
  nand GNAME12172(G12172,G12134,G59430);
  nand GNAME12173(G12173,G12130,G1631);
  nand GNAME12174(G12174,G12125,G8973);
  nand GNAME12175(G12175,G11252,G9102);
  nand GNAME12176(G12176,G8974,G9103);
  nand GNAME12177(G12177,G1644,G9099);
  nand GNAME12178(G12178,G12134,G59429);
  nand GNAME12179(G12179,G12130,G1630);
  nand GNAME12180(G12180,G12125,G8975);
  nand GNAME12181(G12181,G11261,G9102);
  nand GNAME12182(G12182,G8976,G9103);
  nand GNAME12183(G12183,G9105,G8794,G8799);
  or GNAME12184(G12184,G59795,G59796);
  nand GNAME12185(G12185,G8801,G12183);
  nand GNAME12186(G12186,G8789,G8786);
  nand GNAME12187(G12187,G8814,G9106);
  nand GNAME12188(G12188,G1588,G59427);
  nand GNAME12189(G12189,G8835,G9955,G9977);
  nand GNAME12190(G12190,G59425,G21598,G8802);
  nand GNAME12191(G12191,G8787,G12190);
  or GNAME12192(G12192,G9106,G9798);
  nand GNAME12193(G12193,G21598,G8907);
  nand GNAME12194(G12194,G12193,G12191,G12192);
  nand GNAME12195(G12195,G9108,G8749,G59428);
  nand GNAME12196(G12196,G12195,G9804);
  nand GNAME12197(G12197,G9810,G9107);
  nand GNAME12198(G12198,G12197,G59427);
  nand GNAME12199(G12199,G9107,G12196);
  nand GNAME12200(G12200,G8839,G8749,G59427);
  nand GNAME12201(G12201,G8787,G8940);
  or GNAME12202(G12202,G8834,G9107);
  or GNAME12203(G12203,G59390,G59392);
  nand GNAME12204(G12204,G12203,G9771);
  nand GNAME12205(G12205,G8748,G59798);
  nand GNAME12206(G12206,G8806,G34);
  nand GNAME12207(G12207,G59798,G9110,G12206);
  or GNAME12208(G12208,G8749,G8805);
  nand GNAME12209(G12209,G8749,G59390);
  or GNAME12210(G12210,G1588,G33);
  nand GNAME12211(G12211,G8812,G59390);
  nand GNAME12212(G12212,G8748,G12205);
  nand GNAME12213(G12213,G59392,G9109,G12212);
  nand GNAME12214(G12214,G12213,G8817);
  or GNAME12215(G12215,G9110,G8812,G8748);
  nand GNAME12216(G12216,G9784,G59389);
  nand GNAME12217(G12217,G59760,G9111);
  nand GNAME12218(G12218,G59759,G9112);
  nand GNAME12219(G12219,G9784,G59388);
  nand GNAME12220(G12220,G59760,G9112);
  nand GNAME12221(G12221,G59761,G9111);
  nand GNAME12222(G12222,G9784,G59387);
  nand GNAME12223(G12223,G59761,G9112);
  nand GNAME12224(G12224,G59762,G9111);
  nand GNAME12225(G12225,G9784,G59386);
  nand GNAME12226(G12226,G59762,G9112);
  nand GNAME12227(G12227,G59763,G9111);
  nand GNAME12228(G12228,G9784,G59385);
  nand GNAME12229(G12229,G59763,G9112);
  nand GNAME12230(G12230,G59764,G9111);
  nand GNAME12231(G12231,G9784,G59384);
  nand GNAME12232(G12232,G59764,G9112);
  nand GNAME12233(G12233,G59765,G9111);
  nand GNAME12234(G12234,G9784,G59383);
  nand GNAME12235(G12235,G59765,G9112);
  nand GNAME12236(G12236,G59766,G9111);
  nand GNAME12237(G12237,G9784,G59382);
  nand GNAME12238(G12238,G59766,G9112);
  nand GNAME12239(G12239,G59767,G9111);
  nand GNAME12240(G12240,G9784,G59381);
  nand GNAME12241(G12241,G59767,G9112);
  nand GNAME12242(G12242,G59768,G9111);
  nand GNAME12243(G12243,G9784,G59380);
  nand GNAME12244(G12244,G59768,G9112);
  nand GNAME12245(G12245,G59769,G9111);
  nand GNAME12246(G12246,G9784,G59379);
  nand GNAME12247(G12247,G59769,G9112);
  nand GNAME12248(G12248,G59770,G9111);
  nand GNAME12249(G12249,G9784,G59378);
  nand GNAME12250(G12250,G59770,G9112);
  nand GNAME12251(G12251,G59771,G9111);
  nand GNAME12252(G12252,G9784,G59377);
  nand GNAME12253(G12253,G59771,G9112);
  nand GNAME12254(G12254,G59772,G9111);
  nand GNAME12255(G12255,G9784,G59376);
  nand GNAME12256(G12256,G59772,G9112);
  nand GNAME12257(G12257,G59773,G9111);
  nand GNAME12258(G12258,G9784,G59375);
  nand GNAME12259(G12259,G59773,G9112);
  nand GNAME12260(G12260,G59774,G9111);
  nand GNAME12261(G12261,G9784,G59374);
  nand GNAME12262(G12262,G59774,G9112);
  nand GNAME12263(G12263,G59775,G9111);
  nand GNAME12264(G12264,G9784,G59373);
  nand GNAME12265(G12265,G59775,G9112);
  nand GNAME12266(G12266,G59776,G9111);
  nand GNAME12267(G12267,G9784,G59372);
  nand GNAME12268(G12268,G59776,G9112);
  nand GNAME12269(G12269,G59777,G9111);
  nand GNAME12270(G12270,G9784,G59371);
  nand GNAME12271(G12271,G59777,G9112);
  nand GNAME12272(G12272,G59778,G9111);
  nand GNAME12273(G12273,G9784,G59370);
  nand GNAME12274(G12274,G59778,G9112);
  nand GNAME12275(G12275,G59779,G9111);
  nand GNAME12276(G12276,G9784,G59369);
  nand GNAME12277(G12277,G59779,G9112);
  nand GNAME12278(G12278,G59780,G9111);
  nand GNAME12279(G12279,G9784,G59368);
  nand GNAME12280(G12280,G59780,G9112);
  nand GNAME12281(G12281,G59781,G9111);
  nand GNAME12282(G12282,G9784,G59367);
  nand GNAME12283(G12283,G59781,G9112);
  nand GNAME12284(G12284,G59782,G9111);
  nand GNAME12285(G12285,G9784,G59366);
  nand GNAME12286(G12286,G59782,G9112);
  nand GNAME12287(G12287,G59783,G9111);
  nand GNAME12288(G12288,G9784,G59365);
  nand GNAME12289(G12289,G59783,G9112);
  nand GNAME12290(G12290,G59784,G9111);
  nand GNAME12291(G12291,G9784,G59364);
  nand GNAME12292(G12292,G59784,G9112);
  nand GNAME12293(G12293,G59785,G9111);
  nand GNAME12294(G12294,G9784,G59363);
  nand GNAME12295(G12295,G59785,G9112);
  nand GNAME12296(G12296,G59786,G9111);
  nand GNAME12297(G12297,G9784,G59362);
  nand GNAME12298(G12298,G59786,G9112);
  nand GNAME12299(G12299,G59787,G9111);
  nand GNAME12300(G12300,G9784,G59361);
  nand GNAME12301(G12301,G59787,G9112);
  nand GNAME12302(G12302,G59788,G9111);
  nand GNAME12303(G12303,G9784,G59360);
  nand GNAME12304(G12304,G59788,G9112);
  nand GNAME12305(G12305,G59789,G9111);
  nand GNAME12306(G12306,G59541,G9115);
  nand GNAME12307(G12307,G59533,G9118);
  nand GNAME12308(G12308,G59525,G9119);
  nand GNAME12309(G12309,G59517,G9121);
  nand GNAME12310(G12310,G59509,G9122);
  nand GNAME12311(G12311,G59501,G9124);
  nand GNAME12312(G12312,G59493,G9125);
  nand GNAME12313(G12313,G59485,G9127);
  nand GNAME12314(G12314,G59477,G9129);
  nand GNAME12315(G12315,G59469,G9130);
  nand GNAME12316(G12316,G59461,G9131);
  nand GNAME12317(G12317,G59453,G9132);
  nand GNAME12318(G12318,G59445,G9133);
  nand GNAME12319(G12319,G59437,G9134);
  nand GNAME12320(G12320,G59429,G9135);
  nand GNAME12321(G12321,G59549,G9136);
  nand GNAME12322(G12322,G59542,G9115);
  nand GNAME12323(G12323,G59534,G9118);
  nand GNAME12324(G12324,G59526,G9119);
  nand GNAME12325(G12325,G59518,G9121);
  nand GNAME12326(G12326,G59510,G9122);
  nand GNAME12327(G12327,G59502,G9124);
  nand GNAME12328(G12328,G59494,G9125);
  nand GNAME12329(G12329,G59486,G9127);
  nand GNAME12330(G12330,G59478,G9129);
  nand GNAME12331(G12331,G59470,G9130);
  nand GNAME12332(G12332,G59462,G9131);
  nand GNAME12333(G12333,G59454,G9132);
  nand GNAME12334(G12334,G59446,G9133);
  nand GNAME12335(G12335,G59438,G9134);
  nand GNAME12336(G12336,G59430,G9135);
  nand GNAME12337(G12337,G59550,G9136);
  nand GNAME12338(G12338,G59543,G9115);
  nand GNAME12339(G12339,G59535,G9118);
  nand GNAME12340(G12340,G59527,G9119);
  nand GNAME12341(G12341,G59519,G9121);
  nand GNAME12342(G12342,G59511,G9122);
  nand GNAME12343(G12343,G59503,G9124);
  nand GNAME12344(G12344,G59495,G9125);
  nand GNAME12345(G12345,G59487,G9127);
  nand GNAME12346(G12346,G59479,G9129);
  nand GNAME12347(G12347,G59471,G9130);
  nand GNAME12348(G12348,G59463,G9131);
  nand GNAME12349(G12349,G59455,G9132);
  nand GNAME12350(G12350,G59447,G9133);
  nand GNAME12351(G12351,G59439,G9134);
  nand GNAME12352(G12352,G59431,G9135);
  nand GNAME12353(G12353,G59551,G9136);
  nand GNAME12354(G12354,G59544,G9115);
  nand GNAME12355(G12355,G59536,G9118);
  nand GNAME12356(G12356,G59528,G9119);
  nand GNAME12357(G12357,G59520,G9121);
  nand GNAME12358(G12358,G59512,G9122);
  nand GNAME12359(G12359,G59504,G9124);
  nand GNAME12360(G12360,G59496,G9125);
  nand GNAME12361(G12361,G59488,G9127);
  nand GNAME12362(G12362,G59480,G9129);
  nand GNAME12363(G12363,G59472,G9130);
  nand GNAME12364(G12364,G59464,G9131);
  nand GNAME12365(G12365,G59456,G9132);
  nand GNAME12366(G12366,G59448,G9133);
  nand GNAME12367(G12367,G59440,G9134);
  nand GNAME12368(G12368,G59432,G9135);
  nand GNAME12369(G12369,G59552,G9136);
  nand GNAME12370(G12370,G59545,G9115);
  nand GNAME12371(G12371,G59537,G9118);
  nand GNAME12372(G12372,G59529,G9119);
  nand GNAME12373(G12373,G59521,G9121);
  nand GNAME12374(G12374,G59513,G9122);
  nand GNAME12375(G12375,G59505,G9124);
  nand GNAME12376(G12376,G59497,G9125);
  nand GNAME12377(G12377,G59489,G9127);
  nand GNAME12378(G12378,G59481,G9129);
  nand GNAME12379(G12379,G59473,G9130);
  nand GNAME12380(G12380,G59465,G9131);
  nand GNAME12381(G12381,G59457,G9132);
  nand GNAME12382(G12382,G59449,G9133);
  nand GNAME12383(G12383,G59441,G9134);
  nand GNAME12384(G12384,G59433,G9135);
  nand GNAME12385(G12385,G59553,G9136);
  nand GNAME12386(G12386,G59554,G9136);
  nand GNAME12387(G12387,G59546,G9115);
  nand GNAME12388(G12388,G59538,G9118);
  nand GNAME12389(G12389,G59530,G9119);
  nand GNAME12390(G12390,G59522,G9121);
  nand GNAME12391(G12391,G59514,G9122);
  nand GNAME12392(G12392,G59506,G9124);
  nand GNAME12393(G12393,G59498,G9125);
  nand GNAME12394(G12394,G59490,G9127);
  nand GNAME12395(G12395,G59482,G9129);
  nand GNAME12396(G12396,G59474,G9130);
  nand GNAME12397(G12397,G59466,G9131);
  nand GNAME12398(G12398,G59458,G9132);
  nand GNAME12399(G12399,G59450,G9133);
  nand GNAME12400(G12400,G59442,G9134);
  nand GNAME12401(G12401,G59434,G9135);
  nand GNAME12402(G12402,G59555,G9136);
  nand GNAME12403(G12403,G59547,G9115);
  nand GNAME12404(G12404,G59539,G9118);
  nand GNAME12405(G12405,G59531,G9119);
  nand GNAME12406(G12406,G59523,G9121);
  nand GNAME12407(G12407,G59515,G9122);
  nand GNAME12408(G12408,G59507,G9124);
  nand GNAME12409(G12409,G59499,G9125);
  nand GNAME12410(G12410,G59491,G9127);
  nand GNAME12411(G12411,G59483,G9129);
  nand GNAME12412(G12412,G59475,G9130);
  nand GNAME12413(G12413,G59467,G9131);
  nand GNAME12414(G12414,G59459,G9132);
  nand GNAME12415(G12415,G59451,G9133);
  nand GNAME12416(G12416,G59443,G9134);
  nand GNAME12417(G12417,G59435,G9135);
  nand GNAME12418(G12418,G59556,G9136);
  nand GNAME12419(G12419,G59548,G9115);
  nand GNAME12420(G12420,G59540,G9118);
  nand GNAME12421(G12421,G59532,G9119);
  nand GNAME12422(G12422,G59524,G9121);
  nand GNAME12423(G12423,G59516,G9122);
  nand GNAME12424(G12424,G59508,G9124);
  nand GNAME12425(G12425,G59500,G9125);
  nand GNAME12426(G12426,G59492,G9127);
  nand GNAME12427(G12427,G59484,G9129);
  nand GNAME12428(G12428,G59476,G9130);
  nand GNAME12429(G12429,G59468,G9131);
  nand GNAME12430(G12430,G59460,G9132);
  nand GNAME12431(G12431,G59452,G9133);
  nand GNAME12432(G12432,G59444,G9134);
  nand GNAME12433(G12433,G59436,G9135);
  not GNAME12434(G12434,G9137);
  nand GNAME12435(G12435,G59541,G9139);
  nand GNAME12436(G12436,G59533,G9140);
  nand GNAME12437(G12437,G59525,G9141);
  nand GNAME12438(G12438,G59517,G9143);
  nand GNAME12439(G12439,G59509,G9144);
  nand GNAME12440(G12440,G59501,G9145);
  nand GNAME12441(G12441,G59493,G9146);
  nand GNAME12442(G12442,G59485,G9148);
  nand GNAME12443(G12443,G59477,G9149);
  nand GNAME12444(G12444,G59469,G9150);
  nand GNAME12445(G12445,G59461,G9151);
  nand GNAME12446(G12446,G59453,G9153);
  nand GNAME12447(G12447,G59445,G9154);
  nand GNAME12448(G12448,G59437,G9155);
  nand GNAME12449(G12449,G59429,G9156);
  nand GNAME12450(G12450,G59549,G9157);
  nand GNAME12451(G12451,G59542,G9139);
  nand GNAME12452(G12452,G59534,G9140);
  nand GNAME12453(G12453,G59526,G9141);
  nand GNAME12454(G12454,G59518,G9143);
  nand GNAME12455(G12455,G59510,G9144);
  nand GNAME12456(G12456,G59502,G9145);
  nand GNAME12457(G12457,G59494,G9146);
  nand GNAME12458(G12458,G59486,G9148);
  nand GNAME12459(G12459,G59478,G9149);
  nand GNAME12460(G12460,G59470,G9150);
  nand GNAME12461(G12461,G59462,G9151);
  nand GNAME12462(G12462,G59454,G9153);
  nand GNAME12463(G12463,G59446,G9154);
  nand GNAME12464(G12464,G59438,G9155);
  nand GNAME12465(G12465,G59430,G9156);
  nand GNAME12466(G12466,G59550,G9157);
  nand GNAME12467(G12467,G59543,G9139);
  nand GNAME12468(G12468,G59535,G9140);
  nand GNAME12469(G12469,G59527,G9141);
  nand GNAME12470(G12470,G59519,G9143);
  nand GNAME12471(G12471,G59511,G9144);
  nand GNAME12472(G12472,G59503,G9145);
  nand GNAME12473(G12473,G59495,G9146);
  nand GNAME12474(G12474,G59487,G9148);
  nand GNAME12475(G12475,G59479,G9149);
  nand GNAME12476(G12476,G59471,G9150);
  nand GNAME12477(G12477,G59463,G9151);
  nand GNAME12478(G12478,G59455,G9153);
  nand GNAME12479(G12479,G59447,G9154);
  nand GNAME12480(G12480,G59439,G9155);
  nand GNAME12481(G12481,G59431,G9156);
  nand GNAME12482(G12482,G59551,G9157);
  nand GNAME12483(G12483,G59544,G9139);
  nand GNAME12484(G12484,G59536,G9140);
  nand GNAME12485(G12485,G59528,G9141);
  nand GNAME12486(G12486,G59520,G9143);
  nand GNAME12487(G12487,G59512,G9144);
  nand GNAME12488(G12488,G59504,G9145);
  nand GNAME12489(G12489,G59496,G9146);
  nand GNAME12490(G12490,G59488,G9148);
  nand GNAME12491(G12491,G59480,G9149);
  nand GNAME12492(G12492,G59472,G9150);
  nand GNAME12493(G12493,G59464,G9151);
  nand GNAME12494(G12494,G59456,G9153);
  nand GNAME12495(G12495,G59448,G9154);
  nand GNAME12496(G12496,G59440,G9155);
  nand GNAME12497(G12497,G59432,G9156);
  nand GNAME12498(G12498,G59552,G9157);
  nand GNAME12499(G12499,G59545,G9139);
  nand GNAME12500(G12500,G59537,G9140);
  nand GNAME12501(G12501,G59529,G9141);
  nand GNAME12502(G12502,G59521,G9143);
  nand GNAME12503(G12503,G59513,G9144);
  nand GNAME12504(G12504,G59505,G9145);
  nand GNAME12505(G12505,G59497,G9146);
  nand GNAME12506(G12506,G59489,G9148);
  nand GNAME12507(G12507,G59481,G9149);
  nand GNAME12508(G12508,G59473,G9150);
  nand GNAME12509(G12509,G59465,G9151);
  nand GNAME12510(G12510,G59457,G9153);
  nand GNAME12511(G12511,G59449,G9154);
  nand GNAME12512(G12512,G59441,G9155);
  nand GNAME12513(G12513,G59433,G9156);
  nand GNAME12514(G12514,G59553,G9157);
  nand GNAME12515(G12515,G59554,G9157);
  nand GNAME12516(G12516,G59546,G9139);
  nand GNAME12517(G12517,G59538,G9140);
  nand GNAME12518(G12518,G59530,G9141);
  nand GNAME12519(G12519,G59522,G9143);
  nand GNAME12520(G12520,G59514,G9144);
  nand GNAME12521(G12521,G59506,G9145);
  nand GNAME12522(G12522,G59498,G9146);
  nand GNAME12523(G12523,G59490,G9148);
  nand GNAME12524(G12524,G59482,G9149);
  nand GNAME12525(G12525,G59474,G9150);
  nand GNAME12526(G12526,G59466,G9151);
  nand GNAME12527(G12527,G59458,G9153);
  nand GNAME12528(G12528,G59450,G9154);
  nand GNAME12529(G12529,G59442,G9155);
  nand GNAME12530(G12530,G59434,G9156);
  nand GNAME12531(G12531,G59555,G9157);
  nand GNAME12532(G12532,G59547,G9139);
  nand GNAME12533(G12533,G59539,G9140);
  nand GNAME12534(G12534,G59531,G9141);
  nand GNAME12535(G12535,G59523,G9143);
  nand GNAME12536(G12536,G59515,G9144);
  nand GNAME12537(G12537,G59507,G9145);
  nand GNAME12538(G12538,G59499,G9146);
  nand GNAME12539(G12539,G59491,G9148);
  nand GNAME12540(G12540,G59483,G9149);
  nand GNAME12541(G12541,G59475,G9150);
  nand GNAME12542(G12542,G59467,G9151);
  nand GNAME12543(G12543,G59459,G9153);
  nand GNAME12544(G12544,G59451,G9154);
  nand GNAME12545(G12545,G59443,G9155);
  nand GNAME12546(G12546,G59435,G9156);
  nand GNAME12547(G12547,G59556,G9157);
  nand GNAME12548(G12548,G59548,G9139);
  nand GNAME12549(G12549,G59540,G9140);
  nand GNAME12550(G12550,G59532,G9141);
  nand GNAME12551(G12551,G59524,G9143);
  nand GNAME12552(G12552,G59516,G9144);
  nand GNAME12553(G12553,G59508,G9145);
  nand GNAME12554(G12554,G59500,G9146);
  nand GNAME12555(G12555,G59492,G9148);
  nand GNAME12556(G12556,G59484,G9149);
  nand GNAME12557(G12557,G59476,G9150);
  nand GNAME12558(G12558,G59468,G9151);
  nand GNAME12559(G12559,G59460,G9153);
  nand GNAME12560(G12560,G59452,G9154);
  nand GNAME12561(G12561,G59444,G9155);
  nand GNAME12562(G12562,G59436,G9156);
  nand GNAME12563(G12563,G59541,G8987);
  nand GNAME12564(G12564,G59533,G8998);
  nand GNAME12565(G12565,G59525,G9006);
  nand GNAME12566(G12566,G59517,G9016);
  nand GNAME12567(G12567,G59509,G9025);
  nand GNAME12568(G12568,G59501,G9032);
  nand GNAME12569(G12569,G59493,G9039);
  nand GNAME12570(G12570,G59485,G9050);
  nand GNAME12571(G12571,G59477,G9057);
  nand GNAME12572(G12572,G59469,G9066);
  nand GNAME12573(G12573,G59461,G9073);
  nand GNAME12574(G12574,G59453,G9082);
  nand GNAME12575(G12575,G59445,G9089);
  nand GNAME12576(G12576,G59437,G9096);
  nand GNAME12577(G12577,G59429,G9103);
  nand GNAME12578(G12578,G59549,G8960);
  nand GNAME12579(G12579,G9597,G9598,G9599,G9600);
  nand GNAME12580(G12580,G59542,G8987);
  nand GNAME12581(G12581,G59534,G8998);
  nand GNAME12582(G12582,G59526,G9006);
  nand GNAME12583(G12583,G59518,G9016);
  nand GNAME12584(G12584,G59510,G9025);
  nand GNAME12585(G12585,G59502,G9032);
  nand GNAME12586(G12586,G59494,G9039);
  nand GNAME12587(G12587,G59486,G9050);
  nand GNAME12588(G12588,G59478,G9057);
  nand GNAME12589(G12589,G59470,G9066);
  nand GNAME12590(G12590,G59462,G9073);
  nand GNAME12591(G12591,G59454,G9082);
  nand GNAME12592(G12592,G59446,G9089);
  nand GNAME12593(G12593,G59438,G9096);
  nand GNAME12594(G12594,G59430,G9103);
  nand GNAME12595(G12595,G59550,G8960);
  nand GNAME12596(G12596,G9601,G9602,G9603,G9604);
  nand GNAME12597(G12597,G59543,G8987);
  nand GNAME12598(G12598,G59535,G8998);
  nand GNAME12599(G12599,G59527,G9006);
  nand GNAME12600(G12600,G59519,G9016);
  nand GNAME12601(G12601,G59511,G9025);
  nand GNAME12602(G12602,G59503,G9032);
  nand GNAME12603(G12603,G59495,G9039);
  nand GNAME12604(G12604,G59487,G9050);
  nand GNAME12605(G12605,G59479,G9057);
  nand GNAME12606(G12606,G59471,G9066);
  nand GNAME12607(G12607,G59463,G9073);
  nand GNAME12608(G12608,G59455,G9082);
  nand GNAME12609(G12609,G59447,G9089);
  nand GNAME12610(G12610,G59439,G9096);
  nand GNAME12611(G12611,G59431,G9103);
  nand GNAME12612(G12612,G59551,G8960);
  nand GNAME12613(G12613,G9605,G9606,G9607,G9608);
  nand GNAME12614(G12614,G59544,G8987);
  nand GNAME12615(G12615,G59536,G8998);
  nand GNAME12616(G12616,G59528,G9006);
  nand GNAME12617(G12617,G59520,G9016);
  nand GNAME12618(G12618,G59512,G9025);
  nand GNAME12619(G12619,G59504,G9032);
  nand GNAME12620(G12620,G59496,G9039);
  nand GNAME12621(G12621,G59488,G9050);
  nand GNAME12622(G12622,G59480,G9057);
  nand GNAME12623(G12623,G59472,G9066);
  nand GNAME12624(G12624,G59464,G9073);
  nand GNAME12625(G12625,G59456,G9082);
  nand GNAME12626(G12626,G59448,G9089);
  nand GNAME12627(G12627,G59440,G9096);
  nand GNAME12628(G12628,G59432,G9103);
  nand GNAME12629(G12629,G59552,G8960);
  nand GNAME12630(G12630,G9609,G9610,G9611,G9612);
  nand GNAME12631(G12631,G59545,G8987);
  nand GNAME12632(G12632,G59537,G8998);
  nand GNAME12633(G12633,G59529,G9006);
  nand GNAME12634(G12634,G59521,G9016);
  nand GNAME12635(G12635,G59513,G9025);
  nand GNAME12636(G12636,G59505,G9032);
  nand GNAME12637(G12637,G59497,G9039);
  nand GNAME12638(G12638,G59489,G9050);
  nand GNAME12639(G12639,G59481,G9057);
  nand GNAME12640(G12640,G59473,G9066);
  nand GNAME12641(G12641,G59465,G9073);
  nand GNAME12642(G12642,G59457,G9082);
  nand GNAME12643(G12643,G59449,G9089);
  nand GNAME12644(G12644,G59441,G9096);
  nand GNAME12645(G12645,G59433,G9103);
  nand GNAME12646(G12646,G59553,G8960);
  nand GNAME12647(G12647,G9613,G9614,G9615,G9616);
  nand GNAME12648(G12648,G59554,G8960);
  nand GNAME12649(G12649,G59546,G8987);
  nand GNAME12650(G12650,G59538,G8998);
  nand GNAME12651(G12651,G59530,G9006);
  nand GNAME12652(G12652,G59522,G9016);
  nand GNAME12653(G12653,G59514,G9025);
  nand GNAME12654(G12654,G59506,G9032);
  nand GNAME12655(G12655,G59498,G9039);
  nand GNAME12656(G12656,G59490,G9050);
  nand GNAME12657(G12657,G59482,G9057);
  nand GNAME12658(G12658,G59474,G9066);
  nand GNAME12659(G12659,G59466,G9073);
  nand GNAME12660(G12660,G59458,G9082);
  nand GNAME12661(G12661,G59450,G9089);
  nand GNAME12662(G12662,G59442,G9096);
  nand GNAME12663(G12663,G59434,G9103);
  nand GNAME12664(G12664,G9617,G9618,G9619,G9620);
  nand GNAME12665(G12665,G59555,G8960);
  nand GNAME12666(G12666,G59547,G8987);
  nand GNAME12667(G12667,G59539,G8998);
  nand GNAME12668(G12668,G59531,G9006);
  nand GNAME12669(G12669,G59523,G9016);
  nand GNAME12670(G12670,G59515,G9025);
  nand GNAME12671(G12671,G59507,G9032);
  nand GNAME12672(G12672,G59499,G9039);
  nand GNAME12673(G12673,G59491,G9050);
  nand GNAME12674(G12674,G59483,G9057);
  nand GNAME12675(G12675,G59475,G9066);
  nand GNAME12676(G12676,G59467,G9073);
  nand GNAME12677(G12677,G59459,G9082);
  nand GNAME12678(G12678,G59451,G9089);
  nand GNAME12679(G12679,G59443,G9096);
  nand GNAME12680(G12680,G59435,G9103);
  nand GNAME12681(G12681,G9621,G9622,G9623,G9624);
  nand GNAME12682(G12682,G59556,G8960);
  nand GNAME12683(G12683,G59548,G8987);
  nand GNAME12684(G12684,G59540,G8998);
  nand GNAME12685(G12685,G59532,G9006);
  nand GNAME12686(G12686,G59524,G9016);
  nand GNAME12687(G12687,G59516,G9025);
  nand GNAME12688(G12688,G59508,G9032);
  nand GNAME12689(G12689,G59500,G9039);
  nand GNAME12690(G12690,G59492,G9050);
  nand GNAME12691(G12691,G59484,G9057);
  nand GNAME12692(G12692,G59476,G9066);
  nand GNAME12693(G12693,G59468,G9073);
  nand GNAME12694(G12694,G59460,G9082);
  nand GNAME12695(G12695,G59452,G9089);
  nand GNAME12696(G12696,G59444,G9096);
  nand GNAME12697(G12697,G59436,G9103);
  nand GNAME12698(G12698,G9625,G9626,G9627,G9628);
  nand GNAME12699(G12699,G59541,G9160);
  nand GNAME12700(G12700,G59533,G9163);
  nand GNAME12701(G12701,G59525,G9165);
  nand GNAME12702(G12702,G59517,G9168);
  nand GNAME12703(G12703,G59509,G9169);
  nand GNAME12704(G12704,G59501,G9170);
  nand GNAME12705(G12705,G59493,G9171);
  nand GNAME12706(G12706,G59485,G9173);
  nand GNAME12707(G12707,G59477,G9174);
  nand GNAME12708(G12708,G59469,G9175);
  nand GNAME12709(G12709,G59461,G9176);
  nand GNAME12710(G12710,G59453,G9178);
  nand GNAME12711(G12711,G59445,G9179);
  nand GNAME12712(G12712,G59437,G9180);
  nand GNAME12713(G12713,G59429,G9181);
  nand GNAME12714(G12714,G59549,G9182);
  nand GNAME12715(G12715,G9629,G9630,G9631,G9632);
  nand GNAME12716(G12716,G59542,G9160);
  nand GNAME12717(G12717,G59534,G9163);
  nand GNAME12718(G12718,G59526,G9165);
  nand GNAME12719(G12719,G59518,G9168);
  nand GNAME12720(G12720,G59510,G9169);
  nand GNAME12721(G12721,G59502,G9170);
  nand GNAME12722(G12722,G59494,G9171);
  nand GNAME12723(G12723,G59486,G9173);
  nand GNAME12724(G12724,G59478,G9174);
  nand GNAME12725(G12725,G59470,G9175);
  nand GNAME12726(G12726,G59462,G9176);
  nand GNAME12727(G12727,G59454,G9178);
  nand GNAME12728(G12728,G59446,G9179);
  nand GNAME12729(G12729,G59438,G9180);
  nand GNAME12730(G12730,G59430,G9181);
  nand GNAME12731(G12731,G59550,G9182);
  nand GNAME12732(G12732,G9633,G9634,G9635,G9636);
  nand GNAME12733(G12733,G59543,G9160);
  nand GNAME12734(G12734,G59535,G9163);
  nand GNAME12735(G12735,G59527,G9165);
  nand GNAME12736(G12736,G59519,G9168);
  nand GNAME12737(G12737,G59511,G9169);
  nand GNAME12738(G12738,G59503,G9170);
  nand GNAME12739(G12739,G59495,G9171);
  nand GNAME12740(G12740,G59487,G9173);
  nand GNAME12741(G12741,G59479,G9174);
  nand GNAME12742(G12742,G59471,G9175);
  nand GNAME12743(G12743,G59463,G9176);
  nand GNAME12744(G12744,G59455,G9178);
  nand GNAME12745(G12745,G59447,G9179);
  nand GNAME12746(G12746,G59439,G9180);
  nand GNAME12747(G12747,G59431,G9181);
  nand GNAME12748(G12748,G59551,G9182);
  nand GNAME12749(G12749,G9637,G9638,G9639,G9640);
  nand GNAME12750(G12750,G59544,G9160);
  nand GNAME12751(G12751,G59536,G9163);
  nand GNAME12752(G12752,G59528,G9165);
  nand GNAME12753(G12753,G59520,G9168);
  nand GNAME12754(G12754,G59512,G9169);
  nand GNAME12755(G12755,G59504,G9170);
  nand GNAME12756(G12756,G59496,G9171);
  nand GNAME12757(G12757,G59488,G9173);
  nand GNAME12758(G12758,G59480,G9174);
  nand GNAME12759(G12759,G59472,G9175);
  nand GNAME12760(G12760,G59464,G9176);
  nand GNAME12761(G12761,G59456,G9178);
  nand GNAME12762(G12762,G59448,G9179);
  nand GNAME12763(G12763,G59440,G9180);
  nand GNAME12764(G12764,G59432,G9181);
  nand GNAME12765(G12765,G59552,G9182);
  nand GNAME12766(G12766,G9641,G9642,G9643,G9644);
  nand GNAME12767(G12767,G59545,G9160);
  nand GNAME12768(G12768,G59537,G9163);
  nand GNAME12769(G12769,G59529,G9165);
  nand GNAME12770(G12770,G59521,G9168);
  nand GNAME12771(G12771,G59513,G9169);
  nand GNAME12772(G12772,G59505,G9170);
  nand GNAME12773(G12773,G59497,G9171);
  nand GNAME12774(G12774,G59489,G9173);
  nand GNAME12775(G12775,G59481,G9174);
  nand GNAME12776(G12776,G59473,G9175);
  nand GNAME12777(G12777,G59465,G9176);
  nand GNAME12778(G12778,G59457,G9178);
  nand GNAME12779(G12779,G59449,G9179);
  nand GNAME12780(G12780,G59441,G9180);
  nand GNAME12781(G12781,G59433,G9181);
  nand GNAME12782(G12782,G59553,G9182);
  nand GNAME12783(G12783,G9645,G9646,G9647,G9648);
  nand GNAME12784(G12784,G59554,G9182);
  nand GNAME12785(G12785,G59546,G9160);
  nand GNAME12786(G12786,G59538,G9163);
  nand GNAME12787(G12787,G59530,G9165);
  nand GNAME12788(G12788,G59522,G9168);
  nand GNAME12789(G12789,G59514,G9169);
  nand GNAME12790(G12790,G59506,G9170);
  nand GNAME12791(G12791,G59498,G9171);
  nand GNAME12792(G12792,G59490,G9173);
  nand GNAME12793(G12793,G59482,G9174);
  nand GNAME12794(G12794,G59474,G9175);
  nand GNAME12795(G12795,G59466,G9176);
  nand GNAME12796(G12796,G59458,G9178);
  nand GNAME12797(G12797,G59450,G9179);
  nand GNAME12798(G12798,G59442,G9180);
  nand GNAME12799(G12799,G59434,G9181);
  nand GNAME12800(G12800,G9649,G9650,G9651,G9652);
  nand GNAME12801(G12801,G59555,G9182);
  nand GNAME12802(G12802,G59547,G9160);
  nand GNAME12803(G12803,G59539,G9163);
  nand GNAME12804(G12804,G59531,G9165);
  nand GNAME12805(G12805,G59523,G9168);
  nand GNAME12806(G12806,G59515,G9169);
  nand GNAME12807(G12807,G59507,G9170);
  nand GNAME12808(G12808,G59499,G9171);
  nand GNAME12809(G12809,G59491,G9173);
  nand GNAME12810(G12810,G59483,G9174);
  nand GNAME12811(G12811,G59475,G9175);
  nand GNAME12812(G12812,G59467,G9176);
  nand GNAME12813(G12813,G59459,G9178);
  nand GNAME12814(G12814,G59451,G9179);
  nand GNAME12815(G12815,G59443,G9180);
  nand GNAME12816(G12816,G59435,G9181);
  nand GNAME12817(G12817,G9653,G9654,G9655,G9656);
  nand GNAME12818(G12818,G59556,G9182);
  nand GNAME12819(G12819,G59548,G9160);
  nand GNAME12820(G12820,G59540,G9163);
  nand GNAME12821(G12821,G59532,G9165);
  nand GNAME12822(G12822,G59524,G9168);
  nand GNAME12823(G12823,G59516,G9169);
  nand GNAME12824(G12824,G59508,G9170);
  nand GNAME12825(G12825,G59500,G9171);
  nand GNAME12826(G12826,G59492,G9173);
  nand GNAME12827(G12827,G59484,G9174);
  nand GNAME12828(G12828,G59476,G9175);
  nand GNAME12829(G12829,G59468,G9176);
  nand GNAME12830(G12830,G59460,G9178);
  nand GNAME12831(G12831,G59452,G9179);
  nand GNAME12832(G12832,G59444,G9180);
  nand GNAME12833(G12833,G59436,G9181);
  nand GNAME12834(G12834,G9657,G9658,G9659,G9660);
  nand GNAME12835(G12835,G9805,G9782,G9791);
  or GNAME12836(G12836,G9236,G9237);
  nand GNAME12837(G12837,G8824,G22755);
  nand GNAME12838(G12838,G12836,G21971);
  nand GNAME12839(G12839,G12835,G59576);
  nand GNAME12840(G12840,G21709,G9184);
  nand GNAME12841(G12841,G59767,G9186);
  nand GNAME12842(G12842,G8824,G22756);
  nand GNAME12843(G12843,G12836,G22006);
  nand GNAME12844(G12844,G12835,G59575);
  nand GNAME12845(G12845,G21666,G9184);
  nand GNAME12846(G12846,G59766,G9186);
  nand GNAME12847(G12847,G8824,G21996);
  nand GNAME12848(G12848,G12836,G21996);
  nand GNAME12849(G12849,G12835,G59574);
  nand GNAME12850(G12850,G21667,G9184);
  nand GNAME12851(G12851,G59765,G9186);
  nand GNAME12852(G12852,G8824,G21938);
  nand GNAME12853(G12853,G12836,G21938);
  nand GNAME12854(G12854,G12835,G59573);
  nand GNAME12855(G12855,G21633,G9184);
  nand GNAME12856(G12856,G59764,G9186);
  nand GNAME12857(G12857,G8824,G22010);
  nand GNAME12858(G12858,G12836,G22010);
  nand GNAME12859(G12859,G12835,G59572);
  nand GNAME12860(G12860,G21668,G9184);
  nand GNAME12861(G12861,G59763,G9186);
  nand GNAME12862(G12862,G8824,G22013);
  nand GNAME12863(G12863,G12836,G22013);
  nand GNAME12864(G12864,G12835,G59571);
  nand GNAME12865(G12865,G21669,G9184);
  nand GNAME12866(G12866,G59762,G9186);
  nand GNAME12867(G12867,G12836,G21998);
  nand GNAME12868(G12868,G12835,G59598);
  nand GNAME12869(G12869,G21700,G9184);
  nand GNAME12870(G12870,G59789,G9186);
  nand GNAME12871(G12871,G8824,G22757);
  nand GNAME12872(G12872,G12836,G21937);
  nand GNAME12873(G12873,G12835,G59597);
  nand GNAME12874(G12874,G21632,G9184);
  nand GNAME12875(G12875,G59788,G9186);
  nand GNAME12876(G12876,G8824,G21997);
  nand GNAME12877(G12877,G12836,G21997);
  nand GNAME12878(G12878,G12835,G59570);
  nand GNAME12879(G12879,G59761,G9186);
  nand GNAME12880(G12880,G21670,G9184);
  nand GNAME12881(G12881,G8824,G22758);
  nand GNAME12882(G12882,G12836,G21985);
  nand GNAME12883(G12883,G12835,G59596);
  nand GNAME12884(G12884,G21686,G9184);
  nand GNAME12885(G12885,G59787,G9186);
  nand GNAME12886(G12886,G8824,G22759);
  nand GNAME12887(G12887,G12836,G21986);
  nand GNAME12888(G12888,G12835,G59595);
  nand GNAME12889(G12889,G21687,G9184);
  nand GNAME12890(G12890,G59786,G9186);
  nand GNAME12891(G12891,G8824,G22760);
  nand GNAME12892(G12892,G12836,G21987);
  nand GNAME12893(G12893,G12835,G59594);
  nand GNAME12894(G12894,G21688,G9184);
  nand GNAME12895(G12895,G59785,G9186);
  nand GNAME12896(G12896,G8824,G22761);
  nand GNAME12897(G12897,G12836,G21988);
  nand GNAME12898(G12898,G12835,G59593);
  nand GNAME12899(G12899,G21689,G9184);
  nand GNAME12900(G12900,G59784,G9186);
  nand GNAME12901(G12901,G8824,G22762);
  nand GNAME12902(G12902,G12836,G21989);
  nand GNAME12903(G12903,G12835,G59592);
  nand GNAME12904(G12904,G21690,G9184);
  nand GNAME12905(G12905,G59783,G9186);
  nand GNAME12906(G12906,G8824,G22763);
  nand GNAME12907(G12907,G12836,G22027);
  nand GNAME12908(G12908,G12835,G59591);
  nand GNAME12909(G12909,G21691,G9184);
  nand GNAME12910(G12910,G59782,G9186);
  nand GNAME12911(G12911,G8824,G22764);
  nand GNAME12912(G12912,G12836,G22030);
  nand GNAME12913(G12913,G12835,G59590);
  nand GNAME12914(G12914,G21692,G9184);
  nand GNAME12915(G12915,G59781,G9186);
  nand GNAME12916(G12916,G8824,G22765);
  nand GNAME12917(G12917,G12836,G22033);
  nand GNAME12918(G12918,G12835,G59589);
  nand GNAME12919(G12919,G21693,G9184);
  nand GNAME12920(G12920,G59780,G9186);
  nand GNAME12921(G12921,G8824,G22766);
  nand GNAME12922(G12922,G12836,G22036);
  nand GNAME12923(G12923,G12835,G59588);
  nand GNAME12924(G12924,G21694,G9184);
  nand GNAME12925(G12925,G59779,G9186);
  nand GNAME12926(G12926,G8824,G22767);
  nand GNAME12927(G12927,G12836,G22039);
  nand GNAME12928(G12928,G12835,G59587);
  nand GNAME12929(G12929,G21695,G9184);
  nand GNAME12930(G12930,G59778,G9186);
  nand GNAME12931(G12931,G8824,G21936);
  nand GNAME12932(G12932,G12836,G21936);
  nand GNAME12933(G12933,G12835,G59569);
  nand GNAME12934(G12934,G59760,G9186);
  nand GNAME12935(G12935,G21631,G9184);
  nand GNAME12936(G12936,G8824,G22768);
  nand GNAME12937(G12937,G12836,G22045);
  nand GNAME12938(G12938,G12835,G59586);
  nand GNAME12939(G12939,G21696,G9184);
  nand GNAME12940(G12940,G59777,G9186);
  nand GNAME12941(G12941,G8824,G22769);
  nand GNAME12942(G12942,G12836,G22048);
  nand GNAME12943(G12943,G12835,G59585);
  nand GNAME12944(G12944,G21697,G9184);
  nand GNAME12945(G12945,G59776,G9186);
  nand GNAME12946(G12946,G8824,G22770);
  nand GNAME12947(G12947,G12836,G22051);
  nand GNAME12948(G12948,G12835,G59584);
  nand GNAME12949(G12949,G21698,G9184);
  nand GNAME12950(G12950,G59775,G9186);
  nand GNAME12951(G12951,G8824,G22783);
  nand GNAME12952(G12952,G12836,G21990);
  nand GNAME12953(G12953,G12835,G59583);
  nand GNAME12954(G12954,G21726,G9184);
  nand GNAME12955(G12955,G59774,G9186);
  nand GNAME12956(G12956,G8824,G22720);
  nand GNAME12957(G12957,G12836,G21991);
  nand GNAME12958(G12958,G12835,G59582);
  nand GNAME12959(G12959,G21729,G9184);
  nand GNAME12960(G12960,G59773,G9186);
  nand GNAME12961(G12961,G8824,G22785);
  nand GNAME12962(G12962,G12836,G21935);
  nand GNAME12963(G12963,G12835,G59581);
  nand GNAME12964(G12964,G21701,G9184);
  nand GNAME12965(G12965,G59772,G9186);
  nand GNAME12966(G12966,G8824,G22786);
  nand GNAME12967(G12967,G12836,G21992);
  nand GNAME12968(G12968,G12835,G59580);
  nand GNAME12969(G12969,G21733,G9184);
  nand GNAME12970(G12970,G59771,G9186);
  nand GNAME12971(G12971,G8824,G22787);
  nand GNAME12972(G12972,G12836,G21993);
  nand GNAME12973(G12973,G12835,G59579);
  nand GNAME12974(G12974,G21736,G9184);
  nand GNAME12975(G12975,G59770,G9186);
  nand GNAME12976(G12976,G8824,G22788);
  nand GNAME12977(G12977,G12836,G21994);
  nand GNAME12978(G12978,G12835,G59578);
  nand GNAME12979(G12979,G21702,G9184);
  nand GNAME12980(G12980,G59769,G9186);
  nand GNAME12981(G12981,G8824,G22789);
  nand GNAME12982(G12982,G12836,G21934);
  nand GNAME12983(G12983,G12835,G59577);
  nand GNAME12984(G12984,G21630,G9184);
  nand GNAME12985(G12985,G59768,G9186);
  nand GNAME12986(G12986,G8824,G22042);
  nand GNAME12987(G12987,G12836,G22042);
  nand GNAME12988(G12988,G12835,G59568);
  nand GNAME12989(G12989,G21723,G9184);
  nand GNAME12990(G12990,G59759,G9186);
  nand GNAME12991(G12991,G8824,G21995);
  nand GNAME12992(G12992,G12836,G21995);
  nand GNAME12993(G12993,G12835,G59567);
  nand GNAME12994(G12994,G21699,G9184);
  nand GNAME12995(G12995,G59758,G9186);
  nand GNAME12996(G12996,G59541,G11268);
  nand GNAME12997(G12997,G59533,G11329);
  nand GNAME12998(G12998,G59525,G11390);
  nand GNAME12999(G12999,G59517,G11451);
  nand GNAME13000(G13000,G59509,G11512);
  nand GNAME13001(G13001,G59501,G11573);
  nand GNAME13002(G13002,G59493,G11634);
  nand GNAME13003(G13003,G59485,G11695);
  nand GNAME13004(G13004,G59477,G11756);
  nand GNAME13005(G13005,G59469,G11817);
  nand GNAME13006(G13006,G59461,G11878);
  nand GNAME13007(G13007,G59453,G11939);
  nand GNAME13008(G13008,G59445,G12000);
  nand GNAME13009(G13009,G59437,G12061);
  nand GNAME13010(G13010,G59429,G12122);
  nand GNAME13011(G13011,G59549,G11186);
  nand GNAME13012(G13012,G9670,G9671,G9672,G9673);
  nand GNAME13013(G13013,G59541,G9214);
  nand GNAME13014(G13014,G59533,G9216);
  nand GNAME13015(G13015,G59525,G9218);
  nand GNAME13016(G13016,G59517,G9221);
  nand GNAME13017(G13017,G59509,G9222);
  nand GNAME13018(G13018,G59501,G9223);
  nand GNAME13019(G13019,G59493,G9224);
  nand GNAME13020(G13020,G59485,G9226);
  nand GNAME13021(G13021,G59477,G9227);
  nand GNAME13022(G13022,G59469,G9228);
  nand GNAME13023(G13023,G59461,G9229);
  nand GNAME13024(G13024,G59453,G9231);
  nand GNAME13025(G13025,G59445,G9232);
  nand GNAME13026(G13026,G59437,G9233);
  nand GNAME13027(G13027,G59429,G9234);
  nand GNAME13028(G13028,G59549,G9235);
  nand GNAME13029(G13029,G9666,G9667,G9668,G9669);
  nand GNAME13030(G13030,G59541,G9190);
  nand GNAME13031(G13031,G59533,G9193);
  nand GNAME13032(G13032,G59525,G9194);
  nand GNAME13033(G13033,G59517,G9196);
  nand GNAME13034(G13034,G59509,G9198);
  nand GNAME13035(G13035,G59501,G9199);
  nand GNAME13036(G13036,G59493,G9200);
  nand GNAME13037(G13037,G59485,G9202);
  nand GNAME13038(G13038,G59477,G9203);
  nand GNAME13039(G13039,G59469,G9205);
  nand GNAME13040(G13040,G59461,G9206);
  nand GNAME13041(G13041,G59453,G9207);
  nand GNAME13042(G13042,G59445,G9208);
  nand GNAME13043(G13043,G59437,G9209);
  nand GNAME13044(G13044,G59429,G9210);
  nand GNAME13045(G13045,G59549,G9211);
  nand GNAME13046(G13046,G9662,G9663,G9664,G9665);
  nand GNAME13047(G13047,G9184,G21928);
  nand GNAME13048(G13048,G13046,G8824);
  nand GNAME13049(G13049,G13029,G9236);
  nand GNAME13050(G13050,G13012,G9237);
  nand GNAME13051(G13051,G59542,G11268);
  nand GNAME13052(G13052,G59534,G11329);
  nand GNAME13053(G13053,G59526,G11390);
  nand GNAME13054(G13054,G59518,G11451);
  nand GNAME13055(G13055,G59510,G11512);
  nand GNAME13056(G13056,G59502,G11573);
  nand GNAME13057(G13057,G59494,G11634);
  nand GNAME13058(G13058,G59486,G11695);
  nand GNAME13059(G13059,G59478,G11756);
  nand GNAME13060(G13060,G59470,G11817);
  nand GNAME13061(G13061,G59462,G11878);
  nand GNAME13062(G13062,G59454,G11939);
  nand GNAME13063(G13063,G59446,G12000);
  nand GNAME13064(G13064,G59438,G12061);
  nand GNAME13065(G13065,G59430,G12122);
  nand GNAME13066(G13066,G59550,G11186);
  nand GNAME13067(G13067,G9682,G9683,G9684,G9685);
  nand GNAME13068(G13068,G59542,G9214);
  nand GNAME13069(G13069,G59534,G9216);
  nand GNAME13070(G13070,G59526,G9218);
  nand GNAME13071(G13071,G59518,G9221);
  nand GNAME13072(G13072,G59510,G9222);
  nand GNAME13073(G13073,G59502,G9223);
  nand GNAME13074(G13074,G59494,G9224);
  nand GNAME13075(G13075,G59486,G9226);
  nand GNAME13076(G13076,G59478,G9227);
  nand GNAME13077(G13077,G59470,G9228);
  nand GNAME13078(G13078,G59462,G9229);
  nand GNAME13079(G13079,G59454,G9231);
  nand GNAME13080(G13080,G59446,G9232);
  nand GNAME13081(G13081,G59438,G9233);
  nand GNAME13082(G13082,G59430,G9234);
  nand GNAME13083(G13083,G59550,G9235);
  nand GNAME13084(G13084,G9678,G9679,G9680,G9681);
  nand GNAME13085(G13085,G59542,G9190);
  nand GNAME13086(G13086,G59534,G9193);
  nand GNAME13087(G13087,G59526,G9194);
  nand GNAME13088(G13088,G59518,G9196);
  nand GNAME13089(G13089,G59510,G9198);
  nand GNAME13090(G13090,G59502,G9199);
  nand GNAME13091(G13091,G59494,G9200);
  nand GNAME13092(G13092,G59486,G9202);
  nand GNAME13093(G13093,G59478,G9203);
  nand GNAME13094(G13094,G59470,G9205);
  nand GNAME13095(G13095,G59462,G9206);
  nand GNAME13096(G13096,G59454,G9207);
  nand GNAME13097(G13097,G59446,G9208);
  nand GNAME13098(G13098,G59438,G9209);
  nand GNAME13099(G13099,G59430,G9210);
  nand GNAME13100(G13100,G59550,G9211);
  nand GNAME13101(G13101,G9674,G9675,G9676,G9677);
  nand GNAME13102(G13102,G9184,G21926);
  nand GNAME13103(G13103,G13101,G8824);
  nand GNAME13104(G13104,G13084,G9236);
  nand GNAME13105(G13105,G13067,G9237);
  nand GNAME13106(G13106,G59543,G11268);
  nand GNAME13107(G13107,G59535,G11329);
  nand GNAME13108(G13108,G59527,G11390);
  nand GNAME13109(G13109,G59519,G11451);
  nand GNAME13110(G13110,G59511,G11512);
  nand GNAME13111(G13111,G59503,G11573);
  nand GNAME13112(G13112,G59495,G11634);
  nand GNAME13113(G13113,G59487,G11695);
  nand GNAME13114(G13114,G59479,G11756);
  nand GNAME13115(G13115,G59471,G11817);
  nand GNAME13116(G13116,G59463,G11878);
  nand GNAME13117(G13117,G59455,G11939);
  nand GNAME13118(G13118,G59447,G12000);
  nand GNAME13119(G13119,G59439,G12061);
  nand GNAME13120(G13120,G59431,G12122);
  nand GNAME13121(G13121,G59551,G11186);
  nand GNAME13122(G13122,G9694,G9695,G9696,G9697);
  nand GNAME13123(G13123,G59543,G9214);
  nand GNAME13124(G13124,G59535,G9216);
  nand GNAME13125(G13125,G59527,G9218);
  nand GNAME13126(G13126,G59519,G9221);
  nand GNAME13127(G13127,G59511,G9222);
  nand GNAME13128(G13128,G59503,G9223);
  nand GNAME13129(G13129,G59495,G9224);
  nand GNAME13130(G13130,G59487,G9226);
  nand GNAME13131(G13131,G59479,G9227);
  nand GNAME13132(G13132,G59471,G9228);
  nand GNAME13133(G13133,G59463,G9229);
  nand GNAME13134(G13134,G59455,G9231);
  nand GNAME13135(G13135,G59447,G9232);
  nand GNAME13136(G13136,G59439,G9233);
  nand GNAME13137(G13137,G59431,G9234);
  nand GNAME13138(G13138,G59551,G9235);
  nand GNAME13139(G13139,G9690,G9691,G9692,G9693);
  nand GNAME13140(G13140,G59543,G9190);
  nand GNAME13141(G13141,G59535,G9193);
  nand GNAME13142(G13142,G59527,G9194);
  nand GNAME13143(G13143,G59519,G9196);
  nand GNAME13144(G13144,G59511,G9198);
  nand GNAME13145(G13145,G59503,G9199);
  nand GNAME13146(G13146,G59495,G9200);
  nand GNAME13147(G13147,G59487,G9202);
  nand GNAME13148(G13148,G59479,G9203);
  nand GNAME13149(G13149,G59471,G9205);
  nand GNAME13150(G13150,G59463,G9206);
  nand GNAME13151(G13151,G59455,G9207);
  nand GNAME13152(G13152,G59447,G9208);
  nand GNAME13153(G13153,G59439,G9209);
  nand GNAME13154(G13154,G59431,G9210);
  nand GNAME13155(G13155,G59551,G9211);
  nand GNAME13156(G13156,G9686,G9687,G9688,G9689);
  nand GNAME13157(G13157,G9184,G21929);
  nand GNAME13158(G13158,G13156,G8824);
  nand GNAME13159(G13159,G13139,G9236);
  nand GNAME13160(G13160,G13122,G9237);
  nand GNAME13161(G13161,G59544,G9214);
  nand GNAME13162(G13162,G59536,G9216);
  nand GNAME13163(G13163,G59528,G9218);
  nand GNAME13164(G13164,G59520,G9221);
  nand GNAME13165(G13165,G59512,G9222);
  nand GNAME13166(G13166,G59504,G9223);
  nand GNAME13167(G13167,G59496,G9224);
  nand GNAME13168(G13168,G59488,G9226);
  nand GNAME13169(G13169,G59480,G9227);
  nand GNAME13170(G13170,G59472,G9228);
  nand GNAME13171(G13171,G59464,G9229);
  nand GNAME13172(G13172,G59456,G9231);
  nand GNAME13173(G13173,G59448,G9232);
  nand GNAME13174(G13174,G59440,G9233);
  nand GNAME13175(G13175,G59432,G9234);
  nand GNAME13176(G13176,G59552,G9235);
  nand GNAME13177(G13177,G9706,G9707,G9708,G9709);
  nand GNAME13178(G13178,G59544,G9190);
  nand GNAME13179(G13179,G59536,G9193);
  nand GNAME13180(G13180,G59528,G9194);
  nand GNAME13181(G13181,G59520,G9196);
  nand GNAME13182(G13182,G59512,G9198);
  nand GNAME13183(G13183,G59504,G9199);
  nand GNAME13184(G13184,G59496,G9200);
  nand GNAME13185(G13185,G59488,G9202);
  nand GNAME13186(G13186,G59480,G9203);
  nand GNAME13187(G13187,G59472,G9205);
  nand GNAME13188(G13188,G59464,G9206);
  nand GNAME13189(G13189,G59456,G9207);
  nand GNAME13190(G13190,G59448,G9208);
  nand GNAME13191(G13191,G59440,G9209);
  nand GNAME13192(G13192,G59432,G9210);
  nand GNAME13193(G13193,G59552,G9211);
  nand GNAME13194(G13194,G9702,G9703,G9704,G9705);
  nand GNAME13195(G13195,G59544,G11268);
  nand GNAME13196(G13196,G59536,G11329);
  nand GNAME13197(G13197,G59528,G11390);
  nand GNAME13198(G13198,G59520,G11451);
  nand GNAME13199(G13199,G59512,G11512);
  nand GNAME13200(G13200,G59504,G11573);
  nand GNAME13201(G13201,G59496,G11634);
  nand GNAME13202(G13202,G59488,G11695);
  nand GNAME13203(G13203,G59480,G11756);
  nand GNAME13204(G13204,G59472,G11817);
  nand GNAME13205(G13205,G59464,G11878);
  nand GNAME13206(G13206,G59456,G11939);
  nand GNAME13207(G13207,G59448,G12000);
  nand GNAME13208(G13208,G59440,G12061);
  nand GNAME13209(G13209,G59432,G12122);
  nand GNAME13210(G13210,G59552,G11186);
  nand GNAME13211(G13211,G9698,G9699,G9700,G9701);
  or GNAME13212(G13212,G9883,G13982);
  nand GNAME13213(G13213,G9184,G21933);
  nand GNAME13214(G13214,G13211,G9237);
  nand GNAME13215(G13215,G13194,G8824);
  nand GNAME13216(G13216,G13177,G9236);
  nand GNAME13217(G13217,G59545,G9214);
  nand GNAME13218(G13218,G59537,G9216);
  nand GNAME13219(G13219,G59529,G9218);
  nand GNAME13220(G13220,G59521,G9221);
  nand GNAME13221(G13221,G59513,G9222);
  nand GNAME13222(G13222,G59505,G9223);
  nand GNAME13223(G13223,G59497,G9224);
  nand GNAME13224(G13224,G59489,G9226);
  nand GNAME13225(G13225,G59481,G9227);
  nand GNAME13226(G13226,G59473,G9228);
  nand GNAME13227(G13227,G59465,G9229);
  nand GNAME13228(G13228,G59457,G9231);
  nand GNAME13229(G13229,G59449,G9232);
  nand GNAME13230(G13230,G59441,G9233);
  nand GNAME13231(G13231,G59433,G9234);
  nand GNAME13232(G13232,G59553,G9235);
  nand GNAME13233(G13233,G9718,G9719,G9720,G9721);
  nand GNAME13234(G13234,G59545,G9190);
  nand GNAME13235(G13235,G59537,G9193);
  nand GNAME13236(G13236,G59529,G9194);
  nand GNAME13237(G13237,G59521,G9196);
  nand GNAME13238(G13238,G59513,G9198);
  nand GNAME13239(G13239,G59505,G9199);
  nand GNAME13240(G13240,G59497,G9200);
  nand GNAME13241(G13241,G59489,G9202);
  nand GNAME13242(G13242,G59481,G9203);
  nand GNAME13243(G13243,G59473,G9205);
  nand GNAME13244(G13244,G59465,G9206);
  nand GNAME13245(G13245,G59457,G9207);
  nand GNAME13246(G13246,G59449,G9208);
  nand GNAME13247(G13247,G59441,G9209);
  nand GNAME13248(G13248,G59433,G9210);
  nand GNAME13249(G13249,G59553,G9211);
  nand GNAME13250(G13250,G9714,G9715,G9716,G9717);
  nand GNAME13251(G13251,G59545,G11268);
  nand GNAME13252(G13252,G59537,G11329);
  nand GNAME13253(G13253,G59529,G11390);
  nand GNAME13254(G13254,G59521,G11451);
  nand GNAME13255(G13255,G59513,G11512);
  nand GNAME13256(G13256,G59505,G11573);
  nand GNAME13257(G13257,G59497,G11634);
  nand GNAME13258(G13258,G59489,G11695);
  nand GNAME13259(G13259,G59481,G11756);
  nand GNAME13260(G13260,G59473,G11817);
  nand GNAME13261(G13261,G59465,G11878);
  nand GNAME13262(G13262,G59457,G11939);
  nand GNAME13263(G13263,G59449,G12000);
  nand GNAME13264(G13264,G59441,G12061);
  nand GNAME13265(G13265,G59433,G12122);
  nand GNAME13266(G13266,G59553,G11186);
  nand GNAME13267(G13267,G9710,G9711,G9712,G9713);
  nand GNAME13268(G13268,G9184,G21931);
  nand GNAME13269(G13269,G13267,G9237);
  nand GNAME13270(G13270,G13250,G8824);
  nand GNAME13271(G13271,G13233,G9236);
  nand GNAME13272(G13272,G8781,G59558);
  nand GNAME13273(G13273,G59554,G9235);
  nand GNAME13274(G13274,G59546,G9214);
  nand GNAME13275(G13275,G59538,G9216);
  nand GNAME13276(G13276,G59530,G9218);
  nand GNAME13277(G13277,G59522,G9221);
  nand GNAME13278(G13278,G59514,G9222);
  nand GNAME13279(G13279,G59506,G9223);
  nand GNAME13280(G13280,G59498,G9224);
  nand GNAME13281(G13281,G59490,G9226);
  nand GNAME13282(G13282,G59482,G9227);
  nand GNAME13283(G13283,G59474,G9228);
  nand GNAME13284(G13284,G59466,G9229);
  nand GNAME13285(G13285,G59458,G9231);
  nand GNAME13286(G13286,G59450,G9232);
  nand GNAME13287(G13287,G59442,G9233);
  nand GNAME13288(G13288,G59434,G9234);
  nand GNAME13289(G13289,G9730,G9731,G9732,G9733);
  nand GNAME13290(G13290,G59554,G9211);
  nand GNAME13291(G13291,G59546,G9190);
  nand GNAME13292(G13292,G59538,G9193);
  nand GNAME13293(G13293,G59530,G9194);
  nand GNAME13294(G13294,G59522,G9196);
  nand GNAME13295(G13295,G59514,G9198);
  nand GNAME13296(G13296,G59506,G9199);
  nand GNAME13297(G13297,G59498,G9200);
  nand GNAME13298(G13298,G59490,G9202);
  nand GNAME13299(G13299,G59482,G9203);
  nand GNAME13300(G13300,G59474,G9205);
  nand GNAME13301(G13301,G59466,G9206);
  nand GNAME13302(G13302,G59458,G9207);
  nand GNAME13303(G13303,G59450,G9208);
  nand GNAME13304(G13304,G59442,G9209);
  nand GNAME13305(G13305,G59434,G9210);
  nand GNAME13306(G13306,G9726,G9727,G9728,G9729);
  nand GNAME13307(G13307,G59554,G11186);
  nand GNAME13308(G13308,G59546,G11268);
  nand GNAME13309(G13309,G59538,G11329);
  nand GNAME13310(G13310,G59530,G11390);
  nand GNAME13311(G13311,G59522,G11451);
  nand GNAME13312(G13312,G59514,G11512);
  nand GNAME13313(G13313,G59506,G11573);
  nand GNAME13314(G13314,G59498,G11634);
  nand GNAME13315(G13315,G59490,G11695);
  nand GNAME13316(G13316,G59482,G11756);
  nand GNAME13317(G13317,G59474,G11817);
  nand GNAME13318(G13318,G59466,G11878);
  nand GNAME13319(G13319,G59458,G11939);
  nand GNAME13320(G13320,G59450,G12000);
  nand GNAME13321(G13321,G59442,G12061);
  nand GNAME13322(G13322,G59434,G12122);
  nand GNAME13323(G13323,G9722,G9723,G9724,G9725);
  nand GNAME13324(G13324,G9184,G21932);
  nand GNAME13325(G13325,G13323,G9237);
  nand GNAME13326(G13326,G13306,G8824);
  nand GNAME13327(G13327,G13289,G9236);
  nand GNAME13328(G13328,G8781,G59559);
  nand GNAME13329(G13329,G59555,G9235);
  nand GNAME13330(G13330,G59547,G9214);
  nand GNAME13331(G13331,G59539,G9216);
  nand GNAME13332(G13332,G59531,G9218);
  nand GNAME13333(G13333,G59523,G9221);
  nand GNAME13334(G13334,G59515,G9222);
  nand GNAME13335(G13335,G59507,G9223);
  nand GNAME13336(G13336,G59499,G9224);
  nand GNAME13337(G13337,G59491,G9226);
  nand GNAME13338(G13338,G59483,G9227);
  nand GNAME13339(G13339,G59475,G9228);
  nand GNAME13340(G13340,G59467,G9229);
  nand GNAME13341(G13341,G59459,G9231);
  nand GNAME13342(G13342,G59451,G9232);
  nand GNAME13343(G13343,G59443,G9233);
  nand GNAME13344(G13344,G59435,G9234);
  nand GNAME13345(G13345,G9743,G9744,G9745,G9746);
  nand GNAME13346(G13346,G59555,G9211);
  nand GNAME13347(G13347,G59547,G9190);
  nand GNAME13348(G13348,G59539,G9193);
  nand GNAME13349(G13349,G59531,G9194);
  nand GNAME13350(G13350,G59523,G9196);
  nand GNAME13351(G13351,G59515,G9198);
  nand GNAME13352(G13352,G59507,G9199);
  nand GNAME13353(G13353,G59499,G9200);
  nand GNAME13354(G13354,G59491,G9202);
  nand GNAME13355(G13355,G59483,G9203);
  nand GNAME13356(G13356,G59475,G9205);
  nand GNAME13357(G13357,G59467,G9206);
  nand GNAME13358(G13358,G59459,G9207);
  nand GNAME13359(G13359,G59451,G9208);
  nand GNAME13360(G13360,G59443,G9209);
  nand GNAME13361(G13361,G59435,G9210);
  nand GNAME13362(G13362,G9739,G9740,G9741,G9742);
  nand GNAME13363(G13363,G59555,G11186);
  nand GNAME13364(G13364,G59547,G11268);
  nand GNAME13365(G13365,G59539,G11329);
  nand GNAME13366(G13366,G59531,G11390);
  nand GNAME13367(G13367,G59523,G11451);
  nand GNAME13368(G13368,G59515,G11512);
  nand GNAME13369(G13369,G59507,G11573);
  nand GNAME13370(G13370,G59499,G11634);
  nand GNAME13371(G13371,G59491,G11695);
  nand GNAME13372(G13372,G59483,G11756);
  nand GNAME13373(G13373,G59475,G11817);
  nand GNAME13374(G13374,G59467,G11878);
  nand GNAME13375(G13375,G59459,G11939);
  nand GNAME13376(G13376,G59451,G12000);
  nand GNAME13377(G13377,G59443,G12061);
  nand GNAME13378(G13378,G59435,G12122);
  nand GNAME13379(G13379,G9735,G9736,G9737,G9738);
  nand GNAME13380(G13380,G9184,G21927);
  nand GNAME13381(G13381,G13379,G9237);
  nand GNAME13382(G13382,G13362,G8824);
  nand GNAME13383(G13383,G13345,G9236);
  nand GNAME13384(G13384,G8781,G59560);
  nand GNAME13385(G13385,G59556,G9235);
  nand GNAME13386(G13386,G59548,G9214);
  nand GNAME13387(G13387,G59540,G9216);
  nand GNAME13388(G13388,G59532,G9218);
  nand GNAME13389(G13389,G59524,G9221);
  nand GNAME13390(G13390,G59516,G9222);
  nand GNAME13391(G13391,G59508,G9223);
  nand GNAME13392(G13392,G59500,G9224);
  nand GNAME13393(G13393,G59492,G9226);
  nand GNAME13394(G13394,G59484,G9227);
  nand GNAME13395(G13395,G59476,G9228);
  nand GNAME13396(G13396,G59468,G9229);
  nand GNAME13397(G13397,G59460,G9231);
  nand GNAME13398(G13398,G59452,G9232);
  nand GNAME13399(G13399,G59444,G9233);
  nand GNAME13400(G13400,G59436,G9234);
  nand GNAME13401(G13401,G9756,G9757,G9758,G9759);
  nand GNAME13402(G13402,G59556,G9211);
  nand GNAME13403(G13403,G59548,G9190);
  nand GNAME13404(G13404,G59540,G9193);
  nand GNAME13405(G13405,G59532,G9194);
  nand GNAME13406(G13406,G59524,G9196);
  nand GNAME13407(G13407,G59516,G9198);
  nand GNAME13408(G13408,G59508,G9199);
  nand GNAME13409(G13409,G59500,G9200);
  nand GNAME13410(G13410,G59492,G9202);
  nand GNAME13411(G13411,G59484,G9203);
  nand GNAME13412(G13412,G59476,G9205);
  nand GNAME13413(G13413,G59468,G9206);
  nand GNAME13414(G13414,G59460,G9207);
  nand GNAME13415(G13415,G59452,G9208);
  nand GNAME13416(G13416,G59444,G9209);
  nand GNAME13417(G13417,G59436,G9210);
  nand GNAME13418(G13418,G9752,G9753,G9754,G9755);
  nand GNAME13419(G13419,G59556,G11186);
  nand GNAME13420(G13420,G59548,G11268);
  nand GNAME13421(G13421,G59540,G11329);
  nand GNAME13422(G13422,G59532,G11390);
  nand GNAME13423(G13423,G59524,G11451);
  nand GNAME13424(G13424,G59516,G11512);
  nand GNAME13425(G13425,G59508,G11573);
  nand GNAME13426(G13426,G59500,G11634);
  nand GNAME13427(G13427,G59492,G11695);
  nand GNAME13428(G13428,G59484,G11756);
  nand GNAME13429(G13429,G59476,G11817);
  nand GNAME13430(G13430,G59468,G11878);
  nand GNAME13431(G13431,G59460,G11939);
  nand GNAME13432(G13432,G59452,G12000);
  nand GNAME13433(G13433,G59444,G12061);
  nand GNAME13434(G13434,G59436,G12122);
  nand GNAME13435(G13435,G9748,G9749,G9750,G9751);
  nand GNAME13436(G13436,G9184,G21930);
  nand GNAME13437(G13437,G13435,G9237);
  nand GNAME13438(G13438,G13418,G8824);
  nand GNAME13439(G13439,G13401,G9236);
  nand GNAME13440(G13440,G8781,G59561);
  nand GNAME13441(G13441,G8798,G9237,G59428,G8782,G9900);
  nand GNAME13442(G13442,G59554,G8856);
  or GNAME13443(G13443,G8787,G9917,G8750);
  nand GNAME13444(G13444,G8784,G59428,G8798,G13987);
  nand GNAME13445(G13445,G59555,G8856);
  nand GNAME13446(G13446,G8781,G9832);
  nand GNAME13447(G13447,G8791,G8887);
  nand GNAME13448(G13448,G9762,G13832,G13967,G8892,G9240);
  nand GNAME13449(G13449,G13448,G59428);
  nand GNAME13450(G13450,G59556,G8856);
  nand GNAME13451(G13451,G8852,G8860);
  nand GNAME13452(G13452,G9849,G8853);
  nand GNAME13453(G13453,G8780,G9951);
  nand GNAME13454(G13454,G13453,G13451,G13452);
  nand GNAME13455(G13455,G8746,G8792);
  nand GNAME13456(G13456,G8743,G8782);
  nand GNAME13457(G13457,G13456,G9783);
  nand GNAME13458(G13458,G13457,G8887);
  nand GNAME13459(G13459,G13455,G8827);
  nand GNAME13460(G13460,G8853,G8894);
  nand GNAME13461(G13461,G8792,G13454);
  nand GNAME13462(G13462,G8821,G8824);
  nand GNAME13463(G13463,G9763,G8895,G13461,G13462);
  nand GNAME13464(G13464,G13463,G59428);
  or GNAME13465(G13465,G8899,G8787);
  nand GNAME13466(G13466,G9807,G13441,G13465,G9241);
  nand GNAME13467(G13467,G9796,G9779);
  nand GNAME13468(G13468,G13467,G21709);
  nand GNAME13469(G13469,G13466,G59576);
  nand GNAME13470(G13470,G9780,G59608);
  nand GNAME13471(G13471,G8788,G59767);
  nand GNAME13472(G13472,G13467,G21666);
  nand GNAME13473(G13473,G13466,G59575);
  nand GNAME13474(G13474,G9780,G59607);
  nand GNAME13475(G13475,G8788,G59766);
  nand GNAME13476(G13476,G13467,G21667);
  nand GNAME13477(G13477,G13466,G59574);
  nand GNAME13478(G13478,G9780,G59606);
  nand GNAME13479(G13479,G8788,G59765);
  nand GNAME13480(G13480,G13467,G21633);
  nand GNAME13481(G13481,G13466,G59573);
  nand GNAME13482(G13482,G9780,G59605);
  nand GNAME13483(G13483,G8788,G59764);
  nand GNAME13484(G13484,G13467,G21668);
  nand GNAME13485(G13485,G13466,G59572);
  nand GNAME13486(G13486,G9780,G59604);
  nand GNAME13487(G13487,G8788,G59763);
  nand GNAME13488(G13488,G59428,G8871);
  nand GNAME13489(G13489,G13488,G8863);
  nand GNAME13490(G13490,G13489,G59557);
  nand GNAME13491(G13491,G13467,G21669);
  nand GNAME13492(G13492,G13466,G59571);
  nand GNAME13493(G13493,G9780,G59603);
  nand GNAME13494(G13494,G8788,G59762);
  nand GNAME13495(G13495,G13466,G59598);
  nand GNAME13496(G13496,G9780,G59630);
  nand GNAME13497(G13497,G8833,G21700);
  nand GNAME13498(G13498,G8788,G59789);
  nand GNAME13499(G13499,G13467,G21632);
  nand GNAME13500(G13500,G13466,G59597);
  nand GNAME13501(G13501,G9780,G59629);
  nand GNAME13502(G13502,G8788,G59788);
  nand GNAME13503(G13503,G12579,G8864);
  nand GNAME13504(G13504,G10830,G10831);
  nand GNAME13505(G13505,G13504,G59428);
  nand GNAME13506(G13506,G9183,G9238);
  or GNAME13507(G13507,G8902,G8787);
  nand GNAME13508(G13508,G13507,G9242,G13506,G9797,G10320);
  nand GNAME13509(G13509,G13508,G59558);
  nand GNAME13510(G13510,G13467,G21670);
  nand GNAME13511(G13511,G13466,G59570);
  nand GNAME13512(G13512,G9780,G59602);
  nand GNAME13513(G13513,G8788,G59761);
  nand GNAME13514(G13514,G13467,G21686);
  nand GNAME13515(G13515,G13466,G59596);
  nand GNAME13516(G13516,G9780,G59628);
  nand GNAME13517(G13517,G8788,G59787);
  nand GNAME13518(G13518,G12596,G8864);
  nand GNAME13519(G13519,G13467,G21687);
  nand GNAME13520(G13520,G13466,G59595);
  nand GNAME13521(G13521,G9780,G59627);
  nand GNAME13522(G13522,G8788,G59786);
  nand GNAME13523(G13523,G12613,G8864);
  nand GNAME13524(G13524,G13467,G21688);
  nand GNAME13525(G13525,G13466,G59594);
  nand GNAME13526(G13526,G9780,G59626);
  nand GNAME13527(G13527,G8788,G59785);
  nand GNAME13528(G13528,G12630,G8864);
  nand GNAME13529(G13529,G13467,G21689);
  nand GNAME13530(G13530,G13466,G59593);
  nand GNAME13531(G13531,G9780,G59625);
  nand GNAME13532(G13532,G8788,G59784);
  nand GNAME13533(G13533,G12647,G8864);
  nand GNAME13534(G13534,G13467,G21690);
  nand GNAME13535(G13535,G13466,G59592);
  nand GNAME13536(G13536,G9780,G59624);
  nand GNAME13537(G13537,G8788,G59783);
  nand GNAME13538(G13538,G12664,G8864);
  nand GNAME13539(G13539,G13467,G21691);
  nand GNAME13540(G13540,G13466,G59591);
  nand GNAME13541(G13541,G9780,G59623);
  nand GNAME13542(G13542,G8788,G59782);
  nand GNAME13543(G13543,G12681,G8864);
  nand GNAME13544(G13544,G13467,G21692);
  nand GNAME13545(G13545,G13466,G59590);
  nand GNAME13546(G13546,G9780,G59622);
  nand GNAME13547(G13547,G8788,G59781);
  nand GNAME13548(G13548,G12698,G8864);
  nand GNAME13549(G13549,G13467,G21693);
  nand GNAME13550(G13550,G13466,G59589);
  nand GNAME13551(G13551,G9780,G59621);
  nand GNAME13552(G13552,G8788,G59780);
  nand GNAME13553(G13553,G13467,G21694);
  nand GNAME13554(G13554,G13466,G59588);
  nand GNAME13555(G13555,G9780,G59620);
  nand GNAME13556(G13556,G8788,G59779);
  nand GNAME13557(G13557,G13467,G21695);
  nand GNAME13558(G13558,G13466,G59587);
  nand GNAME13559(G13559,G9780,G59619);
  nand GNAME13560(G13560,G8788,G59778);
  nand GNAME13561(G13561,G13508,G59559);
  nand GNAME13562(G13562,G13467,G21631);
  nand GNAME13563(G13563,G13466,G59569);
  nand GNAME13564(G13564,G9780,G59601);
  nand GNAME13565(G13565,G8788,G59760);
  nand GNAME13566(G13566,G13467,G21696);
  nand GNAME13567(G13567,G13466,G59586);
  nand GNAME13568(G13568,G9780,G59618);
  nand GNAME13569(G13569,G8788,G59777);
  nand GNAME13570(G13570,G13467,G21697);
  nand GNAME13571(G13571,G13466,G59585);
  nand GNAME13572(G13572,G9780,G59617);
  nand GNAME13573(G13573,G8788,G59776);
  nand GNAME13574(G13574,G13467,G21698);
  nand GNAME13575(G13575,G13466,G59584);
  nand GNAME13576(G13576,G9780,G59616);
  nand GNAME13577(G13577,G8788,G59775);
  nand GNAME13578(G13578,G13467,G21726);
  nand GNAME13579(G13579,G13466,G59583);
  nand GNAME13580(G13580,G9780,G59615);
  nand GNAME13581(G13581,G8788,G59774);
  nand GNAME13582(G13582,G13467,G21729);
  nand GNAME13583(G13583,G13466,G59582);
  nand GNAME13584(G13584,G9780,G59614);
  nand GNAME13585(G13585,G8788,G59773);
  nand GNAME13586(G13586,G13467,G21701);
  nand GNAME13587(G13587,G13466,G59581);
  nand GNAME13588(G13588,G9780,G59613);
  nand GNAME13589(G13589,G8788,G59772);
  nand GNAME13590(G13590,G13467,G21733);
  nand GNAME13591(G13591,G13466,G59580);
  nand GNAME13592(G13592,G9780,G59612);
  nand GNAME13593(G13593,G8788,G59771);
  nand GNAME13594(G13594,G13467,G21736);
  nand GNAME13595(G13595,G13466,G59579);
  nand GNAME13596(G13596,G9780,G59611);
  nand GNAME13597(G13597,G8788,G59770);
  nand GNAME13598(G13598,G13467,G21702);
  nand GNAME13599(G13599,G13466,G59578);
  nand GNAME13600(G13600,G9780,G59610);
  nand GNAME13601(G13601,G8788,G59769);
  nand GNAME13602(G13602,G13467,G21630);
  nand GNAME13603(G13603,G13466,G59577);
  nand GNAME13604(G13604,G9780,G59609);
  nand GNAME13605(G13605,G8788,G59768);
  nand GNAME13606(G13606,G13508,G59560);
  nand GNAME13607(G13607,G13467,G21723);
  nand GNAME13608(G13608,G13466,G59568);
  nand GNAME13609(G13609,G9780,G59600);
  nand GNAME13610(G13610,G8788,G59759);
  nand GNAME13611(G13611,G13508,G59561);
  nand GNAME13612(G13612,G13467,G21699);
  nand GNAME13613(G13613,G13466,G59567);
  nand GNAME13614(G13614,G9780,G59599);
  nand GNAME13615(G13615,G8788,G59758);
  nand GNAME13616(G13616,G8783,G13970,G13971);
  or GNAME13617(G13617,G9951,G8823);
  nand GNAME13618(G13618,G9883,G8791);
  nand GNAME13619(G13619,G9764,G9240,G13972,G13973);
  nand GNAME13620(G13620,G13619,G59428);
  nand GNAME13621(G13621,G8801,G9238);
  nand GNAME13622(G13622,G59428,G8896);
  nand GNAME13623(G13623,G9809,G13621,G13622,G9242);
  nand GNAME13624(G13624,G10221,G9953);
  nand GNAME13625(G13625,G13624,G59735);
  nand GNAME13626(G13626,G13623,G59576);
  nand GNAME13627(G13627,G59703,G9244);
  nand GNAME13628(G13628,G8833,G59608);
  nand GNAME13629(G13629,G8856,G22924);
  nand GNAME13630(G13630,G13624,G59734);
  nand GNAME13631(G13631,G13623,G59575);
  nand GNAME13632(G13632,G59702,G9244);
  nand GNAME13633(G13633,G8833,G59607);
  nand GNAME13634(G13634,G8856,G22925);
  nand GNAME13635(G13635,G13624,G59733);
  nand GNAME13636(G13636,G13623,G59574);
  nand GNAME13637(G13637,G59701,G9244);
  nand GNAME13638(G13638,G8833,G59606);
  nand GNAME13639(G13639,G8856,G22926);
  nand GNAME13640(G13640,G13624,G59732);
  nand GNAME13641(G13641,G13623,G59573);
  nand GNAME13642(G13642,G59700,G9244);
  nand GNAME13643(G13643,G8833,G59605);
  nand GNAME13644(G13644,G8856,G22927);
  nand GNAME13645(G13645,G13624,G59731);
  nand GNAME13646(G13646,G13623,G59572);
  nand GNAME13647(G13647,G59699,G9244);
  nand GNAME13648(G13648,G8833,G59604);
  nand GNAME13649(G13649,G8856,G22928);
  nand GNAME13650(G13650,G13624,G59730);
  nand GNAME13651(G13651,G13623,G59571);
  nand GNAME13652(G13652,G59698,G9244);
  nand GNAME13653(G13653,G8833,G59603);
  nand GNAME13654(G13654,G8856,G22929);
  nand GNAME13655(G13655,G13624,G59757);
  nand GNAME13656(G13656,G13623,G59598);
  nand GNAME13657(G13657,G59725,G9244);
  nand GNAME13658(G13658,G8833,G59630);
  nand GNAME13659(G13659,G13624,G59756);
  nand GNAME13660(G13660,G13623,G59597);
  nand GNAME13661(G13661,G59724,G9244);
  nand GNAME13662(G13662,G8833,G59629);
  nand GNAME13663(G13663,G8856,G22932);
  nand GNAME13664(G13664,G21598,G9238);
  nand GNAME13665(G13665,G9241,G9991,G13664);
  nand GNAME13666(G13666,G13665,G59558);
  nand GNAME13667(G13667,G13624,G59729);
  nand GNAME13668(G13668,G13623,G59570);
  nand GNAME13669(G13669,G59697,G9244);
  nand GNAME13670(G13670,G8833,G59602);
  nand GNAME13671(G13671,G8856,G22930);
  nand GNAME13672(G13672,G8813,G13879);
  nand GNAME13673(G13673,G8941,G8940);
  nand GNAME13674(G13674,G8802,G59563);
  nand GNAME13675(G13675,G13624,G59755);
  nand GNAME13676(G13676,G13623,G59596);
  nand GNAME13677(G13677,G59723,G9244);
  nand GNAME13678(G13678,G8833,G59628);
  nand GNAME13679(G13679,G8856,G22883);
  nand GNAME13680(G13680,G13624,G59754);
  nand GNAME13681(G13681,G13623,G59595);
  nand GNAME13682(G13682,G59722,G9244);
  nand GNAME13683(G13683,G8833,G59627);
  nand GNAME13684(G13684,G8856,G22882);
  nand GNAME13685(G13685,G13624,G59753);
  nand GNAME13686(G13686,G13623,G59594);
  nand GNAME13687(G13687,G59721,G9244);
  nand GNAME13688(G13688,G8833,G59626);
  nand GNAME13689(G13689,G8856,G22934);
  nand GNAME13690(G13690,G13624,G59752);
  nand GNAME13691(G13691,G13623,G59593);
  nand GNAME13692(G13692,G59720,G9244);
  nand GNAME13693(G13693,G8833,G59625);
  nand GNAME13694(G13694,G8856,G22881);
  nand GNAME13695(G13695,G13624,G59751);
  nand GNAME13696(G13696,G13623,G59592);
  nand GNAME13697(G13697,G59719,G9244);
  nand GNAME13698(G13698,G8833,G59624);
  nand GNAME13699(G13699,G8856,G22880);
  nand GNAME13700(G13700,G13624,G59750);
  nand GNAME13701(G13701,G13623,G59591);
  nand GNAME13702(G13702,G59718,G9244);
  nand GNAME13703(G13703,G8833,G59623);
  nand GNAME13704(G13704,G8856,G22958);
  nand GNAME13705(G13705,G13624,G59749);
  nand GNAME13706(G13706,G13623,G59590);
  nand GNAME13707(G13707,G59717,G9244);
  nand GNAME13708(G13708,G8833,G59622);
  nand GNAME13709(G13709,G8856,G22959);
  nand GNAME13710(G13710,G13624,G59748);
  nand GNAME13711(G13711,G13623,G59589);
  nand GNAME13712(G13712,G59716,G9244);
  nand GNAME13713(G13713,G8833,G59621);
  nand GNAME13714(G13714,G8856,G22960);
  nand GNAME13715(G13715,G13624,G59747);
  nand GNAME13716(G13716,G13623,G59588);
  nand GNAME13717(G13717,G59715,G9244);
  nand GNAME13718(G13718,G8833,G59620);
  nand GNAME13719(G13719,G8856,G22961);
  nand GNAME13720(G13720,G13624,G59746);
  nand GNAME13721(G13721,G13623,G59587);
  nand GNAME13722(G13722,G59714,G9244);
  nand GNAME13723(G13723,G8833,G59619);
  nand GNAME13724(G13724,G8856,G22962);
  nand GNAME13725(G13725,G13665,G59559);
  nand GNAME13726(G13726,G13624,G59728);
  nand GNAME13727(G13727,G13623,G59569);
  nand GNAME13728(G13728,G59696,G9244);
  nand GNAME13729(G13729,G8833,G59601);
  nand GNAME13730(G13730,G8856,G22933);
  nand GNAME13731(G13731,G13892,G8940);
  nand GNAME13732(G13732,G8813,G11066);
  nand GNAME13733(G13733,G8802,G59564);
  nand GNAME13734(G13734,G13624,G59745);
  nand GNAME13735(G13735,G13623,G59586);
  nand GNAME13736(G13736,G59713,G9244);
  nand GNAME13737(G13737,G8833,G59618);
  nand GNAME13738(G13738,G8856,G22964);
  nand GNAME13739(G13739,G13624,G59744);
  nand GNAME13740(G13740,G13623,G59585);
  nand GNAME13741(G13741,G59712,G9244);
  nand GNAME13742(G13742,G8833,G59617);
  nand GNAME13743(G13743,G8856,G22965);
  nand GNAME13744(G13744,G13624,G59743);
  nand GNAME13745(G13745,G13623,G59584);
  nand GNAME13746(G13746,G59711,G9244);
  nand GNAME13747(G13747,G8833,G59616);
  nand GNAME13748(G13748,G8856,G22966);
  nand GNAME13749(G13749,G13624,G59742);
  nand GNAME13750(G13750,G13623,G59583);
  nand GNAME13751(G13751,G59710,G9244);
  nand GNAME13752(G13752,G8833,G59615);
  nand GNAME13753(G13753,G8856,G22936);
  nand GNAME13754(G13754,G13624,G59741);
  nand GNAME13755(G13755,G13623,G59582);
  nand GNAME13756(G13756,G59709,G9244);
  nand GNAME13757(G13757,G8833,G59614);
  nand GNAME13758(G13758,G8856,G22937);
  nand GNAME13759(G13759,G13624,G59740);
  nand GNAME13760(G13760,G13623,G59581);
  nand GNAME13761(G13761,G59708,G9244);
  nand GNAME13762(G13762,G8833,G59613);
  nand GNAME13763(G13763,G8856,G22938);
  nand GNAME13764(G13764,G13624,G59739);
  nand GNAME13765(G13765,G13623,G59580);
  nand GNAME13766(G13766,G59707,G9244);
  nand GNAME13767(G13767,G8833,G59612);
  nand GNAME13768(G13768,G8856,G22939);
  nand GNAME13769(G13769,G13624,G59738);
  nand GNAME13770(G13770,G13623,G59579);
  nand GNAME13771(G13771,G59706,G9244);
  nand GNAME13772(G13772,G8833,G59611);
  nand GNAME13773(G13773,G8856,G22940);
  nand GNAME13774(G13774,G13624,G59737);
  nand GNAME13775(G13775,G13623,G59578);
  nand GNAME13776(G13776,G59705,G9244);
  nand GNAME13777(G13777,G8833,G59610);
  nand GNAME13778(G13778,G8856,G22941);
  nand GNAME13779(G13779,G13624,G59736);
  nand GNAME13780(G13780,G13623,G59577);
  nand GNAME13781(G13781,G59704,G9244);
  nand GNAME13782(G13782,G8833,G59609);
  nand GNAME13783(G13783,G8856,G22942);
  nand GNAME13784(G13784,G13665,G59560);
  nand GNAME13785(G13785,G13624,G59727);
  nand GNAME13786(G13786,G13623,G59568);
  nand GNAME13787(G13787,G59695,G9244);
  nand GNAME13788(G13788,G8833,G59600);
  nand GNAME13789(G13789,G8856,G22935);
  nand GNAME13790(G13790,G9250,G8813);
  nand GNAME13791(G13791,G13886,G8940);
  nand GNAME13792(G13792,G8802,G59565);
  nand GNAME13793(G13793,G13665,G59561);
  nand GNAME13794(G13794,G13624,G59726);
  nand GNAME13795(G13795,G13623,G59567);
  nand GNAME13796(G13796,G59694,G9244);
  nand GNAME13797(G13797,G8833,G59599);
  nand GNAME13798(G13798,G8856,G22943);
  nand GNAME13799(G13799,G11096,G8940);
  nand GNAME13800(G13800,G8813,G11044);
  nand GNAME13801(G13801,G8802,G59566);
  not GNAME13802(G13802,G9245);
  or GNAME13803(G13803,G8834,G13982);
  nand GNAME13804(G13804,G13211,G13802);
  nand GNAME13805(G13805,G13267,G13802);
  nand GNAME13806(G13806,G59558,G59425);
  nand GNAME13807(G13807,G8780,G9917);
  nand GNAME13808(G13808,G13807,G9790);
  nand GNAME13809(G13809,G13808,G9108);
  nand GNAME13810(G13810,G13323,G13802);
  nand GNAME13811(G13811,G59559,G59425);
  nand GNAME13812(G13812,G8780,G13974,G13975);
  nand GNAME13813(G13813,G13379,G13802);
  nand GNAME13814(G13814,G13435,G13802);
  nand GNAME13815(G13815,G9790,G9246);
  nand GNAME13816(G13816,G22294,G9247);
  nand GNAME13817(G13817,G59427,G8115);
  nand GNAME13818(G13818,G9247,G22308);
  nand GNAME13819(G13819,G59427,G22878);
  nand GNAME13820(G13820,G9247,G22309);
  nand GNAME13821(G13821,G59427,G22879);
  nand GNAME13822(G13822,G9247,G22310);
  nand GNAME13823(G13823,G59427,G22876);
  nand GNAME13824(G13824,G9247,G22307);
  nand GNAME13825(G13825,G59427,G22877);
  nand GNAME13826(G13826,G9247,G22295);
  nand GNAME13827(G13827,G8782,G9246);
  nand GNAME13828(G13828,G8834,G13827);
  nand GNAME13829(G13829,G59391,G12209,G12210);
  nand GNAME13830(G13830,G59798,G9110,G59392);
  nand GNAME13831(G13831,G59391,G1588,G12214);
  nand GNAME13832(G13832,G8782,G9183);
  nand GNAME13833(G13833,G13981,G59804);
  nand GNAME13834(G13834,G9769,G9958);
  nand GNAME13835(G13835,G59803,G13981);
  nand GNAME13836(G13836,G9769,G9959);
  nand GNAME13837(G13837,G9784,G59800);
  nand GNAME13838(G13838,G8811,G59804);
  or GNAME13839(G13839,G59801,G9784);
  nand GNAME13840(G13840,G9784,G59799);
  nand GNAME13841(G13841,G59798,G9770);
  or GNAME13842(G13842,G9770,G9987);
  nand GNAME13843(G13843,G8807,G35);
  nand GNAME13844(G13844,G9961,G59797);
  nand GNAME13845(G13845,G8781,G9849);
  nand GNAME13846(G13846,G8796,G9883);
  not GNAME13847(G13847,G9249);
  nand GNAME13848(G13848,G9784,G59794);
  or GNAME13849(G13849,G59803,G9784);
  nand GNAME13850(G13850,G13985,G59793);
  nand GNAME13851(G13851,G8829,G59758);
  nand GNAME13852(G13852,G8780,G8783,G8782);
  nand GNAME13853(G13853,G9832,G8783,G8746);
  nand GNAME13854(G13854,G8783,G8894);
  nand GNAME13855(G13855,G10841,G9900);
  nand GNAME13856(G13856,G8792,G10833,G9951);
  nand GNAME13857(G13857,G8745,G9866);
  nand GNAME13858(G13858,G8814,G8813);
  nand GNAME13859(G13859,G59427,G8751,G8787);
  nand GNAME13860(G13860,G8917,G59428,G21598);
  nand GNAME13861(G13861,G59566,G11040);
  nand GNAME13862(G13862,G8838,G59567);
  nand GNAME13863(G13863,G9282,G59567);
  nand GNAME13864(G13864,G13862,G13863);
  or GNAME13865(G13865,G59566,G59426);
  nand GNAME13866(G13866,G8813,G59566);
  or GNAME13867(G13867,G9282,G59568);
  or GNAME13868(G13868,G8838,G23082);
  nand GNAME13869(G13869,G8920,G9801);
  nand GNAME13870(G13870,G8919,G11051);
  nand GNAME13871(G13871,G11055,G9399);
  or GNAME13872(G13872,G11055,G9399);
  not GNAME13873(G13873,G9250);
  or GNAME13874(G13874,G8923,G8922);
  nand GNAME13875(G13875,G8922,G8923);
  not GNAME13876(G13876,G9251);
  or GNAME13877(G13877,G9773,G9772);
  nand GNAME13878(G13878,G9772,G9773);
  not GNAME13879(G13879,G9252);
  or GNAME13880(G13880,G8752,G9774);
  nand GNAME13881(G13881,G9774,G11116);
  or GNAME13882(G13882,G11094,G9775);
  nand GNAME13883(G13883,G9775,G11094);
  nand GNAME13884(G13884,G11119,G9400);
  or GNAME13885(G13885,G11119,G9400);
  not GNAME13886(G13886,G9253);
  or GNAME13887(G13887,G8756,G9774);
  nand GNAME13888(G13888,G9774,G11134);
  nand GNAME13889(G13889,G11160,G11163);
  nand GNAME13890(G13890,G8936,G13889);
  nand GNAME13891(G13891,G11138,G11160,G11163);
  not GNAME13892(G13892,G9264);
  nand GNAME13893(G13893,G8792,G59559);
  nand GNAME13894(G13894,G8761,G9866);
  not GNAME13895(G13895,G9255);
  nand GNAME13896(G13896,G11144,G59559);
  nand GNAME13897(G13897,G8761,G9776);
  not GNAME13898(G13898,G9254);
  or GNAME13899(G13899,G8761,G9774);
  nand GNAME13900(G13900,G9774,G11155);
  or GNAME13901(G13901,G8768,G9777);
  nand GNAME13902(G13902,G9777,G11170);
  or GNAME13903(G13903,G8768,G9774);
  nand GNAME13904(G13904,G9774,G11182);
  nand GNAME13905(G13905,G9774,G8862,G8790,G22013);
  or GNAME13906(G13906,G13982,G9774);
  nand GNAME13907(G13907,G12187,G59428);
  nand GNAME13908(G13908,G8787,G12188);
  or GNAME13909(G13909,G8787,G9107);
  nand GNAME13910(G13910,G9107,G12194);
  nand GNAME13911(G13911,G9961,G59394);
  nand GNAME13912(G13912,G8807,G12204);
  nand GNAME13913(G13913,G8807,G9771,G12203);
  nand GNAME13914(G13914,G9961,G59393);
  nand GNAME13915(G13915,G8804,G12207);
  nand GNAME13916(G13916,G59391,G12205,G59392);
  or GNAME13917(G13917,G8806,G8748,G59391,G59798);
  nand GNAME13918(G13918,G8806,G9109,G59390);
  nand GNAME13919(G13919,G9784,G59359);
  nand GNAME13920(G13920,G8811,G59793);
  nand GNAME13921(G13921,G9784,G59358);
  nand GNAME13922(G13922,G8811,G59792);
  nand GNAME13923(G13923,G9784,G59357);
  nand GNAME13924(G13924,G8811,G59791);
  nand GNAME13925(G13925,G9784,G59356);
  nand GNAME13926(G13926,G8811,G59790);
  nand GNAME13927(G13927,G8761,G59560);
  nand GNAME13928(G13928,G8756,G59559);
  not GNAME13929(G13929,G9256);
  nand GNAME13930(G13930,G8756,G59558);
  nand GNAME13931(G13931,G59560,G8762);
  or GNAME13932(G13932,G59795,G8761);
  nand GNAME13933(G13933,G59795,G13864,G11066);
  or GNAME13934(G13934,G59795,G8756);
  nand GNAME13935(G13935,G59795,G13864,G9250);
  or GNAME13936(G13936,G59795,G8752);
  nand GNAME13937(G13937,G11112,G59795);
  nand GNAME13938(G13938,G9778,G22013,G8862);
  or GNAME13939(G13939,G13982,G9778);
  or GNAME13940(G13940,G8768,G9778);
  nand GNAME13941(G13941,G9778,G11179);
  or GNAME13942(G13942,G8761,G9778);
  nand GNAME13943(G13943,G9778,G11151);
  or GNAME13944(G13944,G8756,G9778);
  nand GNAME13945(G13945,G9778,G11130);
  or GNAME13946(G13946,G8752,G9778);
  nand GNAME13947(G13947,G9778,G11111);
  nand GNAME13948(G13948,G8814,G59757);
  nand GNAME13949(G13949,G59427,G59598);
  nand GNAME13950(G13950,G9866,G59597);
  nand GNAME13951(G13951,G8792,G12715);
  nand GNAME13952(G13952,G9866,G59596);
  nand GNAME13953(G13953,G8792,G12732);
  nand GNAME13954(G13954,G9866,G59595);
  nand GNAME13955(G13955,G8792,G12749);
  nand GNAME13956(G13956,G9866,G59594);
  nand GNAME13957(G13957,G8792,G12766);
  nand GNAME13958(G13958,G9866,G59593);
  nand GNAME13959(G13959,G8792,G12783);
  nand GNAME13960(G13960,G9866,G59592);
  nand GNAME13961(G13961,G8792,G12800);
  nand GNAME13962(G13962,G9866,G59591);
  nand GNAME13963(G13963,G8792,G12817);
  nand GNAME13964(G13964,G9866,G59590);
  nand GNAME13965(G13965,G8792,G12834);
  nand GNAME13966(G13966,G9951,G9917);
  nand GNAME13967(G13967,G8746,G8860);
  nand GNAME13968(G13968,G8792,G9951);
  nand GNAME13969(G13969,G8784,G9866);
  nand GNAME13970(G13970,G8782,G9832);
  nand GNAME13971(G13971,G8780,G8746);
  nand GNAME13972(G13972,G8796,G8887);
  nand GNAME13973(G13973,G9849,G9934);
  nand GNAME13974(G13974,G8782,G9849);
  nand GNAME13975(G13975,G8796,G9951);
  nand GNAME13976(G13976,G59560,G59425);
  nand GNAME13977(G13977,G8834,G13812);
  nand GNAME13978(G13978,G59561,G59425);
  nand GNAME13979(G13979,G8834,G13808);
  not GNAME13980(G13980,G8803);
  not GNAME13981(G13981,G9769);
  not GNAME13982(G13982,G59557);
  not GNAME13983(G13983,G8944);
  not GNAME13984(G13984,G8908);
  not GNAME13985(G13985,G8829);
  not GNAME13986(G13986,G8794);
  not GNAME13987(G13987,G9185);
  nand GNAME13988(G13988,G8031,G8030);
  and GNAME13989(G13989,G15281,G13990);
  and GNAME13990(G13990,G13991,G15283,G15282);
  and GNAME13991(G13991,G15284,G13992);
  and GNAME13992(G13992,G15285,G8082,G15286);
  not GNAME13993(G13993,G14300);
  and GNAME13994(G13994,G8043,G8042);
  not GNAME13995(G13995,G14301);
  and GNAME13996(G13996,G8046,G8045);
  not GNAME13997(G13997,G14302);
  and GNAME13998(G13998,G8049,G8048);
  not GNAME13999(G13999,G14303);
  and GNAME14000(G14000,G8052,G8051);
  not GNAME14001(G14001,G14304);
  and GNAME14002(G14002,G8055,G8054);
  not GNAME14003(G14003,G14305);
  and GNAME14004(G14004,G8058,G8057);
  not GNAME14005(G14005,G14306);
  and GNAME14006(G14006,G8061,G8060);
  not GNAME14007(G14007,G14283);
  and GNAME14008(G14008,G14284,G14285,G14010);
  not GNAME14009(G14009,G14284);
  and GNAME14010(G14010,G14286,G14287,G14012);
  not GNAME14011(G14011,G14286);
  and GNAME14012(G14012,G14288,G8063,G14289);
  not GNAME14013(G14013,G14288);
  not GNAME14014(G14014,G14289);
  nand GNAME14015(G14015,G14017,G14290);
  not GNAME14016(G14016,G14290);
  and GNAME14017(G14017,G14292,G14020,G14291);
  not GNAME14018(G14018,G14292);
  not GNAME14019(G14019,G14291);
  and GNAME14020(G14020,G14293,G14021);
  and GNAME14021(G14021,G14294,G14024,G14295);
  not GNAME14022(G14022,G14294);
  not GNAME14023(G14023,G14295);
  and GNAME14024(G14024,G8064,G14296);
  not GNAME14025(G14025,G14296);
  not GNAME14026(G14026,G14299);
  not GNAME14027(G14027,G14298);
  nand GNAME14028(G14028,G8065,G15863);
  and GNAME14029(G14029,G2085,G8038);
  nor GNAME14030(G14030,G13990,G8036);
  and GNAME14031(G14031,G8066,G8035);
  nor GNAME14032(G14032,G13992,G8033);
  not GNAME14033(G14033,G15271);
  not GNAME14034(G14034,G14113);
  not GNAME14035(G14035,G15273);
  not GNAME14036(G14036,G15272);
  not GNAME14037(G14037,G20036);
  not GNAME14038(G14038,G20042);
  not GNAME14039(G14039,G20046);
  not GNAME14040(G14040,G19993);
  or GNAME14041(G14041,G20061,G20009);
  nand GNAME14042(G14042,G20061,G20009);
  or GNAME14043(G14043,G23424,G20060);
  nand GNAME14044(G14044,G20060,G23424);
  or GNAME14045(G14045,G20059,G20010);
  nand GNAME14046(G14046,G20059,G20010);
  or GNAME14047(G14047,G23484,G20058);
  nand GNAME14048(G14048,G20058,G23484);
  or GNAME14049(G14049,G20057,G20011);
  nand GNAME14050(G14050,G20057,G20011);
  or GNAME14051(G14051,G23483,G20056);
  nand GNAME14052(G14052,G20056,G23483);
  or GNAME14053(G14053,G20055,G20012);
  nand GNAME14054(G14054,G20055,G20012);
  or GNAME14055(G14055,G23482,G20054);
  nand GNAME14056(G14056,G20054,G23482);
  or GNAME14057(G14057,G20052,G20013);
  nand GNAME14058(G14058,G20052,G20013);
  or GNAME14059(G14059,G23425,G20053);
  or GNAME14060(G14060,G14123,G20001);
  or GNAME14061(G14061,G23480,G19995);
  or GNAME14062(G14062,G20003,G20050);
  nand GNAME14063(G14063,G20047,G20049);
  or GNAME14064(G14064,G20049,G20047);
  nand GNAME14065(G14065,G20048,G20004);
  or GNAME14066(G14066,G20004,G20048);
  nand GNAME14067(G14067,G20046,G23535);
  or GNAME14068(G14068,G23535,G20046);
  nand GNAME14069(G14069,G20043,G20045);
  or GNAME14070(G14070,G20045,G20043);
  nand GNAME14071(G14071,G20044,G20005);
  or GNAME14072(G14072,G20005,G20044);
  nand GNAME14073(G14073,G20042,G23523);
  or GNAME14074(G14074,G23523,G20042);
  nand GNAME14075(G14075,G20039,G20041);
  or GNAME14076(G14076,G20041,G20039);
  nand GNAME14077(G14077,G20040,G20006);
  or GNAME14078(G14078,G20006,G20040);
  nand GNAME14079(G14079,G20037,G23479);
  or GNAME14080(G14080,G23479,G20037);
  nand GNAME14081(G14081,G20038,G20007);
  or GNAME14082(G14082,G20007,G20038);
  nand GNAME14083(G14083,G20036,G23477);
  or GNAME14084(G14084,G23477,G20036);
  nand GNAME14085(G14085,G20034,G20035);
  or GNAME14086(G14086,G20035,G20034);
  nand GNAME14087(G14087,G20032,G20033);
  or GNAME14088(G14088,G20033,G20032);
  or GNAME14089(G14089,G23427,G20008);
  nand GNAME14090(G14090,G20008,G23427);
  nand GNAME14091(G14091,G20064,G14129);
  or GNAME14092(G14092,G14129,G20064);
  or GNAME14093(G14093,G20062,G20014);
  nand GNAME14094(G14094,G20062,G20014);
  or GNAME14095(G14095,G23461,G20063);
  nand GNAME14096(G14096,G20063,G23461);
  nand GNAME14097(G14097,G19993,G20031);
  or GNAME14098(G14098,G14099,G20051);
  and GNAME14099(G14099,G19993,G14100);
  or GNAME14100(G14100,G14122,G23481);
  or GNAME14101(G14101,G14123,G14104);
  nand GNAME14102(G14102,G20001,G14103);
  or GNAME14103(G14103,G20052,G20053);
  not GNAME14104(G14104,G20052);
  or GNAME14105(G14105,G20055,G20054);
  nand GNAME14106(G14106,G14107,G23482);
  nand GNAME14107(G14107,G20054,G20055);
  or GNAME14108(G14108,G20057,G20056);
  nand GNAME14109(G14109,G14110,G23483);
  nand GNAME14110(G14110,G20056,G20057);
  or GNAME14111(G14111,G20059,G20058);
  nor GNAME14112(G14112,G60244,G19979);
  nor GNAME14113(G14113,G60244,G14765);
  nand GNAME14114(G14114,G15530,G15531,G15532,G15533);
  nand GNAME14115(G14115,G15534,G15535,G15536,G15537);
  nand GNAME14116(G14116,G15538,G15539,G15540,G15541);
  nand GNAME14117(G14117,G15542,G15543,G15544,G15545);
  nand GNAME14118(G14118,G15546,G15547,G15548,G15549);
  nand GNAME14119(G14119,G15550,G15551,G15552,G15553);
  nand GNAME14120(G14120,G15554,G15555,G15556,G15557);
  nand GNAME14121(G14121,G15558,G15559,G15560,G15561);
  nand GNAME14122(G14122,G15562,G15563,G15564,G15565);
  nand GNAME14123(G14123,G15566,G15567,G15568,G15569);
  nand GNAME14124(G14124,G15570,G15571,G15572,G15573);
  nand GNAME14125(G14125,G15574,G15575,G15576,G15577);
  nand GNAME14126(G14126,G15578,G15579,G15580,G15581);
  nand GNAME14127(G14127,G15582,G15583,G15584,G15585);
  nand GNAME14128(G14128,G15586,G15587,G15588,G15589);
  nand GNAME14129(G14129,G15590,G15591,G15592,G15593);
  nand GNAME14130(G14130,G19825,G14811);
  nand GNAME14131(G14131,G19813,G19814);
  or GNAME14132(G14132,G14131,G19799);
  nand GNAME14133(G14133,G19815,G15242,G19814);
  nand GNAME14134(G14134,G15245,G19816,G19817);
  nand GNAME14135(G14135,G15245,G19818,G19819);
  nand GNAME14136(G14136,G15245,G19820,G19821);
  nand GNAME14137(G14137,G15245,G19822,G19823);
  and GNAME14138(G14138,G19009,G19799);
  and GNAME14139(G14139,G19064,G19799);
  and GNAME14140(G14140,G19119,G19799);
  nand GNAME14141(G14141,G19800,G19801);
  nand GNAME14142(G14142,G19802,G19803);
  nand GNAME14143(G14143,G19808,G19806,G19807);
  nand GNAME14144(G14144,G19973,G19974,G14811,G19810);
  nand GNAME14145(G14145,G19975,G19976,G14811,G19811);
  nand GNAME14146(G14146,G19652,G19653,G19654,G19655);
  nand GNAME14147(G14147,G19659,G19660,G19658,G19656,G19657);
  nand GNAME14148(G14148,G19675,G19676,G19674,G19672,G19673);
  nand GNAME14149(G14149,G19680,G19681,G19679,G19677,G19678);
  nand GNAME14150(G14150,G19685,G19686,G19684,G19682,G19683);
  nand GNAME14151(G14151,G19690,G19691,G19689,G19687,G19688);
  nand GNAME14152(G14152,G19695,G19696,G19694,G19692,G19693);
  nand GNAME14153(G14153,G19700,G19701,G19699,G19697,G19698);
  nand GNAME14154(G14154,G19705,G19706,G19704,G19702,G19703);
  nand GNAME14155(G14155,G19710,G19711,G19709,G19707,G19708);
  nand GNAME14156(G14156,G19715,G19716,G19714,G19712,G19713);
  nand GNAME14157(G14157,G19720,G19721,G19719,G19717,G19718);
  nand GNAME14158(G14158,G19734,G19735,G19733,G19731,G19732);
  nand GNAME14159(G14159,G19739,G19740,G19738,G19736,G19737);
  nand GNAME14160(G14160,G19744,G19745,G19743,G19741,G19742);
  nand GNAME14161(G14161,G19749,G19750,G19748,G19746,G19747);
  nand GNAME14162(G14162,G19754,G19755,G19753,G19751,G19752);
  nand GNAME14163(G14163,G19759,G19760,G19758,G19756,G19757);
  nand GNAME14164(G14164,G19764,G19765,G19763,G19761,G19762);
  nand GNAME14165(G14165,G19769,G19770,G19768,G19766,G19767);
  nand GNAME14166(G14166,G19774,G19775,G19773,G19771,G19772);
  nand GNAME14167(G14167,G19779,G19780,G19778,G19776,G19777);
  nand GNAME14168(G14168,G19625,G19626,G19624,G19622,G19623);
  nand GNAME14169(G14169,G19630,G19631,G19629,G19627,G19628);
  nand GNAME14170(G14170,G19635,G19636,G19634,G19632,G19633);
  nand GNAME14171(G14171,G19640,G19641,G19639,G19637,G19638);
  nand GNAME14172(G14172,G19645,G19646,G19644,G19642,G19643);
  nand GNAME14173(G14173,G19650,G19651,G19649,G19647,G19648);
  nand GNAME14174(G14174,G15762,G19663,G19669,G19670,G19665);
  nand GNAME14175(G14175,G15763,G19722,G19728,G19729,G19724);
  nand GNAME14176(G14176,G15764,G19781,G19787,G19788,G19783);
  nand GNAME14177(G14177,G15765,G19790,G19796,G19797,G19792);
  and GNAME14178(G14178,G14122,G14853);
  and GNAME14179(G14179,G14123,G14853);
  and GNAME14180(G14180,G14124,G14853);
  and GNAME14181(G14181,G14125,G14853);
  and GNAME14182(G14182,G14126,G14853);
  and GNAME14183(G14183,G14127,G14853);
  and GNAME14184(G14184,G14128,G14853);
  and GNAME14185(G14185,G14129,G14853);
  nand GNAME14186(G14186,G14869,G15236,G15988,G15793,G15806);
  nand GNAME14187(G14187,G15794,G15988,G19617,G15240);
  nand GNAME14188(G14188,G19492,G19493,G19494,G19495);
  nand GNAME14189(G14189,G19499,G19500,G19498,G19496,G19497);
  nand GNAME14190(G14190,G19514,G19515,G19513,G19511,G19512);
  nand GNAME14191(G14191,G19519,G19520,G19518,G19516,G19517);
  nand GNAME14192(G14192,G19524,G19525,G19523,G19521,G19522);
  nand GNAME14193(G14193,G19529,G19530,G19528,G19526,G19527);
  nand GNAME14194(G14194,G19534,G19535,G19533,G19531,G19532);
  nand GNAME14195(G14195,G19539,G19540,G19538,G19536,G19537);
  nand GNAME14196(G14196,G19544,G19545,G19543,G19541,G19542);
  nand GNAME14197(G14197,G19546,G19547,G19548,G19549);
  nand GNAME14198(G14198,G19550,G19551,G19552,G19553);
  nand GNAME14199(G14199,G19554,G19555,G19556,G19557);
  nand GNAME14200(G14200,G19563,G19564,G19565,G19566);
  nand GNAME14201(G14201,G19567,G19568,G19569,G19570);
  nand GNAME14202(G14202,G19571,G19572,G19573,G19574);
  nand GNAME14203(G14203,G19575,G19576,G19577,G19578);
  nand GNAME14204(G14204,G19579,G19580,G19581,G19582);
  nand GNAME14205(G14205,G19583,G19584,G19585,G19586);
  nand GNAME14206(G14206,G19587,G19588,G19589,G19590);
  nand GNAME14207(G14207,G19591,G19592,G19593,G19594);
  nand GNAME14208(G14208,G19595,G19596,G19597,G19598);
  nand GNAME14209(G14209,G19599,G19600,G19601,G19602);
  nand GNAME14210(G14210,G19465,G19466,G19467,G19468);
  nand GNAME14211(G14211,G19469,G19470,G19471,G19472);
  nand GNAME14212(G14212,G19473,G19474,G19475,G19476);
  nand GNAME14213(G14213,G19477,G19478,G19479,G19480);
  nand GNAME14214(G14214,G19481,G19482,G19483,G19484);
  nand GNAME14215(G14215,G19490,G19491,G19489,G19487,G19488);
  nand GNAME14216(G14216,G19509,G19510,G19508,G19506,G19507);
  nand GNAME14217(G14217,G19561,G19562,G19560,G19558,G19559);
  nand GNAME14218(G14218,G19606,G19607,G19605,G19603,G19604);
  nand GNAME14219(G14219,G19611,G19612,G19610,G19608,G19609);
  and GNAME14220(G14220,G19026,G14861);
  and GNAME14221(G14221,G19081,G14861);
  and GNAME14222(G14222,G19136,G14861);
  and GNAME14223(G14223,G19174,G14861);
  and GNAME14224(G14224,G19230,G14861);
  and GNAME14225(G14225,G19286,G14861);
  and GNAME14226(G14226,G19342,G14861);
  and GNAME14227(G14227,G19398,G14861);
  and GNAME14228(G14228,G59998,G14853);
  and GNAME14229(G14229,G59999,G14853);
  and GNAME14230(G14230,G60000,G14853);
  and GNAME14231(G14231,G60001,G14853);
  and GNAME14232(G14232,G60002,G14853);
  nand GNAME14233(G14233,G19439,G15792,G19438);
  nand GNAME14234(G14234,G15236,G15758,G15950,G15796,G15804);
  nand GNAME14235(G14235,G15794,G19438,G19446,G19447);
  nand GNAME14236(G14236,G19044,G19045,G19046,G19047);
  nand GNAME14237(G14237,G19099,G19100,G19101,G19102);
  nand GNAME14238(G14238,G19154,G19155,G19156,G19157);
  nand GNAME14239(G14239,G19212,G19213,G19211,G19209,G19210);
  nand GNAME14240(G14240,G19268,G19269,G19267,G19265,G19266);
  nand GNAME14241(G14241,G15731,G19322,G15788,G19321);
  nand GNAME14242(G14242,G15744,G15779,G15182,G19377,G19378);
  nand GNAME14243(G14243,G15757,G15788,G15802,G19433,G19434);
  nand GNAME14244(G14244,G18864,G18865,G18866,G18867);
  nand GNAME14245(G14245,G18871,G18872,G18870,G18868,G18869);
  nand GNAME14246(G14246,G18881,G18882,G18880,G18878,G18879);
  nand GNAME14247(G14247,G18886,G18887,G18885,G18883,G18884);
  nand GNAME14248(G14248,G18891,G18892,G18890,G18888,G18889);
  nand GNAME14249(G14249,G18896,G18897,G18895,G18893,G18894);
  nand GNAME14250(G14250,G18901,G18902,G18900,G18898,G18899);
  nand GNAME14251(G14251,G18906,G18907,G18905,G18903,G18904);
  nand GNAME14252(G14252,G18911,G18912,G18910,G18908,G18909);
  nand GNAME14253(G14253,G18916,G18917,G18915,G18913,G18914);
  nand GNAME14254(G14254,G18921,G18922,G18920,G18918,G18919);
  nand GNAME14255(G14255,G18926,G18927,G18925,G18923,G18924);
  nand GNAME14256(G14256,G18936,G18937,G18935,G18933,G18934);
  nand GNAME14257(G14257,G18941,G18942,G18940,G18938,G18939);
  nand GNAME14258(G14258,G18946,G18947,G18945,G18943,G18944);
  nand GNAME14259(G14259,G18951,G18952,G18950,G18948,G18949);
  nand GNAME14260(G14260,G18956,G18957,G18955,G18953,G18954);
  nand GNAME14261(G14261,G18961,G18962,G18960,G18958,G18959);
  nand GNAME14262(G14262,G18966,G18967,G18965,G18963,G18964);
  nand GNAME14263(G14263,G18971,G18972,G18970,G18968,G18969);
  nand GNAME14264(G14264,G18976,G18977,G18975,G18973,G18974);
  nand GNAME14265(G14265,G18981,G18982,G18980,G18978,G18979);
  nand GNAME14266(G14266,G18837,G18838,G18836,G18834,G18835);
  nand GNAME14267(G14267,G18842,G18843,G18841,G18839,G18840);
  nand GNAME14268(G14268,G18847,G18848,G18846,G18844,G18845);
  nand GNAME14269(G14269,G18852,G18853,G18851,G18849,G18850);
  nand GNAME14270(G14270,G18857,G18858,G18856,G18854,G18855);
  nand GNAME14271(G14271,G18862,G18863,G18861,G18859,G18860);
  nand GNAME14272(G14272,G18876,G18877,G18875,G18873,G18874);
  nand GNAME14273(G14273,G18931,G18932,G18930,G18928,G18929);
  nand GNAME14274(G14274,G18986,G18987,G18985,G18983,G18984);
  nand GNAME14275(G14275,G15658,G18990,G18988,G18989);
  and GNAME14276(G14276,G15863,G60047);
  and GNAME14277(G14277,G15863,G60038);
  and GNAME14278(G14278,G15863,G60037);
  and GNAME14279(G14279,G15863,G60036);
  and GNAME14280(G14280,G15863,G60035);
  and GNAME14281(G14281,G15863,G60034);
  and GNAME14282(G14282,G15863,G60033);
  and GNAME14283(G14283,G15863,G60032);
  and GNAME14284(G14284,G15863,G60031);
  and GNAME14285(G14285,G15863,G60030);
  and GNAME14286(G14286,G15863,G60029);
  and GNAME14287(G14287,G15863,G60028);
  and GNAME14288(G14288,G15863,G60027);
  and GNAME14289(G14289,G15863,G60026);
  and GNAME14290(G14290,G15863,G60025);
  and GNAME14291(G14291,G15863,G60024);
  and GNAME14292(G14292,G15863,G60023);
  and GNAME14293(G14293,G15863,G60022);
  and GNAME14294(G14294,G15863,G60021);
  and GNAME14295(G14295,G15863,G60020);
  and GNAME14296(G14296,G15863,G60019);
  and GNAME14297(G14297,G15863,G60018);
  and GNAME14298(G14298,G15863,G60017);
  and GNAME14299(G14299,G15863,G60016);
  and GNAME14300(G14300,G14789,G18576);
  and GNAME14301(G14301,G14789,G18593);
  and GNAME14302(G14302,G14789,G18610);
  and GNAME14303(G14303,G14789,G18627);
  and GNAME14304(G14304,G14789,G18644);
  and GNAME14305(G14305,G14789,G18661);
  and GNAME14306(G14306,G14789,G18678);
  and GNAME14307(G14307,G14789,G18695);
  nand GNAME14308(G14308,G18302,G18300,G18301);
  nand GNAME14309(G14309,G18299,G18297,G18298);
  nand GNAME14310(G14310,G18296,G18294,G18295);
  nand GNAME14311(G14311,G18293,G18291,G18292);
  nand GNAME14312(G14312,G18290,G18288,G18289);
  nand GNAME14313(G14313,G18287,G18285,G18286);
  nand GNAME14314(G14314,G18284,G18282,G18283);
  nand GNAME14315(G14315,G18281,G18279,G18280);
  nand GNAME14316(G14316,G18278,G18276,G18277);
  nand GNAME14317(G14317,G18275,G18273,G18274);
  nand GNAME14318(G14318,G18272,G18270,G18271);
  nand GNAME14319(G14319,G18269,G18267,G18268);
  nand GNAME14320(G14320,G18266,G18264,G18265);
  nand GNAME14321(G14321,G18263,G18261,G18262);
  nand GNAME14322(G14322,G18260,G18258,G18259);
  nand GNAME14323(G14323,G18257,G18255,G18256);
  nand GNAME14324(G14324,G18254,G18252,G18253);
  nand GNAME14325(G14325,G18251,G18249,G18250);
  nand GNAME14326(G14326,G18248,G18246,G18247);
  nand GNAME14327(G14327,G18245,G18243,G18244);
  nand GNAME14328(G14328,G18242,G18240,G18241);
  nand GNAME14329(G14329,G18239,G18237,G18238);
  nand GNAME14330(G14330,G18236,G18234,G18235);
  nand GNAME14331(G14331,G18233,G18231,G18232);
  nand GNAME14332(G14332,G18230,G18228,G18229);
  nand GNAME14333(G14333,G18227,G18225,G18226);
  nand GNAME14334(G14334,G18224,G18222,G18223);
  nand GNAME14335(G14335,G18221,G18219,G18220);
  nand GNAME14336(G14336,G18218,G18216,G18217);
  nand GNAME14337(G14337,G18215,G18213,G18214);
  nand GNAME14338(G14338,G15783,G18212,G19828,G19914,G19915);
  nand GNAME14339(G14339,G15782,G18208,G19826,G19827);
  nand GNAME14340(G14340,G19912,G19913,G18200,G18205);
  and GNAME14341(G14341,G15958,G59844);
  and GNAME14342(G14342,G15958,G59845);
  and GNAME14343(G14343,G15958,G59846);
  and GNAME14344(G14344,G15958,G59847);
  and GNAME14345(G14345,G15958,G59848);
  and GNAME14346(G14346,G15958,G59849);
  and GNAME14347(G14347,G15958,G59850);
  and GNAME14348(G14348,G15958,G59851);
  and GNAME14349(G14349,G15958,G59852);
  and GNAME14350(G14350,G15958,G59853);
  and GNAME14351(G14351,G15958,G59854);
  and GNAME14352(G14352,G15958,G59855);
  and GNAME14353(G14353,G15958,G59856);
  and GNAME14354(G14354,G15958,G59857);
  and GNAME14355(G14355,G15958,G59858);
  and GNAME14356(G14356,G15958,G59859);
  and GNAME14357(G14357,G15958,G59860);
  and GNAME14358(G14358,G15958,G59861);
  and GNAME14359(G14359,G15958,G59862);
  and GNAME14360(G14360,G15958,G59863);
  and GNAME14361(G14361,G15958,G59864);
  and GNAME14362(G14362,G15958,G59865);
  and GNAME14363(G14363,G15958,G59866);
  and GNAME14364(G14364,G15958,G59867);
  and GNAME14365(G14365,G15958,G59868);
  and GNAME14366(G14366,G15958,G59869);
  and GNAME14367(G14367,G15958,G59870);
  and GNAME14368(G14368,G15958,G59871);
  and GNAME14369(G14369,G15958,G59872);
  and GNAME14370(G14370,G15958,G59873);
  nand GNAME14371(G14371,G18199,G14906,G19981);
  nand GNAME14372(G14372,G15795,G15796,G18197,G18198);
  nand GNAME14373(G14373,G18196,G15808,G18195);
  nand GNAME14374(G14374,G19906,G19907,G15807,G15809);
  nand GNAME14375(G14375,G15528,G18176,G18174,G18175);
  nand GNAME14376(G14376,G15527,G18170,G18168,G18169);
  nand GNAME14377(G14377,G15526,G18164,G18162,G18163);
  nand GNAME14378(G14378,G15525,G18158,G18156,G18157);
  nand GNAME14379(G14379,G15524,G18152,G18150,G18151);
  nand GNAME14380(G14380,G15523,G18146,G18144,G18145);
  nand GNAME14381(G14381,G15522,G18140,G18138,G18139);
  nand GNAME14382(G14382,G15521,G18134,G18132,G18133);
  nand GNAME14383(G14383,G15520,G18115,G18113,G18114);
  nand GNAME14384(G14384,G15519,G18109,G18107,G18108);
  nand GNAME14385(G14385,G15518,G18103,G18101,G18102);
  nand GNAME14386(G14386,G15517,G18097,G18095,G18096);
  nand GNAME14387(G14387,G15516,G18091,G18089,G18090);
  nand GNAME14388(G14388,G15515,G18085,G18083,G18084);
  nand GNAME14389(G14389,G15514,G18079,G18077,G18078);
  nand GNAME14390(G14390,G15513,G18073,G18071,G18072);
  nand GNAME14391(G14391,G15512,G18054,G18052,G18053);
  nand GNAME14392(G14392,G15511,G18048,G18046,G18047);
  nand GNAME14393(G14393,G15510,G18042,G18040,G18041);
  nand GNAME14394(G14394,G15509,G18036,G18034,G18035);
  nand GNAME14395(G14395,G15508,G18030,G18028,G18029);
  nand GNAME14396(G14396,G15507,G18024,G18022,G18023);
  nand GNAME14397(G14397,G15506,G18018,G18016,G18017);
  nand GNAME14398(G14398,G15505,G18012,G18010,G18011);
  nand GNAME14399(G14399,G15504,G17993,G17991,G17992);
  nand GNAME14400(G14400,G15503,G17987,G17985,G17986);
  nand GNAME14401(G14401,G15502,G17981,G17979,G17980);
  nand GNAME14402(G14402,G15501,G17975,G17973,G17974);
  nand GNAME14403(G14403,G15500,G17969,G17967,G17968);
  nand GNAME14404(G14404,G15499,G17963,G17961,G17962);
  nand GNAME14405(G14405,G15498,G17957,G17955,G17956);
  nand GNAME14406(G14406,G15497,G17951,G17949,G17950);
  nand GNAME14407(G14407,G15496,G17932,G17930,G17931);
  nand GNAME14408(G14408,G15495,G17926,G17924,G17925);
  nand GNAME14409(G14409,G15494,G17920,G17918,G17919);
  nand GNAME14410(G14410,G15493,G17914,G17912,G17913);
  nand GNAME14411(G14411,G15492,G17908,G17906,G17907);
  nand GNAME14412(G14412,G15491,G17902,G17900,G17901);
  nand GNAME14413(G14413,G15490,G17896,G17894,G17895);
  nand GNAME14414(G14414,G15489,G17890,G17888,G17889);
  nand GNAME14415(G14415,G15488,G17871,G17869,G17870);
  nand GNAME14416(G14416,G15487,G17865,G17863,G17864);
  nand GNAME14417(G14417,G15486,G17859,G17857,G17858);
  nand GNAME14418(G14418,G15485,G17853,G17851,G17852);
  nand GNAME14419(G14419,G15484,G17847,G17845,G17846);
  nand GNAME14420(G14420,G15483,G17841,G17839,G17840);
  nand GNAME14421(G14421,G15482,G17835,G17833,G17834);
  nand GNAME14422(G14422,G15481,G17829,G17827,G17828);
  nand GNAME14423(G14423,G15480,G17810,G17808,G17809);
  nand GNAME14424(G14424,G15479,G17804,G17802,G17803);
  nand GNAME14425(G14425,G15478,G17798,G17796,G17797);
  nand GNAME14426(G14426,G15477,G17792,G17790,G17791);
  nand GNAME14427(G14427,G15476,G17786,G17784,G17785);
  nand GNAME14428(G14428,G15475,G17780,G17778,G17779);
  nand GNAME14429(G14429,G15474,G17774,G17772,G17773);
  nand GNAME14430(G14430,G15473,G17768,G17766,G17767);
  nand GNAME14431(G14431,G15472,G17749,G17747,G17748);
  nand GNAME14432(G14432,G15471,G17743,G17741,G17742);
  nand GNAME14433(G14433,G15470,G17737,G17735,G17736);
  nand GNAME14434(G14434,G15469,G17731,G17729,G17730);
  nand GNAME14435(G14435,G15468,G17725,G17723,G17724);
  nand GNAME14436(G14436,G15467,G17719,G17717,G17718);
  nand GNAME14437(G14437,G15466,G17713,G17711,G17712);
  nand GNAME14438(G14438,G15465,G17707,G17705,G17706);
  nand GNAME14439(G14439,G15464,G17688,G17686,G17687);
  nand GNAME14440(G14440,G15463,G17682,G17680,G17681);
  nand GNAME14441(G14441,G15462,G17676,G17674,G17675);
  nand GNAME14442(G14442,G15461,G17670,G17668,G17669);
  nand GNAME14443(G14443,G15460,G17664,G17662,G17663);
  nand GNAME14444(G14444,G15459,G17658,G17656,G17657);
  nand GNAME14445(G14445,G15458,G17652,G17650,G17651);
  nand GNAME14446(G14446,G15457,G17646,G17644,G17645);
  nand GNAME14447(G14447,G15456,G17627,G17625,G17626);
  nand GNAME14448(G14448,G15455,G17621,G17619,G17620);
  nand GNAME14449(G14449,G15454,G17615,G17613,G17614);
  nand GNAME14450(G14450,G15453,G17609,G17607,G17608);
  nand GNAME14451(G14451,G15452,G17603,G17601,G17602);
  nand GNAME14452(G14452,G15451,G17597,G17595,G17596);
  nand GNAME14453(G14453,G15450,G17591,G17589,G17590);
  nand GNAME14454(G14454,G15449,G17585,G17583,G17584);
  nand GNAME14455(G14455,G15448,G17566,G17564,G17565);
  nand GNAME14456(G14456,G15447,G17560,G17558,G17559);
  nand GNAME14457(G14457,G15446,G17554,G17552,G17553);
  nand GNAME14458(G14458,G15445,G17548,G17546,G17547);
  nand GNAME14459(G14459,G15444,G17542,G17540,G17541);
  nand GNAME14460(G14460,G15443,G17536,G17534,G17535);
  nand GNAME14461(G14461,G15442,G17530,G17528,G17529);
  nand GNAME14462(G14462,G15441,G17524,G17522,G17523);
  nand GNAME14463(G14463,G15440,G17505,G17503,G17504);
  nand GNAME14464(G14464,G15439,G17499,G17497,G17498);
  nand GNAME14465(G14465,G15438,G17493,G17491,G17492);
  nand GNAME14466(G14466,G15437,G17487,G17485,G17486);
  nand GNAME14467(G14467,G15436,G17481,G17479,G17480);
  nand GNAME14468(G14468,G15435,G17475,G17473,G17474);
  nand GNAME14469(G14469,G15434,G17469,G17467,G17468);
  nand GNAME14470(G14470,G15433,G17463,G17461,G17462);
  nand GNAME14471(G14471,G15432,G17444,G17442,G17443);
  nand GNAME14472(G14472,G15431,G17438,G17436,G17437);
  nand GNAME14473(G14473,G15430,G17432,G17430,G17431);
  nand GNAME14474(G14474,G15429,G17426,G17424,G17425);
  nand GNAME14475(G14475,G15428,G17420,G17418,G17419);
  nand GNAME14476(G14476,G15427,G17414,G17412,G17413);
  nand GNAME14477(G14477,G15426,G17408,G17406,G17407);
  nand GNAME14478(G14478,G15425,G17402,G17400,G17401);
  nand GNAME14479(G14479,G15424,G17383,G17381,G17382);
  nand GNAME14480(G14480,G15423,G17377,G17375,G17376);
  nand GNAME14481(G14481,G15422,G17371,G17369,G17370);
  nand GNAME14482(G14482,G15421,G17365,G17363,G17364);
  nand GNAME14483(G14483,G15420,G17359,G17357,G17358);
  nand GNAME14484(G14484,G15419,G17353,G17351,G17352);
  nand GNAME14485(G14485,G15418,G17347,G17345,G17346);
  nand GNAME14486(G14486,G15417,G17341,G17339,G17340);
  nand GNAME14487(G14487,G15416,G17322,G17320,G17321);
  nand GNAME14488(G14488,G15415,G17316,G17314,G17315);
  nand GNAME14489(G14489,G15414,G17310,G17308,G17309);
  nand GNAME14490(G14490,G15413,G17304,G17302,G17303);
  nand GNAME14491(G14491,G15412,G17298,G17296,G17297);
  nand GNAME14492(G14492,G15411,G17292,G17290,G17291);
  nand GNAME14493(G14493,G15410,G17286,G17284,G17285);
  nand GNAME14494(G14494,G15409,G17280,G17278,G17279);
  nand GNAME14495(G14495,G15408,G17261,G17259,G17260);
  nand GNAME14496(G14496,G15407,G17252,G17250,G17251);
  nand GNAME14497(G14497,G15406,G17243,G17241,G17242);
  nand GNAME14498(G14498,G15405,G17234,G17232,G17233);
  nand GNAME14499(G14499,G15404,G17225,G17223,G17224);
  nand GNAME14500(G14500,G15403,G17216,G17214,G17215);
  nand GNAME14501(G14501,G15402,G17207,G17205,G17206);
  nand GNAME14502(G14502,G15401,G17198,G17196,G17197);
  and GNAME14503(G14503,G17037,G60011);
  nand GNAME14504(G14504,G17073,G17071,G17072);
  nand GNAME14505(G14505,G17066,G17064,G17065);
  nand GNAME14506(G14506,G17055,G17053,G17054);
  nand GNAME14507(G14507,G15395,G17029,G17031,G17032);
  nand GNAME14508(G14508,G15394,G17023,G17025,G17026);
  nand GNAME14509(G14509,G15393,G17017,G17019,G17020);
  nand GNAME14510(G14510,G15392,G17011,G17013,G17014);
  nand GNAME14511(G14511,G15391,G17009,G17007,G17008);
  nand GNAME14512(G14512,G15390,G17003,G17001,G17002);
  nand GNAME14513(G14513,G15389,G16997,G16995,G16996);
  nand GNAME14514(G14514,G15388,G16991,G16989,G16990);
  nand GNAME14515(G14515,G15387,G16985,G16983,G16984);
  nand GNAME14516(G14516,G15386,G16979,G16977,G16978);
  nand GNAME14517(G14517,G15385,G16973,G16971,G16972);
  nand GNAME14518(G14518,G15384,G16967,G16965,G16966);
  nand GNAME14519(G14519,G15383,G16961,G16959,G16960);
  nand GNAME14520(G14520,G15382,G16955,G16953,G16954);
  nand GNAME14521(G14521,G15381,G16949,G16947,G16948);
  nand GNAME14522(G14522,G15380,G16943,G16941,G16942);
  nand GNAME14523(G14523,G15379,G16937,G16935,G16936);
  nand GNAME14524(G14524,G15378,G16931,G16929,G16930);
  nand GNAME14525(G14525,G15377,G16925,G16923,G16924);
  nand GNAME14526(G14526,G15376,G16919,G16917,G16918);
  nand GNAME14527(G14527,G15375,G16913,G16911,G16912);
  nand GNAME14528(G14528,G15374,G16907,G16905,G16906);
  nand GNAME14529(G14529,G15373,G16901,G16899,G16900);
  nand GNAME14530(G14530,G15372,G16895,G16893,G16894);
  nand GNAME14531(G14531,G15371,G16889,G16887,G16888);
  nand GNAME14532(G14532,G15370,G16883,G16881,G16882);
  nand GNAME14533(G14533,G15369,G16877,G16875,G16876);
  nand GNAME14534(G14534,G15368,G16871,G16869,G16870);
  nand GNAME14535(G14535,G15367,G16865,G16863,G16864);
  nand GNAME14536(G14536,G15366,G16859,G16857,G16858);
  nand GNAME14537(G14537,G15365,G16853,G16851,G16852);
  nand GNAME14538(G14538,G15364,G16847,G16845,G16846);
  nand GNAME14539(G14539,G16804,G16805,G16803,G16801,G16802);
  nand GNAME14540(G14540,G16799,G16800,G16798,G16796,G16797);
  nand GNAME14541(G14541,G16794,G16795,G16793,G16791,G16792);
  nand GNAME14542(G14542,G16789,G16790,G16788,G16786,G16787);
  nand GNAME14543(G14543,G16784,G16785,G16783,G16781,G16782);
  nand GNAME14544(G14544,G16779,G16780,G16778,G16776,G16777);
  nand GNAME14545(G14545,G16774,G16775,G16773,G16771,G16772);
  nand GNAME14546(G14546,G16769,G16770,G16768,G16766,G16767);
  nand GNAME14547(G14547,G16764,G16765,G16763,G16761,G16762);
  nand GNAME14548(G14548,G16759,G16760,G16758,G16756,G16757);
  nand GNAME14549(G14549,G16754,G16755,G16753,G16751,G16752);
  nand GNAME14550(G14550,G16749,G16750,G16748,G16746,G16747);
  nand GNAME14551(G14551,G16744,G16745,G16743,G16741,G16742);
  nand GNAME14552(G14552,G16739,G16740,G16738,G16736,G16737);
  nand GNAME14553(G14553,G16734,G16735,G16733,G16731,G16732);
  nand GNAME14554(G14554,G16729,G16730,G16728,G16726,G16727);
  nand GNAME14555(G14555,G16724,G16725,G16723,G16721,G16722);
  nand GNAME14556(G14556,G16719,G16720,G16718,G16716,G16717);
  nand GNAME14557(G14557,G16714,G16715,G16713,G16711,G16712);
  nand GNAME14558(G14558,G16709,G16710,G16708,G16706,G16707);
  nand GNAME14559(G14559,G16704,G16705,G16703,G16701,G16702);
  nand GNAME14560(G14560,G16699,G16700,G16698,G16696,G16697);
  nand GNAME14561(G14561,G16694,G16695,G16693,G16691,G16692);
  nand GNAME14562(G14562,G16689,G16690,G16688,G16686,G16687);
  nand GNAME14563(G14563,G16684,G16685,G16683,G16681,G16682);
  nand GNAME14564(G14564,G16679,G16680,G16678,G16676,G16677);
  nand GNAME14565(G14565,G16674,G16675,G16673,G16671,G16672);
  nand GNAME14566(G14566,G16669,G16670,G16668,G16666,G16667);
  nand GNAME14567(G14567,G16664,G16665,G16663,G16661,G16662);
  nand GNAME14568(G14568,G16659,G16660,G16658,G16656,G16657);
  nand GNAME14569(G14569,G16654,G16655,G16653,G16651,G16652);
  nand GNAME14570(G14570,G16649,G16650,G16648,G16646,G16647);
  nand GNAME14571(G14571,G16644,G16642,G16643);
  nand GNAME14572(G14572,G16641,G16639,G16640);
  nand GNAME14573(G14573,G16638,G16636,G16637);
  nand GNAME14574(G14574,G16635,G16633,G16634);
  nand GNAME14575(G14575,G16632,G16630,G16631);
  nand GNAME14576(G14576,G16629,G16627,G16628);
  nand GNAME14577(G14577,G16626,G16624,G16625);
  nand GNAME14578(G14578,G16623,G16621,G16622);
  nand GNAME14579(G14579,G16620,G16618,G16619);
  nand GNAME14580(G14580,G16617,G16615,G16616);
  nand GNAME14581(G14581,G16614,G16612,G16613);
  nand GNAME14582(G14582,G16611,G16609,G16610);
  nand GNAME14583(G14583,G16608,G16606,G16607);
  nand GNAME14584(G14584,G16605,G16603,G16604);
  nand GNAME14585(G14585,G16602,G16600,G16601);
  nand GNAME14586(G14586,G16599,G16597,G16598);
  nand GNAME14587(G14587,G16596,G16595,G16639);
  nand GNAME14588(G14588,G16594,G16593,G16636);
  nand GNAME14589(G14589,G16592,G16591,G16633);
  nand GNAME14590(G14590,G16590,G16589,G16630);
  nand GNAME14591(G14591,G16588,G16587,G16627);
  nand GNAME14592(G14592,G16586,G16585,G16624);
  nand GNAME14593(G14593,G16584,G16583,G16621);
  nand GNAME14594(G14594,G16620,G16581,G16582);
  nand GNAME14595(G14595,G16617,G16579,G16580);
  nand GNAME14596(G14596,G16614,G16577,G16578);
  nand GNAME14597(G14597,G16611,G16575,G16576);
  nand GNAME14598(G14598,G16608,G16573,G16574);
  nand GNAME14599(G14599,G16605,G16571,G16572);
  nand GNAME14600(G14600,G16602,G16569,G16570);
  nand GNAME14601(G14601,G16599,G16567,G16568);
  nand GNAME14602(G14602,G16564,G16562,G16563);
  nand GNAME14603(G14603,G16561,G16559,G16560);
  nand GNAME14604(G14604,G16558,G16556,G16557);
  nand GNAME14605(G14605,G16555,G16553,G16554);
  nand GNAME14606(G14606,G16552,G16550,G16551);
  nand GNAME14607(G14607,G16549,G16547,G16548);
  nand GNAME14608(G14608,G16546,G16544,G16545);
  nand GNAME14609(G14609,G16543,G16541,G16542);
  nand GNAME14610(G14610,G16540,G16538,G16539);
  nand GNAME14611(G14611,G16537,G16535,G16536);
  nand GNAME14612(G14612,G16534,G16532,G16533);
  nand GNAME14613(G14613,G16531,G16529,G16530);
  nand GNAME14614(G14614,G16528,G16526,G16527);
  nand GNAME14615(G14615,G16525,G16523,G16524);
  nand GNAME14616(G14616,G16522,G16520,G16521);
  nand GNAME14617(G14617,G16519,G16517,G16518);
  nand GNAME14618(G14618,G16516,G16514,G16515);
  nand GNAME14619(G14619,G16513,G16511,G16512);
  nand GNAME14620(G14620,G16510,G16508,G16509);
  nand GNAME14621(G14621,G16507,G16505,G16506);
  nand GNAME14622(G14622,G16504,G16502,G16503);
  nand GNAME14623(G14623,G16501,G16499,G16500);
  nand GNAME14624(G14624,G16498,G16496,G16497);
  nand GNAME14625(G14625,G16495,G16493,G16494);
  nand GNAME14626(G14626,G16492,G16490,G16491);
  nand GNAME14627(G14627,G16489,G16487,G16488);
  nand GNAME14628(G14628,G16486,G16484,G16485);
  nand GNAME14629(G14629,G16483,G16481,G16482);
  nand GNAME14630(G14630,G16480,G16478,G16479);
  nand GNAME14631(G14631,G16477,G16475,G16476);
  nand GNAME14632(G14632,G16474,G16472,G16473);
  and GNAME14633(G14633,G14870,G60142);
  nand GNAME14634(G14634,G16463,G16464,G16465,G16466);
  nand GNAME14635(G14635,G16459,G16460,G16461,G16462);
  nand GNAME14636(G14636,G16455,G16456,G16457,G16458);
  nand GNAME14637(G14637,G16451,G16452,G16453,G16454);
  nand GNAME14638(G14638,G16447,G16448,G16449,G16450);
  nand GNAME14639(G14639,G16443,G16444,G16445,G16446);
  nand GNAME14640(G14640,G16439,G16440,G16441,G16442);
  nand GNAME14641(G14641,G16435,G16436,G16437,G16438);
  nand GNAME14642(G14642,G16431,G16432,G16433,G16434);
  nand GNAME14643(G14643,G16427,G16428,G16429,G16430);
  nand GNAME14644(G14644,G16423,G16424,G16425,G16426);
  nand GNAME14645(G14645,G16419,G16420,G16421,G16422);
  nand GNAME14646(G14646,G16415,G16416,G16417,G16418);
  nand GNAME14647(G14647,G16411,G16412,G16413,G16414);
  nand GNAME14648(G14648,G16407,G16408,G16409,G16410);
  nand GNAME14649(G14649,G16403,G16404,G16405,G16406);
  nand GNAME14650(G14650,G16401,G16402,G16400,G16398,G16399);
  nand GNAME14651(G14651,G16396,G16397,G16395,G16393,G16394);
  nand GNAME14652(G14652,G16391,G16392,G16390,G16388,G16389);
  nand GNAME14653(G14653,G16386,G16387,G16385,G16383,G16384);
  nand GNAME14654(G14654,G16381,G16382,G16380,G16378,G16379);
  nand GNAME14655(G14655,G16376,G16377,G16375,G16373,G16374);
  nand GNAME14656(G14656,G16371,G16372,G16370,G16368,G16369);
  nand GNAME14657(G14657,G16366,G16367,G16365,G16363,G16364);
  nand GNAME14658(G14658,G16361,G16362,G16360,G16358,G16359);
  nand GNAME14659(G14659,G16356,G16357,G16355,G16353,G16354);
  nand GNAME14660(G14660,G16351,G16352,G16350,G16348,G16349);
  nand GNAME14661(G14661,G16346,G16347,G16345,G16343,G16344);
  nand GNAME14662(G14662,G16341,G16342,G16340,G16338,G16339);
  nand GNAME14663(G14663,G16336,G16337,G16335,G16333,G16334);
  nand GNAME14664(G14664,G16331,G16332,G16330,G16328,G16329);
  nand GNAME14665(G14665,G16327,G16325,G16326);
  nand GNAME14666(G14666,G16315,G16313,G16314);
  nand GNAME14667(G14667,G16312,G16310,G16311);
  nand GNAME14668(G14668,G16309,G16307,G16308);
  nand GNAME14669(G14669,G16306,G16304,G16305);
  nand GNAME14670(G14670,G16303,G16301,G16302);
  nand GNAME14671(G14671,G16300,G16298,G16299);
  nand GNAME14672(G14672,G16297,G16295,G16296);
  nand GNAME14673(G14673,G16294,G16292,G16293);
  nand GNAME14674(G14674,G16291,G16289,G16290);
  nand GNAME14675(G14675,G16288,G16286,G16287);
  nand GNAME14676(G14676,G16285,G16283,G16284);
  nand GNAME14677(G14677,G16282,G16280,G16281);
  nand GNAME14678(G14678,G16279,G16277,G16278);
  nand GNAME14679(G14679,G16276,G16274,G16275);
  nand GNAME14680(G14680,G16273,G16271,G16272);
  nand GNAME14681(G14681,G16270,G16268,G16269);
  nand GNAME14682(G14682,G16267,G16265,G16266);
  nand GNAME14683(G14683,G16264,G16262,G16263);
  nand GNAME14684(G14684,G16261,G16259,G16260);
  nand GNAME14685(G14685,G16258,G16256,G16257);
  nand GNAME14686(G14686,G16255,G16253,G16254);
  nand GNAME14687(G14687,G16252,G16250,G16251);
  nand GNAME14688(G14688,G16249,G16247,G16248);
  nand GNAME14689(G14689,G16246,G16244,G16245);
  nand GNAME14690(G14690,G16243,G16241,G16242);
  nand GNAME14691(G14691,G16240,G16238,G16239);
  nand GNAME14692(G14692,G16237,G16235,G16236);
  nand GNAME14693(G14693,G16234,G16232,G16233);
  nand GNAME14694(G14694,G16231,G16229,G16230);
  nand GNAME14695(G14695,G16228,G16226,G16227);
  nand GNAME14696(G14696,G16225,G16223,G16224);
  nand GNAME14697(G14697,G16221,G16222);
  nand GNAME14698(G14698,G15359,G16212,G16214,G16215);
  nand GNAME14699(G14699,G15358,G16206,G16208,G16209);
  nand GNAME14700(G14700,G16204,G15357,G16201,G16199,G16200);
  nand GNAME14701(G14701,G16198,G15356,G16195,G16193,G16194);
  nand GNAME14702(G14702,G15355,G16188,G16190,G16191);
  nand GNAME14703(G14703,G15354,G16182,G16184,G16185);
  nand GNAME14704(G14704,G15353,G16174,G16171,G16172,G16173);
  nand GNAME14705(G14705,G15352,G16168,G16165,G16166,G16167);
  nand GNAME14706(G14706,G15351,G16162,G16159,G16160,G16161);
  nand GNAME14707(G14707,G15350,G16156,G16153,G16154,G16157);
  nand GNAME14708(G14708,G15349,G16151,G16147,G16148,G16149);
  nand GNAME14709(G14709,G15348,G16145,G16141,G16142,G16143);
  nand GNAME14710(G14710,G15347,G16139,G16135,G16136,G16137);
  nand GNAME14711(G14711,G15346,G16133,G16129,G16130,G16131);
  nand GNAME14712(G14712,G15345,G16127,G16123,G16124,G16125);
  nand GNAME14713(G14713,G15344,G16121,G16117,G16118,G16119);
  nand GNAME14714(G14714,G15343,G16115,G16111,G16112,G16113);
  nand GNAME14715(G14715,G15342,G16109,G16105,G16106,G16107);
  nand GNAME14716(G14716,G15341,G16103,G16099,G16100,G16101);
  nand GNAME14717(G14717,G15340,G16097,G16093,G16094,G16095);
  nand GNAME14718(G14718,G15339,G16090,G16086,G16087);
  nand GNAME14719(G14719,G15338,G16084,G16080,G16081);
  nand GNAME14720(G14720,G15337,G16078,G16074,G16075);
  nand GNAME14721(G14721,G15336,G16072,G16068,G16069);
  nand GNAME14722(G14722,G15335,G16066,G16062,G16063);
  nand GNAME14723(G14723,G15334,G16060,G16056,G16057);
  nand GNAME14724(G14724,G15333,G16054,G16050,G16051);
  nand GNAME14725(G14725,G15332,G16048,G16044,G16045);
  nand GNAME14726(G14726,G15331,G16042,G16038,G16039);
  nand GNAME14727(G14727,G15330,G16036,G16032,G16033);
  nand GNAME14728(G14728,G15329,G16030,G16026,G16027);
  nand GNAME14729(G14729,G15328,G16024,G16020,G16021);
  nand GNAME14730(G14730,G16008,G15805,G14828);
  nand GNAME14731(G14731,G16007,G16005,G16006);
  nand GNAME14732(G14732,G16003,G15805,G14829);
  nand GNAME14733(G14733,G14829,G19847,G19848);
  nand GNAME14734(G14734,G16001,G16000);
  nand GNAME14735(G14735,G15998,G15999);
  nand GNAME14736(G14736,G15811,G19840,G19841);
  nand GNAME14737(G14737,G15811,G19836,G19837);
  nand GNAME14738(G14738,G15967,G15968);
  nand GNAME14739(G14739,G15959,G15958);
  and GNAME14740(G14740,G14777,G15846);
  nand GNAME14741(G14741,G19857,G19858,G17044,G17045);
  and GNAME14742(G14742,G14793,G15829);
  nand GNAME14743(G14743,G15296,G15297,G15298,G15299);
  and GNAME14744(G14744,G18181,G15101);
  not GNAME14745(G14745,G33);
  not GNAME14746(G14746,G1589);
  nand GNAME14747(G14747,G14888,G15829,G15846);
  not GNAME14748(G14748,G59875);
  not GNAME14749(G14749,G60010);
  and GNAME14750(G14750,G14765,G14758);
  and GNAME14751(G14751,G14753,G60010);
  and GNAME14752(G14752,G14750,G14751);
  not GNAME14753(G14753,G60009);
  and GNAME14754(G14754,G14749,G60009);
  and GNAME14755(G14755,G14750,G14754);
  and GNAME14756(G14756,G60010,G60009);
  and GNAME14757(G14757,G14750,G14756);
  not GNAME14758(G14758,G60008);
  nor GNAME14759(G14759,G60007,G14758);
  nor GNAME14760(G14760,G60010,G60009);
  and GNAME14761(G14761,G14759,G14760);
  and GNAME14762(G14762,G14751,G14759);
  and GNAME14763(G14763,G14754,G14759);
  and GNAME14764(G14764,G14756,G14759);
  not GNAME14765(G14765,G60007);
  and GNAME14766(G14766,G14758,G60007);
  and GNAME14767(G14767,G14760,G14766);
  and GNAME14768(G14768,G14751,G14766);
  and GNAME14769(G14769,G14754,G14766);
  nor GNAME14770(G14770,G15784,G15785);
  nor GNAME14771(G14771,G14758,G14765);
  and GNAME14772(G14772,G14760,G14771);
  and GNAME14773(G14773,G14751,G14771);
  and GNAME14774(G14774,G14754,G14771);
  and GNAME14775(G14775,G14756,G14771);
  and GNAME14776(G14776,G14750,G14760);
  nand GNAME14777(G14777,G15312,G15313,G15314,G15315);
  nand GNAME14778(G14778,G15316,G15317,G15318,G15319);
  nand GNAME14779(G14779,G15300,G15301,G15302,G15303);
  nand GNAME14780(G14780,G15304,G15305,G15306,G15307);
  and GNAME14781(G14781,G15914,G15897);
  and GNAME14782(G14782,G15880,G14742,G14789);
  and GNAME14783(G14783,G14849,G14743,G14781,G14782);
  not GNAME14784(G14784,G59877);
  and GNAME14785(G14785,G14783,G59877);
  not GNAME14786(G14786,G23753);
  and GNAME14787(G14787,G14811,G59875);
  nor GNAME14788(G14788,G15829,G14780);
  nand GNAME14789(G14789,G15288,G15289,G15290,G15291);
  and GNAME14790(G14790,G14788,G14779,G14849);
  nand GNAME14791(G14791,G14778,G15948,G15863,G14790);
  nor GNAME14792(G14792,G59876,G14784);
  nand GNAME14793(G14793,G15308,G15309,G15310,G15311);
  nor GNAME14794(G14794,G14779,G14793);
  nor GNAME14795(G14795,G14778,G15931,G15948);
  nand GNAME14796(G14796,G14794,G14795,G15897,G14789,G15829);
  and GNAME14797(G14797,G59877,G14787);
  not GNAME14798(G14798,G23088);
  and GNAME14799(G14799,G14811,G14748);
  nand GNAME14800(G14800,G14875,G15954);
  not GNAME14801(G14801,G59840);
  nand GNAME14802(G14802,G14814,G59840);
  not GNAME14803(G14803,G59841);
  or GNAME14804(G14804,G15957,G14809);
  and GNAME14805(G14805,G15961,G15802,G14849);
  and GNAME14806(G14806,G15800,G15964,G15965,G14805);
  and GNAME14807(G14807,G14831,G14799);
  and GNAME14808(G14808,G14803,G59840);
  and GNAME14809(G14809,G14801,G14803);
  and GNAME14810(G14810,G14784,G59875);
  not GNAME14811(G14811,G59876);
  nand GNAME14812(G14812,G14810,G59876);
  nor GNAME14813(G14813,G14904,G59874);
  not GNAME14814(G14814,G59839);
  nand GNAME14815(G14815,G15973,G14803);
  not GNAME14816(G14816,G60246);
  and GNAME14817(G14817,G59875,G15846);
  and GNAME14818(G14818,G15880,G14790);
  and GNAME14819(G14819,G14818,G14789,G14743);
  and GNAME14820(G14820,G14849,G15914);
  and GNAME14821(G14821,G14743,G15863);
  and GNAME14822(G14822,G14820,G14821,G15880,G14740,G14780);
  and GNAME14823(G14823,G14789,G14780);
  and GNAME14824(G14824,G14793,G15914);
  and GNAME14825(G14825,G14777,G14795,G14823,G14824);
  and GNAME14826(G14826,G15321,G15323,G15325,G15327);
  not GNAME14827(G14827,G60207);
  or GNAME14828(G14828,G19982,G60208,G59843);
  nand GNAME14829(G14829,G14826,G60208);
  and GNAME14830(G14830,G14816,G59876);
  not GNAME14831(G14831,G59874);
  and GNAME14832(G14832,G14746,G14816);
  nor GNAME14833(G14833,G16009,G14748);
  and GNAME14834(G14834,G16019,G14833);
  not GNAME14835(G14835,G15279);
  nor GNAME14836(G14836,G59875,G14784);
  and GNAME14837(G14837,G14839,G14836);
  and GNAME14838(G14838,G14794,G15974,G14832,G14833);
  nand GNAME14839(G14839,G15808,G15809,G16825,G19977);
  nand GNAME14840(G14840,G16011,G16012);
  not GNAME14841(G14841,G23160);
  not GNAME14842(G14842,G23487);
  not GNAME14843(G14843,G23121);
  not GNAME14844(G14844,G23426);
  not GNAME14845(G14845,G23213);
  not GNAME14846(G14846,G23532);
  not GNAME14847(G14847,G23189);
  not GNAME14848(G14848,G23485);
  nand GNAME14849(G14849,G15292,G15293,G15294,G15295);
  and GNAME14850(G14850,G15948,G15880);
  nor GNAME14851(G14851,G15802,G14780,G14849);
  nand GNAME14852(G14852,G14742,G14789,G14779,G14851);
  and GNAME14853(G14853,G59877,G14825);
  nand GNAME14854(G14854,G16220,G14787);
  nor GNAME14855(G14855,G14743,G14854);
  nor GNAME14856(G14856,G15948,G14854);
  and GNAME14857(G14857,G14779,G15829);
  nand GNAME14858(G14858,G15863,G15846,G14851,G14857);
  and GNAME14859(G14859,G19983,G15846);
  nand GNAME14860(G14860,G59877,G14859);
  and GNAME14861(G14861,G59877,G14822);
  nand GNAME14862(G14862,G16324,G14787);
  nor GNAME14863(G14863,G15802,G14862);
  nor GNAME14864(G14864,G15880,G14862);
  nor GNAME14865(G14865,G15863,G14862);
  nor GNAME14866(G14866,G15786,G14862);
  nor GNAME14867(G14867,G14884,G14862);
  and GNAME14868(G14868,G14793,G19983);
  nand GNAME14869(G14869,G15952,G15973,G59877);
  and GNAME14870(G14870,G14812,G16471);
  nor GNAME14871(G14871,G14870,G59877);
  nor GNAME14872(G14872,G14870,G14784);
  and GNAME14873(G14873,G14789,G14872);
  nand GNAME14874(G14874,G15952,G14797);
  nand GNAME14875(G14875,G14787,G14785,G23753);
  and GNAME14876(G14876,G16565,G16566);
  nor GNAME14877(G14877,G14876,G14793);
  nor GNAME14878(G14878,G14876,G15846);
  and GNAME14879(G14879,G16000,G16645);
  nor GNAME14880(G14880,G15240,G14879);
  nor GNAME14881(G14881,G14879,G15793);
  nor GNAME14882(G14882,G14879,G14784);
  nor GNAME14883(G14883,G14879,G15794);
  and GNAME14884(G14884,G15880,G15863);
  and GNAME14885(G14885,G15360,G14805,G16810,G16811);
  nor GNAME14886(G14886,G14903,G14748);
  and GNAME14887(G14887,G14822,G14886);
  nor GNAME14888(G14888,G15802,G15931,G14789);
  and GNAME14889(G14889,G16806,G19849,G19850);
  and GNAME14890(G14890,G16807,G16831);
  and GNAME14891(G14891,G14793,G15863);
  and GNAME14892(G14892,G15362,G14890,G16836,G14889);
  and GNAME14893(G14893,G15361,G15931,G15897,G14794);
  and GNAME14894(G14894,G14788,G14891,G15948,G14778,G14779);
  and GNAME14895(G14895,G16839,G16840);
  and GNAME14896(G14896,G14852,G14895);
  and GNAME14897(G14897,G15363,G14796,G14892);
  and GNAME14898(G14898,G16841,G14886);
  and GNAME14899(G14899,G17097,G16467);
  and GNAME14900(G14900,G16829,G14886);
  and GNAME14901(G14901,G16826,G14886);
  nor GNAME14902(G14902,G59875,G14903);
  and GNAME14903(G14903,G16824,G16825);
  and GNAME14904(G14904,G59875,G59876);
  and GNAME14905(G14905,G59877,G14904);
  nand GNAME14906(G14906,G14784,G59874);
  nand GNAME14907(G14907,G17034,G19855,G19856);
  not GNAME14908(G14908,G60015);
  nor GNAME14909(G14909,G14929,G17039,G14748,G14784);
  and GNAME14910(G14910,G19862,G19863,G15791,G17038);
  nand GNAME14911(G14911,G17040,G14916);
  nor GNAME14912(G14912,G15793,G59875,G17037);
  and GNAME14913(G14913,G14914,G17043);
  nand GNAME14914(G14914,G17035,G15810,G17036);
  not GNAME14915(G14915,G60014);
  or GNAME14916(G14916,G14910,G14909);
  nand GNAME14917(G14917,G17046,G17047);
  nand GNAME14918(G14918,G17051,G17049,G17050);
  not GNAME14919(G14919,G60013);
  and GNAME14920(G14920,G60015,G60014);
  and GNAME14921(G14921,G17058,G17056,G17057);
  nand GNAME14922(G14922,G17060,G17061);
  nand GNAME14923(G14923,G17062,G15769);
  nor GNAME14924(G14924,G60012,G14919);
  not GNAME14925(G14925,G60012);
  nor GNAME14926(G14926,G59875,G14798);
  nand GNAME14927(G14927,G17086,G60010);
  nand GNAME14928(G14928,G17092,G14930);
  and GNAME14929(G14929,G19861,G59876);
  nand GNAME14930(G14930,G17089,G17090);
  nand GNAME14931(G14931,G17114,G17115);
  nand GNAME14932(G14932,G17136,G17137);
  nand GNAME14933(G14933,G17133,G17134);
  nand GNAME14934(G14934,G17139,G15774);
  nand GNAME14935(G14935,G17168,G19898,G19899);
  nand GNAME14936(G14936,G17163,G17165);
  and GNAME14937(G14937,G59876,G60246);
  nand GNAME14938(G14938,G17161,G17156);
  nor GNAME14939(G14939,G19883,G14938);
  nor GNAME14940(G14940,G17093,G19889);
  nor GNAME14941(G14941,G17035,G15792);
  nor GNAME14942(G14942,G19876,G15247);
  nor GNAME14943(G14943,G17063,G17041);
  nand GNAME14944(G14944,G14942,G14943);
  nor GNAME14945(G14945,G14957,G19980);
  and GNAME14946(G14946,G17183,G14945);
  nor GNAME14947(G14947,G60013,G60012);
  nor GNAME14948(G14948,G60014,G60015);
  or GNAME14949(G14949,G14979,G14990);
  or GNAME14950(G14950,G17067,G15035,G15042);
  nor GNAME14951(G14951,G15248,G14950);
  nor GNAME14952(G14952,G14908,G14949);
  and GNAME14953(G14953,G14951,G14952);
  and GNAME14954(G14954,G14947,G14948);
  nor GNAME14955(G14955,G14953,G17188);
  and GNAME14956(G14956,G14907,G1691);
  and GNAME14957(G14957,G14939,G14940);
  and GNAME14958(G14958,G1675,G14941);
  nor GNAME14959(G14959,G17035,G15794);
  and GNAME14960(G14960,G14907,G1680);
  and GNAME14961(G14961,G1674,G14941);
  and GNAME14962(G14962,G14907,G1669);
  and GNAME14963(G14963,G1673,G14941);
  and GNAME14964(G14964,G14907,G1666);
  and GNAME14965(G14965,G1672,G14941);
  and GNAME14966(G14966,G14907,G1665);
  and GNAME14967(G14967,G1671,G14941);
  and GNAME14968(G14968,G14907,G1664);
  and GNAME14969(G14969,G1670,G14941);
  and GNAME14970(G14970,G14907,G1663);
  and GNAME14971(G14971,G1668,G14941);
  and GNAME14972(G14972,G14907,G1662);
  and GNAME14973(G14973,G1667,G14941);
  nor GNAME14974(G14974,G19889,G14928);
  nor GNAME14975(G14975,G17063,G14911);
  nand GNAME14976(G14976,G14942,G14975);
  nor GNAME14977(G14977,G14984,G19980);
  and GNAME14978(G14978,G17265,G14977);
  and GNAME14979(G14979,G14915,G60015);
  nor GNAME14980(G14980,G60015,G14949);
  and GNAME14981(G14981,G14951,G14980);
  and GNAME14982(G14982,G14947,G14979);
  nor GNAME14983(G14983,G14981,G17270);
  and GNAME14984(G14984,G14939,G14974);
  nor GNAME14985(G14985,G15250,G14938);
  nor GNAME14986(G14986,G19870,G19876);
  nand GNAME14987(G14987,G14943,G14986);
  nor GNAME14988(G14988,G14995,G19980);
  and GNAME14989(G14989,G17326,G14988);
  and GNAME14990(G14990,G14908,G60014);
  and GNAME14991(G14991,G14949,G60015);
  and GNAME14992(G14992,G14951,G14991);
  and GNAME14993(G14993,G14947,G14990);
  nor GNAME14994(G14994,G14992,G17331);
  and GNAME14995(G14995,G14940,G14985);
  nand GNAME14996(G14996,G14975,G14986);
  nor GNAME14997(G14997,G15003,G19980);
  and GNAME14998(G14998,G17387,G14997);
  and GNAME14999(G14999,G14949,G14908);
  and GNAME15000(G15000,G14951,G14999);
  and GNAME15001(G15001,G14920,G14947);
  nor GNAME15002(G15002,G15000,G17392);
  and GNAME15003(G15003,G14974,G14985);
  nor GNAME15004(G15004,G17093,G15261);
  nor GNAME15005(G15005,G17041,G14923);
  nand GNAME15006(G15006,G14942,G15005);
  nor GNAME15007(G15007,G15013,G19980);
  and GNAME15008(G15008,G17448,G15007);
  nor GNAME15009(G15009,G19873,G14950);
  and GNAME15010(G15010,G14952,G15009);
  and GNAME15011(G15011,G14924,G14948);
  nor GNAME15012(G15012,G15010,G17453);
  and GNAME15013(G15013,G14939,G15004);
  nor GNAME15014(G15014,G14928,G15261);
  nor GNAME15015(G15015,G14911,G14923);
  nand GNAME15016(G15016,G14942,G15015);
  nor GNAME15017(G15017,G15022,G19980);
  and GNAME15018(G15018,G17509,G15017);
  and GNAME15019(G15019,G14980,G15009);
  and GNAME15020(G15020,G14924,G14979);
  nor GNAME15021(G15021,G15019,G17514);
  and GNAME15022(G15022,G14939,G15014);
  nand GNAME15023(G15023,G14986,G15005);
  nor GNAME15024(G15024,G15029,G19980);
  and GNAME15025(G15025,G17570,G15024);
  and GNAME15026(G15026,G14991,G15009);
  and GNAME15027(G15027,G14924,G14990);
  nor GNAME15028(G15028,G15026,G17575);
  and GNAME15029(G15029,G14985,G15004);
  nand GNAME15030(G15030,G14986,G15015);
  nor GNAME15031(G15031,G15036,G19980);
  and GNAME15032(G15032,G17631,G15031);
  and GNAME15033(G15033,G14999,G15009);
  nor GNAME15034(G15034,G15033,G17636);
  and GNAME15035(G15035,G14920,G14924);
  and GNAME15036(G15036,G14985,G15014);
  nor GNAME15037(G15037,G17162,G19883);
  nor GNAME15038(G15038,G15249,G15247);
  nand GNAME15039(G15039,G14943,G15038);
  nor GNAME15040(G15040,G15047,G19980);
  and GNAME15041(G15041,G17692,G15040);
  and GNAME15042(G15042,G14919,G60012);
  and GNAME15043(G15043,G14950,G19873);
  and GNAME15044(G15044,G14952,G15043);
  and GNAME15045(G15045,G14948,G15042);
  nor GNAME15046(G15046,G15044,G17697);
  and GNAME15047(G15047,G14940,G15037);
  nand GNAME15048(G15048,G14975,G15038);
  nor GNAME15049(G15049,G15054,G19980);
  and GNAME15050(G15050,G17753,G15049);
  and GNAME15051(G15051,G14980,G15043);
  and GNAME15052(G15052,G14979,G15042);
  nor GNAME15053(G15053,G15051,G17758);
  and GNAME15054(G15054,G14974,G15037);
  nor GNAME15055(G15055,G17162,G15250);
  nor GNAME15056(G15056,G19870,G15249);
  nand GNAME15057(G15057,G14943,G15056);
  nor GNAME15058(G15058,G15063,G19980);
  and GNAME15059(G15059,G17814,G15058);
  and GNAME15060(G15060,G14991,G15043);
  and GNAME15061(G15061,G14990,G15042);
  nor GNAME15062(G15062,G15060,G17819);
  and GNAME15063(G15063,G14940,G15055);
  nand GNAME15064(G15064,G14975,G15056);
  nor GNAME15065(G15065,G15070,G19980);
  and GNAME15066(G15066,G17875,G15065);
  and GNAME15067(G15067,G14999,G15043);
  and GNAME15068(G15068,G14920,G15042);
  nor GNAME15069(G15069,G15067,G17880);
  and GNAME15070(G15070,G14974,G15055);
  nand GNAME15071(G15071,G15005,G15038);
  nor GNAME15072(G15072,G15079,G19980);
  and GNAME15073(G15073,G17936,G15072);
  nor GNAME15074(G15074,G14919,G14925);
  and GNAME15075(G15075,G14950,G15248);
  and GNAME15076(G15076,G14952,G15075);
  and GNAME15077(G15077,G14948,G15074);
  nor GNAME15078(G15078,G15076,G17941);
  and GNAME15079(G15079,G15004,G15037);
  nand GNAME15080(G15080,G15015,G15038);
  nor GNAME15081(G15081,G15086,G19980);
  and GNAME15082(G15082,G17997,G15081);
  and GNAME15083(G15083,G14980,G15075);
  and GNAME15084(G15084,G14979,G15074);
  nor GNAME15085(G15085,G15083,G18002);
  and GNAME15086(G15086,G15014,G15037);
  nand GNAME15087(G15087,G15005,G15056);
  nor GNAME15088(G15088,G15093,G19980);
  and GNAME15089(G15089,G18058,G15088);
  and GNAME15090(G15090,G14991,G15075);
  and GNAME15091(G15091,G14990,G15074);
  nor GNAME15092(G15092,G15090,G18063);
  and GNAME15093(G15093,G15004,G15055);
  nand GNAME15094(G15094,G15015,G15056);
  nor GNAME15095(G15095,G15100,G19980);
  and GNAME15096(G15096,G18119,G15095);
  and GNAME15097(G15097,G14999,G15075);
  nor GNAME15098(G15098,G15097,G18124);
  and GNAME15099(G15099,G14920,G15074);
  and GNAME15100(G15100,G15014,G15055);
  and GNAME15101(G15101,G15986,G14806);
  and GNAME15102(G15102,G15790,G15789);
  nor GNAME15103(G15103,G15529,G14744,G23764,G14819);
  nand GNAME15104(G15104,G19904,G19905,G18186,G59875);
  nor GNAME15105(G15105,G59876,G59874);
  not GNAME15106(G15106,G34);
  nand GNAME15107(G15107,G18202,G59839);
  and GNAME15108(G15108,G14814,G14808);
  and GNAME15109(G15109,G14808,G59839);
  nor GNAME15110(G15110,G23532,G23426);
  nor GNAME15111(G15111,G23487,G14848);
  and GNAME15112(G15112,G15110,G15111);
  nor GNAME15113(G15113,G23426,G14846);
  nor GNAME15114(G15114,G23485,G23487);
  and GNAME15115(G15115,G15113,G15114);
  and GNAME15116(G15116,G15111,G15113);
  nor GNAME15117(G15117,G23532,G14844);
  and GNAME15118(G15118,G15114,G15117);
  and GNAME15119(G15119,G15111,G15117);
  nor GNAME15120(G15120,G14844,G14846);
  and GNAME15121(G15121,G15114,G15120);
  and GNAME15122(G15122,G15111,G15120);
  nor GNAME15123(G15123,G23485,G14842);
  and GNAME15124(G15124,G15110,G15123);
  nor GNAME15125(G15125,G14842,G14848);
  and GNAME15126(G15126,G15110,G15125);
  and GNAME15127(G15127,G15113,G15123);
  and GNAME15128(G15128,G15113,G15125);
  and GNAME15129(G15129,G15117,G15123);
  and GNAME15130(G15130,G15117,G15125);
  and GNAME15131(G15131,G15120,G15123);
  and GNAME15132(G15132,G15120,G15125);
  and GNAME15133(G15133,G15110,G15114);
  nand GNAME15134(G15134,G15785,G19927,G19928);
  nor GNAME15135(G15135,G15253,G15134);
  and GNAME15136(G15136,G14756,G15135);
  and GNAME15137(G15137,G14760,G15135);
  and GNAME15138(G15138,G14751,G15135);
  nor GNAME15139(G15139,G19926,G15134);
  and GNAME15140(G15140,G14754,G15139);
  and GNAME15141(G15141,G14756,G15139);
  and GNAME15142(G15142,G14760,G15139);
  and GNAME15143(G15143,G14751,G15139);
  nor GNAME15144(G15144,G18431,G15253);
  and GNAME15145(G15145,G14754,G15144);
  and GNAME15146(G15146,G14756,G15144);
  and GNAME15147(G15147,G14760,G15144);
  and GNAME15148(G15148,G14751,G15144);
  nor GNAME15149(G15149,G18431,G19926);
  and GNAME15150(G15150,G14754,G15149);
  and GNAME15151(G15151,G14756,G15149);
  and GNAME15152(G15152,G14760,G15149);
  and GNAME15153(G15153,G14751,G15149);
  and GNAME15154(G15154,G14754,G15135);
  nor GNAME15155(G15155,G15803,G19895);
  nor GNAME15156(G15156,G17119,G14749);
  and GNAME15157(G15157,G15155,G15156);
  nand GNAME15158(G15158,G17118,G60009);
  nor GNAME15159(G15159,G60010,G15158);
  and GNAME15160(G15160,G15155,G15159);
  nor GNAME15161(G15161,G14749,G15158);
  and GNAME15162(G15162,G15155,G15161);
  nor GNAME15163(G15163,G15803,G15251);
  nor GNAME15164(G15164,G60010,G17119);
  and GNAME15165(G15165,G15163,G15164);
  and GNAME15166(G15166,G15156,G15163);
  and GNAME15167(G15167,G15159,G15163);
  and GNAME15168(G15168,G15161,G15163);
  nor GNAME15169(G15169,G19895,G14936);
  and GNAME15170(G15170,G15164,G15169);
  and GNAME15171(G15171,G15156,G15169);
  and GNAME15172(G15172,G15159,G15169);
  and GNAME15173(G15173,G15161,G15169);
  nor GNAME15174(G15174,G15251,G14936);
  and GNAME15175(G15175,G15164,G15174);
  and GNAME15176(G15176,G15156,G15174);
  and GNAME15177(G15177,G15159,G15174);
  and GNAME15178(G15178,G15161,G15174);
  and GNAME15179(G15179,G15155,G15164);
  nor GNAME15180(G15180,G23088,G15846);
  and GNAME15181(G15181,G14788,G15180);
  nand GNAME15182(G15182,G15829,G14789,G15973);
  nor GNAME15183(G15183,G14793,G15182);
  or GNAME15184(G15184,G14751,G14754);
  nor GNAME15185(G15185,G17169,G15184);
  nor GNAME15186(G15186,G60010,G17140);
  and GNAME15187(G15187,G15185,G15186);
  nor GNAME15188(G15188,G17117,G17169);
  nor GNAME15189(G15189,G17140,G14749);
  and GNAME15190(G15190,G15188,G15189);
  and GNAME15191(G15191,G15186,G15188);
  nor GNAME15192(G15192,G14749,G14934);
  and GNAME15193(G15193,G15185,G15192);
  nor GNAME15194(G15194,G60010,G14934);
  and GNAME15195(G15195,G15185,G15194);
  and GNAME15196(G15196,G15188,G15192);
  and GNAME15197(G15197,G15188,G15194);
  nor GNAME15198(G15198,G14935,G15184);
  and GNAME15199(G15199,G15189,G15198);
  and GNAME15200(G15200,G15186,G15198);
  nor GNAME15201(G15201,G17117,G14935);
  and GNAME15202(G15202,G15189,G15201);
  and GNAME15203(G15203,G15186,G15201);
  and GNAME15204(G15204,G15192,G15198);
  and GNAME15205(G15205,G15194,G15198);
  and GNAME15206(G15206,G15192,G15201);
  and GNAME15207(G15207,G15194,G15201);
  and GNAME15208(G15208,G15185,G15189);
  nor GNAME15209(G15209,G23121,G23160);
  nor GNAME15210(G15210,G23213,G14847);
  and GNAME15211(G15211,G15209,G15210);
  nor GNAME15212(G15212,G23189,G14845);
  and GNAME15213(G15213,G15209,G15212);
  nor GNAME15214(G15214,G14845,G14847);
  and GNAME15215(G15215,G15209,G15214);
  nor GNAME15216(G15216,G23160,G14843);
  nor GNAME15217(G15217,G23189,G23213);
  and GNAME15218(G15218,G15216,G15217);
  and GNAME15219(G15219,G15210,G15216);
  and GNAME15220(G15220,G15212,G15216);
  and GNAME15221(G15221,G15214,G15216);
  nor GNAME15222(G15222,G23121,G14841);
  and GNAME15223(G15223,G15217,G15222);
  and GNAME15224(G15224,G15210,G15222);
  and GNAME15225(G15225,G15212,G15222);
  and GNAME15226(G15226,G15214,G15222);
  nor GNAME15227(G15227,G14841,G14843);
  and GNAME15228(G15228,G15217,G15227);
  and GNAME15229(G15229,G15210,G15227);
  and GNAME15230(G15230,G15212,G15227);
  and GNAME15231(G15231,G15214,G15227);
  and GNAME15232(G15232,G15209,G15217);
  and GNAME15233(G15233,G23088,G14793,G14788);
  and GNAME15234(G15234,G14740,G14789);
  and GNAME15235(G15235,G59877,G14819);
  and GNAME15236(G15236,G19440,G14860);
  and GNAME15237(G15237,G19965,G19966,G19443,G14890);
  and GNAME15238(G15238,G19461,G14869);
  and GNAME15239(G15239,G14860,G19502);
  and GNAME15240(G15240,G15792,G15796);
  and GNAME15241(G15241,G59877,G16316);
  nand GNAME15242(G15242,G15105,G14779,G14743);
  nor GNAME15243(G15243,G15948,G15829,G15846);
  and GNAME15244(G15244,G19812,G15105);
  nor GNAME15245(G15245,G59874,G19799);
  nand GNAME15246(G15246,G19842,G19843);
  nand GNAME15247(G15247,G19868,G19869);
  nand GNAME15248(G15248,G19871,G19872);
  nand GNAME15249(G15249,G19874,G19875);
  nand GNAME15250(G15250,G19881,G19882);
  nand GNAME15251(G15251,G19893,G19894);
  nand GNAME15252(G15252,G19890,G19891);
  nand GNAME15253(G15253,G19924,G19925);
  nand GNAME15254(G15254,G19830,G19831);
  nand GNAME15255(G15255,G19832,G19833);
  nand GNAME15256(G15256,G19834,G19835);
  nand GNAME15257(G15257,G19838,G19839);
  nand GNAME15258(G15258,G19845,G19846);
  nand GNAME15259(G15259,G19877,G19878);
  nand GNAME15260(G15260,G19884,G19885);
  nand GNAME15261(G15261,G19887,G19888);
  nand GNAME15262(G15262,G19896,G19897);
  nand GNAME15263(G15263,G19900,G19901);
  nand GNAME15264(G15264,G19902,G19903);
  nand GNAME15265(G15265,G19908,G19909);
  nand GNAME15266(G15266,G19910,G19911);
  nand GNAME15267(G15267,G19916,G19917);
  nand GNAME15268(G15268,G19918,G19919);
  nand GNAME15269(G15269,G19920,G19921);
  nand GNAME15270(G15270,G19922,G19923);
  nand GNAME15271(G15271,G19929,G19930);
  nand GNAME15272(G15272,G19931,G19932);
  nand GNAME15273(G15273,G19933,G19934);
  nand GNAME15274(G15274,G19935,G19936);
  nand GNAME15275(G15275,G19937,G19938);
  nand GNAME15276(G15276,G19939,G19940);
  nand GNAME15277(G15277,G19941,G19942);
  nand GNAME15278(G15278,G19943,G19944);
  nand GNAME15279(G15279,G19945,G19946);
  nand GNAME15280(G15280,G19947,G19948);
  nand GNAME15281(G15281,G19949,G19950);
  nand GNAME15282(G15282,G19951,G19952);
  nand GNAME15283(G15283,G19953,G19954);
  nand GNAME15284(G15284,G19955,G19956);
  nand GNAME15285(G15285,G19957,G19958);
  nand GNAME15286(G15286,G19959,G19960);
  nand GNAME15287(G15287,G19961,G19962);
  and GNAME15288(G15288,G15847,G15848,G15849,G15850);
  and GNAME15289(G15289,G15851,G15852,G15853,G15854);
  and GNAME15290(G15290,G15855,G15856,G15857,G15858);
  and GNAME15291(G15291,G15859,G15860,G15861,G15862);
  and GNAME15292(G15292,G15915,G15916,G15917,G15918);
  and GNAME15293(G15293,G15919,G15920,G15921,G15922);
  and GNAME15294(G15294,G15923,G15924,G15925,G15926);
  and GNAME15295(G15295,G15927,G15928,G15929,G15930);
  and GNAME15296(G15296,G15932,G15933,G15934,G15935);
  and GNAME15297(G15297,G15936,G15937,G15938,G15939);
  and GNAME15298(G15298,G15940,G15941,G15942,G15943);
  and GNAME15299(G15299,G15944,G15945,G15946,G15947);
  and GNAME15300(G15300,G15898,G15899,G15900,G15901);
  and GNAME15301(G15301,G15902,G15903,G15904,G15905);
  and GNAME15302(G15302,G15906,G15907,G15908,G15909);
  and GNAME15303(G15303,G15910,G15911,G15912,G15913);
  and GNAME15304(G15304,G15881,G15882,G15883,G15884);
  and GNAME15305(G15305,G15885,G15886,G15887,G15888);
  and GNAME15306(G15306,G15889,G15890,G15891,G15892);
  and GNAME15307(G15307,G15893,G15894,G15895,G15896);
  and GNAME15308(G15308,G15830,G15831,G15832,G15833);
  and GNAME15309(G15309,G15834,G15835,G15836,G15837);
  and GNAME15310(G15310,G15838,G15839,G15840,G15841);
  and GNAME15311(G15311,G15842,G15843,G15844,G15845);
  and GNAME15312(G15312,G15813,G15814,G15815,G15816);
  and GNAME15313(G15313,G15817,G15818,G15819,G15820);
  and GNAME15314(G15314,G15821,G15822,G15823,G15824);
  and GNAME15315(G15315,G15825,G15826,G15827,G15828);
  and GNAME15316(G15316,G15864,G15865,G15866,G15867);
  and GNAME15317(G15317,G15868,G15869,G15870,G15871);
  and GNAME15318(G15318,G15872,G15873,G15874,G15875);
  and GNAME15319(G15319,G15876,G15877,G15878,G15879);
  or GNAME15320(G15320,G59847,G59846,G59845,G59844);
  nor GNAME15321(G15321,G15320,G59848,G59849,G59850,G59851);
  or GNAME15322(G15322,G59855,G59854,G59853,G59852);
  nor GNAME15323(G15323,G15322,G59856,G59857,G59858,G59859);
  or GNAME15324(G15324,G59863,G59862,G59861,G59860);
  nor GNAME15325(G15325,G15324,G59864,G59865,G59866,G59867);
  or GNAME15326(G15326,G59871,G59870,G59869,G59868);
  nor GNAME15327(G15327,G15326,G16002,G59872,G59873);
  and GNAME15328(G15328,G16025,G16023,G16022);
  and GNAME15329(G15329,G16031,G16029,G16028);
  and GNAME15330(G15330,G16037,G16035,G16034);
  and GNAME15331(G15331,G16043,G16041,G16040);
  and GNAME15332(G15332,G16049,G16047,G16046);
  and GNAME15333(G15333,G16055,G16053,G16052);
  and GNAME15334(G15334,G16061,G16059,G16058);
  and GNAME15335(G15335,G16067,G16065,G16064);
  and GNAME15336(G15336,G16073,G16071,G16070);
  and GNAME15337(G15337,G16079,G16077,G16076);
  and GNAME15338(G15338,G16085,G16083,G16082);
  and GNAME15339(G15339,G16091,G16089,G16088);
  and GNAME15340(G15340,G16098,G16096,G16092);
  and GNAME15341(G15341,G16104,G16102,G16092);
  and GNAME15342(G15342,G16110,G16108,G16092);
  and GNAME15343(G15343,G16116,G16114,G16092);
  and GNAME15344(G15344,G16122,G16120,G16092);
  and GNAME15345(G15345,G16128,G16126,G16092);
  and GNAME15346(G15346,G16134,G16132,G16092);
  and GNAME15347(G15347,G16140,G16138,G16092);
  and GNAME15348(G15348,G16146,G16144,G16092);
  and GNAME15349(G15349,G16152,G16150,G16092);
  and GNAME15350(G15350,G16158,G16092,G16155);
  and GNAME15351(G15351,G16164,G16092,G16163);
  and GNAME15352(G15352,G16170,G16092,G16169);
  and GNAME15353(G15353,G16176,G16092,G16175);
  and GNAME15354(G15354,G16092,G16181,G16186,G16183);
  and GNAME15355(G15355,G16092,G16187,G16192,G16189);
  and GNAME15356(G15356,G16196,G16197);
  and GNAME15357(G15357,G16202,G16203);
  and GNAME15358(G15358,G16207,G16205,G16210);
  and GNAME15359(G15359,G16213,G16211,G16216);
  and GNAME15360(G15360,G16809,G16806,G16807);
  and GNAME15361(G15361,G15829,G14778,G15948);
  and GNAME15362(G15362,G16835,G16833,G16834);
  and GNAME15363(G15363,G19851,G19852,G19853,G19854);
  and GNAME15364(G15364,G16844,G16842,G16843);
  and GNAME15365(G15365,G16850,G16848,G16849);
  and GNAME15366(G15366,G16856,G16854,G16855);
  and GNAME15367(G15367,G16862,G16860,G16861);
  and GNAME15368(G15368,G16868,G16866,G16867);
  and GNAME15369(G15369,G16874,G16872,G16873);
  and GNAME15370(G15370,G16880,G16878,G16879);
  and GNAME15371(G15371,G16886,G16884,G16885);
  and GNAME15372(G15372,G16892,G16890,G16891);
  and GNAME15373(G15373,G16898,G16896,G16897);
  and GNAME15374(G15374,G16904,G16902,G16903);
  and GNAME15375(G15375,G16910,G16908,G16909);
  and GNAME15376(G15376,G16916,G16914,G16915);
  and GNAME15377(G15377,G16922,G16920,G16921);
  and GNAME15378(G15378,G16928,G16926,G16927);
  and GNAME15379(G15379,G16934,G16932,G16933);
  and GNAME15380(G15380,G16940,G16938,G16939);
  and GNAME15381(G15381,G16946,G16944,G16945);
  and GNAME15382(G15382,G16952,G16950,G16951);
  and GNAME15383(G15383,G16958,G16956,G16957);
  and GNAME15384(G15384,G16964,G16962,G16963);
  and GNAME15385(G15385,G16970,G16968,G16969);
  and GNAME15386(G15386,G16976,G16974,G16975);
  and GNAME15387(G15387,G16982,G16980,G16981);
  and GNAME15388(G15388,G16988,G16986,G16987);
  and GNAME15389(G15389,G16994,G16992,G16993);
  and GNAME15390(G15390,G17000,G16998,G16999);
  and GNAME15391(G15391,G17006,G17004,G17005);
  and GNAME15392(G15392,G17012,G17010,G17015);
  and GNAME15393(G15393,G17018,G17016,G17021);
  and GNAME15394(G15394,G17024,G17022,G17027);
  and GNAME15395(G15395,G17030,G17028,G17033);
  and GNAME15396(G15396,G19866,G19867);
  and GNAME15397(G15397,G19879,G19880);
  and GNAME15398(G15398,G17126,G17124,G17121);
  and GNAME15399(G15399,G17147,G17143,G17146);
  and GNAME15400(G15400,G17175,G17171,G17174);
  and GNAME15401(G15401,G17201,G17199,G17200);
  and GNAME15402(G15402,G17210,G17208,G17209);
  and GNAME15403(G15403,G17219,G17217,G17218);
  and GNAME15404(G15404,G17228,G17226,G17227);
  and GNAME15405(G15405,G17237,G17235,G17236);
  and GNAME15406(G15406,G17246,G17244,G17245);
  and GNAME15407(G15407,G17255,G17253,G17254);
  and GNAME15408(G15408,G17264,G17262,G17263);
  and GNAME15409(G15409,G17283,G17281,G17282);
  and GNAME15410(G15410,G17289,G17287,G17288);
  and GNAME15411(G15411,G17295,G17293,G17294);
  and GNAME15412(G15412,G17301,G17299,G17300);
  and GNAME15413(G15413,G17307,G17305,G17306);
  and GNAME15414(G15414,G17313,G17311,G17312);
  and GNAME15415(G15415,G17319,G17317,G17318);
  and GNAME15416(G15416,G17325,G17323,G17324);
  and GNAME15417(G15417,G17344,G17342,G17343);
  and GNAME15418(G15418,G17350,G17348,G17349);
  and GNAME15419(G15419,G17356,G17354,G17355);
  and GNAME15420(G15420,G17362,G17360,G17361);
  and GNAME15421(G15421,G17368,G17366,G17367);
  and GNAME15422(G15422,G17374,G17372,G17373);
  and GNAME15423(G15423,G17380,G17378,G17379);
  and GNAME15424(G15424,G17386,G17384,G17385);
  and GNAME15425(G15425,G17405,G17403,G17404);
  and GNAME15426(G15426,G17411,G17409,G17410);
  and GNAME15427(G15427,G17417,G17415,G17416);
  and GNAME15428(G15428,G17423,G17421,G17422);
  and GNAME15429(G15429,G17429,G17427,G17428);
  and GNAME15430(G15430,G17435,G17433,G17434);
  and GNAME15431(G15431,G17441,G17439,G17440);
  and GNAME15432(G15432,G17447,G17445,G17446);
  and GNAME15433(G15433,G17466,G17464,G17465);
  and GNAME15434(G15434,G17472,G17470,G17471);
  and GNAME15435(G15435,G17478,G17476,G17477);
  and GNAME15436(G15436,G17484,G17482,G17483);
  and GNAME15437(G15437,G17490,G17488,G17489);
  and GNAME15438(G15438,G17496,G17494,G17495);
  and GNAME15439(G15439,G17502,G17500,G17501);
  and GNAME15440(G15440,G17508,G17506,G17507);
  and GNAME15441(G15441,G17527,G17525,G17526);
  and GNAME15442(G15442,G17533,G17531,G17532);
  and GNAME15443(G15443,G17539,G17537,G17538);
  and GNAME15444(G15444,G17545,G17543,G17544);
  and GNAME15445(G15445,G17551,G17549,G17550);
  and GNAME15446(G15446,G17557,G17555,G17556);
  and GNAME15447(G15447,G17563,G17561,G17562);
  and GNAME15448(G15448,G17569,G17567,G17568);
  and GNAME15449(G15449,G17588,G17586,G17587);
  and GNAME15450(G15450,G17594,G17592,G17593);
  and GNAME15451(G15451,G17600,G17598,G17599);
  and GNAME15452(G15452,G17606,G17604,G17605);
  and GNAME15453(G15453,G17612,G17610,G17611);
  and GNAME15454(G15454,G17618,G17616,G17617);
  and GNAME15455(G15455,G17624,G17622,G17623);
  and GNAME15456(G15456,G17630,G17628,G17629);
  and GNAME15457(G15457,G17649,G17647,G17648);
  and GNAME15458(G15458,G17655,G17653,G17654);
  and GNAME15459(G15459,G17661,G17659,G17660);
  and GNAME15460(G15460,G17667,G17665,G17666);
  and GNAME15461(G15461,G17673,G17671,G17672);
  and GNAME15462(G15462,G17679,G17677,G17678);
  and GNAME15463(G15463,G17685,G17683,G17684);
  and GNAME15464(G15464,G17691,G17689,G17690);
  and GNAME15465(G15465,G17710,G17708,G17709);
  and GNAME15466(G15466,G17716,G17714,G17715);
  and GNAME15467(G15467,G17722,G17720,G17721);
  and GNAME15468(G15468,G17728,G17726,G17727);
  and GNAME15469(G15469,G17734,G17732,G17733);
  and GNAME15470(G15470,G17740,G17738,G17739);
  and GNAME15471(G15471,G17746,G17744,G17745);
  and GNAME15472(G15472,G17752,G17750,G17751);
  and GNAME15473(G15473,G17771,G17769,G17770);
  and GNAME15474(G15474,G17777,G17775,G17776);
  and GNAME15475(G15475,G17783,G17781,G17782);
  and GNAME15476(G15476,G17789,G17787,G17788);
  and GNAME15477(G15477,G17795,G17793,G17794);
  and GNAME15478(G15478,G17801,G17799,G17800);
  and GNAME15479(G15479,G17807,G17805,G17806);
  and GNAME15480(G15480,G17813,G17811,G17812);
  and GNAME15481(G15481,G17832,G17830,G17831);
  and GNAME15482(G15482,G17838,G17836,G17837);
  and GNAME15483(G15483,G17844,G17842,G17843);
  and GNAME15484(G15484,G17850,G17848,G17849);
  and GNAME15485(G15485,G17856,G17854,G17855);
  and GNAME15486(G15486,G17862,G17860,G17861);
  and GNAME15487(G15487,G17868,G17866,G17867);
  and GNAME15488(G15488,G17874,G17872,G17873);
  and GNAME15489(G15489,G17893,G17891,G17892);
  and GNAME15490(G15490,G17899,G17897,G17898);
  and GNAME15491(G15491,G17905,G17903,G17904);
  and GNAME15492(G15492,G17911,G17909,G17910);
  and GNAME15493(G15493,G17917,G17915,G17916);
  and GNAME15494(G15494,G17923,G17921,G17922);
  and GNAME15495(G15495,G17929,G17927,G17928);
  and GNAME15496(G15496,G17935,G17933,G17934);
  and GNAME15497(G15497,G17954,G17952,G17953);
  and GNAME15498(G15498,G17960,G17958,G17959);
  and GNAME15499(G15499,G17966,G17964,G17965);
  and GNAME15500(G15500,G17972,G17970,G17971);
  and GNAME15501(G15501,G17978,G17976,G17977);
  and GNAME15502(G15502,G17984,G17982,G17983);
  and GNAME15503(G15503,G17990,G17988,G17989);
  and GNAME15504(G15504,G17996,G17994,G17995);
  and GNAME15505(G15505,G18015,G18013,G18014);
  and GNAME15506(G15506,G18021,G18019,G18020);
  and GNAME15507(G15507,G18027,G18025,G18026);
  and GNAME15508(G15508,G18033,G18031,G18032);
  and GNAME15509(G15509,G18039,G18037,G18038);
  and GNAME15510(G15510,G18045,G18043,G18044);
  and GNAME15511(G15511,G18051,G18049,G18050);
  and GNAME15512(G15512,G18057,G18055,G18056);
  and GNAME15513(G15513,G18076,G18074,G18075);
  and GNAME15514(G15514,G18082,G18080,G18081);
  and GNAME15515(G15515,G18088,G18086,G18087);
  and GNAME15516(G15516,G18094,G18092,G18093);
  and GNAME15517(G15517,G18100,G18098,G18099);
  and GNAME15518(G15518,G18106,G18104,G18105);
  and GNAME15519(G15519,G18112,G18110,G18111);
  and GNAME15520(G15520,G18118,G18116,G18117);
  and GNAME15521(G15521,G18137,G18135,G18136);
  and GNAME15522(G15522,G18143,G18141,G18142);
  and GNAME15523(G15523,G18149,G18147,G18148);
  and GNAME15524(G15524,G18155,G18153,G18154);
  and GNAME15525(G15525,G18161,G18159,G18160);
  and GNAME15526(G15526,G18167,G18165,G18166);
  and GNAME15527(G15527,G18173,G18171,G18172);
  and GNAME15528(G15528,G18179,G18177,G18178);
  nand GNAME15529(G15529,G23766,G18182,G18183);
  and GNAME15530(G15530,G18303,G18304,G18305,G18306);
  and GNAME15531(G15531,G18307,G18308,G18309,G18310);
  and GNAME15532(G15532,G18311,G18312,G18313,G18314);
  and GNAME15533(G15533,G18315,G18316,G18317,G18318);
  and GNAME15534(G15534,G18319,G18320,G18321,G18322);
  and GNAME15535(G15535,G18323,G18324,G18325,G18326);
  and GNAME15536(G15536,G18327,G18328,G18329,G18330);
  and GNAME15537(G15537,G18331,G18332,G18333,G18334);
  and GNAME15538(G15538,G18335,G18336,G18337,G18338);
  and GNAME15539(G15539,G18339,G18340,G18341,G18342);
  and GNAME15540(G15540,G18343,G18344,G18345,G18346);
  and GNAME15541(G15541,G18347,G18348,G18349,G18350);
  and GNAME15542(G15542,G18351,G18352,G18353,G18354);
  and GNAME15543(G15543,G18355,G18356,G18357,G18358);
  and GNAME15544(G15544,G18359,G18360,G18361,G18362);
  and GNAME15545(G15545,G18363,G18364,G18365,G18366);
  and GNAME15546(G15546,G18367,G18368,G18369,G18370);
  and GNAME15547(G15547,G18371,G18372,G18373,G18374);
  and GNAME15548(G15548,G18375,G18376,G18377,G18378);
  and GNAME15549(G15549,G18379,G18380,G18381,G18382);
  and GNAME15550(G15550,G18383,G18384,G18385,G18386);
  and GNAME15551(G15551,G18387,G18388,G18389,G18390);
  and GNAME15552(G15552,G18391,G18392,G18393,G18394);
  and GNAME15553(G15553,G18395,G18396,G18397,G18398);
  and GNAME15554(G15554,G18399,G18400,G18401,G18402);
  and GNAME15555(G15555,G18403,G18404,G18405,G18406);
  and GNAME15556(G15556,G18407,G18408,G18409,G18410);
  and GNAME15557(G15557,G18411,G18412,G18413,G18414);
  and GNAME15558(G15558,G18415,G18416,G18417,G18418);
  and GNAME15559(G15559,G18419,G18420,G18421,G18422);
  and GNAME15560(G15560,G18423,G18424,G18425,G18426);
  and GNAME15561(G15561,G18427,G18428,G18429,G18430);
  and GNAME15562(G15562,G18432,G18433,G18434,G18435);
  and GNAME15563(G15563,G18436,G18437,G18438,G18439);
  and GNAME15564(G15564,G18440,G18441,G18442,G18443);
  and GNAME15565(G15565,G18444,G18445,G18446,G18447);
  and GNAME15566(G15566,G18448,G18449,G18450,G18451);
  and GNAME15567(G15567,G18452,G18453,G18454,G18455);
  and GNAME15568(G15568,G18456,G18457,G18458,G18459);
  and GNAME15569(G15569,G18460,G18461,G18462,G18463);
  and GNAME15570(G15570,G18464,G18465,G18466,G18467);
  and GNAME15571(G15571,G18468,G18469,G18470,G18471);
  and GNAME15572(G15572,G18472,G18473,G18474,G18475);
  and GNAME15573(G15573,G18476,G18477,G18478,G18479);
  and GNAME15574(G15574,G18480,G18481,G18482,G18483);
  and GNAME15575(G15575,G18484,G18485,G18486,G18487);
  and GNAME15576(G15576,G18488,G18489,G18490,G18491);
  and GNAME15577(G15577,G18492,G18493,G18494,G18495);
  and GNAME15578(G15578,G18496,G18497,G18498,G18499);
  and GNAME15579(G15579,G18500,G18501,G18502,G18503);
  and GNAME15580(G15580,G18504,G18505,G18506,G18507);
  and GNAME15581(G15581,G18508,G18509,G18510,G18511);
  and GNAME15582(G15582,G18512,G18513,G18514,G18515);
  and GNAME15583(G15583,G18516,G18517,G18518,G18519);
  and GNAME15584(G15584,G18520,G18521,G18522,G18523);
  and GNAME15585(G15585,G18524,G18525,G18526,G18527);
  and GNAME15586(G15586,G18528,G18529,G18530,G18531);
  and GNAME15587(G15587,G18532,G18533,G18534,G18535);
  and GNAME15588(G15588,G18536,G18537,G18538,G18539);
  and GNAME15589(G15589,G18540,G18541,G18542,G18543);
  and GNAME15590(G15590,G18544,G18545,G18546,G18547);
  and GNAME15591(G15591,G18548,G18549,G18550,G18551);
  and GNAME15592(G15592,G18552,G18553,G18554,G18555);
  and GNAME15593(G15593,G18556,G18557,G18558,G18559);
  and GNAME15594(G15594,G18560,G18561,G18562,G18563);
  and GNAME15595(G15595,G18564,G18565,G18566,G18567);
  and GNAME15596(G15596,G18568,G18569,G18570,G18571);
  and GNAME15597(G15597,G18572,G18573,G18574,G18575);
  and GNAME15598(G15598,G18577,G18578,G18579,G18580);
  and GNAME15599(G15599,G18581,G18582,G18583,G18584);
  and GNAME15600(G15600,G18585,G18586,G18587,G18588);
  and GNAME15601(G15601,G18589,G18590,G18591,G18592);
  and GNAME15602(G15602,G18594,G18595,G18596,G18597);
  and GNAME15603(G15603,G18598,G18599,G18600,G18601);
  and GNAME15604(G15604,G18602,G18603,G18604,G18605);
  and GNAME15605(G15605,G18606,G18607,G18608,G18609);
  and GNAME15606(G15606,G18611,G18612,G18613,G18614);
  and GNAME15607(G15607,G18615,G18616,G18617,G18618);
  and GNAME15608(G15608,G18619,G18620,G18621,G18622);
  and GNAME15609(G15609,G18623,G18624,G18625,G18626);
  and GNAME15610(G15610,G18628,G18629,G18630,G18631);
  and GNAME15611(G15611,G18632,G18633,G18634,G18635);
  and GNAME15612(G15612,G18636,G18637,G18638,G18639);
  and GNAME15613(G15613,G18640,G18641,G18642,G18643);
  and GNAME15614(G15614,G18645,G18646,G18647,G18648);
  and GNAME15615(G15615,G18649,G18650,G18651,G18652);
  and GNAME15616(G15616,G18653,G18654,G18655,G18656);
  and GNAME15617(G15617,G18657,G18658,G18659,G18660);
  and GNAME15618(G15618,G18662,G18663,G18664,G18665);
  and GNAME15619(G15619,G18666,G18667,G18668,G18669);
  and GNAME15620(G15620,G18670,G18671,G18672,G18673);
  and GNAME15621(G15621,G18674,G18675,G18676,G18677);
  and GNAME15622(G15622,G18679,G18680,G18681,G18682);
  and GNAME15623(G15623,G18683,G18684,G18685,G18686);
  and GNAME15624(G15624,G18687,G18688,G18689,G18690);
  and GNAME15625(G15625,G18691,G18692,G18693,G18694);
  and GNAME15626(G15626,G18696,G18697,G18698,G18699);
  and GNAME15627(G15627,G18700,G18701,G18702,G18703);
  and GNAME15628(G15628,G18704,G18705,G18706,G18707);
  and GNAME15629(G15629,G18708,G18709,G18710,G18711);
  and GNAME15630(G15630,G18713,G18714,G18715,G18716);
  and GNAME15631(G15631,G18717,G18718,G18719,G18720);
  and GNAME15632(G15632,G18721,G18722,G18723,G18724);
  and GNAME15633(G15633,G18725,G18726,G18727,G18728);
  and GNAME15634(G15634,G18730,G18731,G18732,G18733);
  and GNAME15635(G15635,G18734,G18735,G18736,G18737);
  and GNAME15636(G15636,G18738,G18739,G18740,G18741);
  and GNAME15637(G15637,G18742,G18743,G18744,G18745);
  and GNAME15638(G15638,G18747,G18748,G18749,G18750);
  and GNAME15639(G15639,G18751,G18752,G18753,G18754);
  and GNAME15640(G15640,G18755,G18756,G18757,G18758);
  and GNAME15641(G15641,G18759,G18760,G18761,G18762);
  and GNAME15642(G15642,G18764,G18765,G18766,G18767);
  and GNAME15643(G15643,G18768,G18769,G18770,G18771);
  and GNAME15644(G15644,G18772,G18773,G18774,G18775);
  and GNAME15645(G15645,G18776,G18777,G18778,G18779);
  and GNAME15646(G15646,G18781,G18782,G18783,G18784);
  and GNAME15647(G15647,G18785,G18786,G18787,G18788);
  and GNAME15648(G15648,G18789,G18790,G18791,G18792);
  and GNAME15649(G15649,G18793,G18794,G18795,G18796);
  and GNAME15650(G15650,G18798,G18799,G18800,G18801);
  and GNAME15651(G15651,G18802,G18803,G18804,G18805);
  and GNAME15652(G15652,G18806,G18807,G18808,G18809);
  and GNAME15653(G15653,G18810,G18811,G18812,G18813);
  and GNAME15654(G15654,G18815,G18816,G18817,G18818);
  and GNAME15655(G15655,G18819,G18820,G18821,G18822);
  and GNAME15656(G15656,G18823,G18824,G18825,G18826);
  and GNAME15657(G15657,G18827,G18828,G18829,G18830);
  and GNAME15658(G15658,G15880,G18991,G18992);
  and GNAME15659(G15659,G19027,G19028,G19029,G19030);
  and GNAME15660(G15660,G19031,G19032,G19033,G19034);
  and GNAME15661(G15661,G19035,G19036,G19037,G19038);
  and GNAME15662(G15662,G19039,G19040,G19041,G19042);
  and GNAME15663(G15663,G19010,G19011,G19012,G19013);
  and GNAME15664(G15664,G19014,G19015,G19016,G19017);
  and GNAME15665(G15665,G19018,G19019,G19020,G19021);
  and GNAME15666(G15666,G19022,G19023,G19024,G19025);
  and GNAME15667(G15667,G18993,G18994,G18995,G18996);
  and GNAME15668(G15668,G18997,G18998,G18999,G19000);
  and GNAME15669(G15669,G19001,G19002,G19003,G19004);
  and GNAME15670(G15670,G19005,G19006,G19007,G19008);
  and GNAME15671(G15671,G19082,G19083,G19084,G19085);
  and GNAME15672(G15672,G19086,G19087,G19088,G19089);
  and GNAME15673(G15673,G19090,G19091,G19092,G19093);
  and GNAME15674(G15674,G19094,G19095,G19096,G19097);
  and GNAME15675(G15675,G19065,G19066,G19067,G19068);
  and GNAME15676(G15676,G19069,G19070,G19071,G19072);
  and GNAME15677(G15677,G19073,G19074,G19075,G19076);
  and GNAME15678(G15678,G19077,G19078,G19079,G19080);
  and GNAME15679(G15679,G19048,G19049,G19050,G19051);
  and GNAME15680(G15680,G19052,G19053,G19054,G19055);
  and GNAME15681(G15681,G19056,G19057,G19058,G19059);
  and GNAME15682(G15682,G19060,G19061,G19062,G19063);
  and GNAME15683(G15683,G19137,G19138,G19139,G19140);
  and GNAME15684(G15684,G19141,G19142,G19143,G19144);
  and GNAME15685(G15685,G19145,G19146,G19147,G19148);
  and GNAME15686(G15686,G19149,G19150,G19151,G19152);
  and GNAME15687(G15687,G19120,G19121,G19122,G19123);
  and GNAME15688(G15688,G19124,G19125,G19126,G19127);
  and GNAME15689(G15689,G19128,G19129,G19130,G19131);
  and GNAME15690(G15690,G19132,G19133,G19134,G19135);
  and GNAME15691(G15691,G19103,G19104,G19105,G19106);
  and GNAME15692(G15692,G19107,G19108,G19109,G19110);
  and GNAME15693(G15693,G19111,G19112,G19113,G19114);
  and GNAME15694(G15694,G19115,G19116,G19117,G19118);
  and GNAME15695(G15695,G19192,G19193,G19194,G19195);
  and GNAME15696(G15696,G19196,G19197,G19198,G19199);
  and GNAME15697(G15697,G19200,G19201,G19202,G19203);
  and GNAME15698(G15698,G19204,G19205,G19206,G19207);
  and GNAME15699(G15699,G19175,G19176,G19177,G19178);
  and GNAME15700(G15700,G19179,G19180,G19181,G19182);
  and GNAME15701(G15701,G19183,G19184,G19185,G19186);
  and GNAME15702(G15702,G19187,G19188,G19189,G19190);
  and GNAME15703(G15703,G19158,G19159,G19160,G19161);
  and GNAME15704(G15704,G19162,G19163,G19164,G19165);
  and GNAME15705(G15705,G19166,G19167,G19168,G19169);
  and GNAME15706(G15706,G19170,G19171,G19172,G19173);
  and GNAME15707(G15707,G19248,G19249,G19250,G19251);
  and GNAME15708(G15708,G19252,G19253,G19254,G19255);
  and GNAME15709(G15709,G19256,G19257,G19258,G19259);
  and GNAME15710(G15710,G19260,G19261,G19262,G19263);
  and GNAME15711(G15711,G19231,G19232,G19233,G19234);
  and GNAME15712(G15712,G19235,G19236,G19237,G19238);
  and GNAME15713(G15713,G19239,G19240,G19241,G19242);
  and GNAME15714(G15714,G19243,G19244,G19245,G19246);
  and GNAME15715(G15715,G19214,G19215,G19216,G19217);
  and GNAME15716(G15716,G19218,G19219,G19220,G19221);
  and GNAME15717(G15717,G19222,G19223,G19224,G19225);
  and GNAME15718(G15718,G19226,G19227,G19228,G19229);
  and GNAME15719(G15719,G19304,G19305,G19306,G19307);
  and GNAME15720(G15720,G19308,G19309,G19310,G19311);
  and GNAME15721(G15721,G19312,G19313,G19314,G19315);
  and GNAME15722(G15722,G19316,G19317,G19318,G19319);
  and GNAME15723(G15723,G19287,G19288,G19289,G19290);
  and GNAME15724(G15724,G19291,G19292,G19293,G19294);
  and GNAME15725(G15725,G19295,G19296,G19297,G19298);
  and GNAME15726(G15726,G19299,G19300,G19301,G19302);
  and GNAME15727(G15727,G19270,G19271,G19272,G19273);
  and GNAME15728(G15728,G19274,G19275,G19276,G19277);
  and GNAME15729(G15729,G19278,G19279,G19280,G19281);
  and GNAME15730(G15730,G19282,G19283,G19284,G19285);
  and GNAME15731(G15731,G19325,G19323,G19324);
  and GNAME15732(G15732,G19360,G19361,G19362,G19363);
  and GNAME15733(G15733,G19364,G19365,G19366,G19367);
  and GNAME15734(G15734,G19368,G19369,G19370,G19371);
  and GNAME15735(G15735,G19372,G19373,G19374,G19375);
  and GNAME15736(G15736,G19343,G19344,G19345,G19346);
  and GNAME15737(G15737,G19347,G19348,G19349,G19350);
  and GNAME15738(G15738,G19351,G19352,G19353,G19354);
  and GNAME15739(G15739,G19355,G19356,G19357,G19358);
  and GNAME15740(G15740,G19326,G19327,G19328,G19329);
  and GNAME15741(G15741,G19330,G19331,G19332,G19333);
  and GNAME15742(G15742,G19334,G19335,G19336,G19337);
  and GNAME15743(G15743,G19338,G19339,G19340,G19341);
  and GNAME15744(G15744,G19381,G19379,G19380);
  and GNAME15745(G15745,G19416,G19417,G19418,G19419);
  and GNAME15746(G15746,G19420,G19421,G19422,G19423);
  and GNAME15747(G15747,G19424,G19425,G19426,G19427);
  and GNAME15748(G15748,G19428,G19429,G19430,G19431);
  and GNAME15749(G15749,G19399,G19400,G19401,G19402);
  and GNAME15750(G15750,G19403,G19404,G19405,G19406);
  and GNAME15751(G15751,G19407,G19408,G19409,G19410);
  and GNAME15752(G15752,G19411,G19412,G19413,G19414);
  and GNAME15753(G15753,G19382,G19383,G19384,G19385);
  and GNAME15754(G15754,G19386,G19387,G19388,G19389);
  and GNAME15755(G15755,G19390,G19391,G19392,G19393);
  and GNAME15756(G15756,G19394,G19395,G19396,G19397);
  and GNAME15757(G15757,G19437,G19435,G19436);
  and GNAME15758(G15758,G19441,G19442);
  and GNAME15759(G15759,G15812,G14849,G19444,G19963);
  and GNAME15760(G15760,G19457,G19455,G19456);
  and GNAME15761(G15761,G19615,G19613,G19614);
  and GNAME15762(G15762,G19666,G19667,G19671,G19668,G19664);
  and GNAME15763(G15763,G19725,G19726,G19730,G19727,G19723);
  and GNAME15764(G15764,G19784,G19785,G19789,G19786,G19782);
  and GNAME15765(G15765,G19793,G19794,G19798,G19795,G19791);
  or GNAME15766(G15766,G14807,G14800);
  and GNAME15767(G15767,G19977,G15969,G15971);
  not GNAME15768(G15768,G35);
  or GNAME15769(G15769,G14921,G14922);
  and GNAME15770(G15770,G17070,G17068,G17069);
  nand GNAME15771(G15771,G17082,G15810,G14906);
  nand GNAME15772(G15772,G17084,G59875);
  and GNAME15773(G15773,G14756,G15863);
  nand GNAME15774(G15774,G14756,G19892);
  nand GNAME15775(G15775,G14885,G17080,G17081);
  not GNAME15776(G15776,G14853);
  not GNAME15777(G15777,G15240);
  not GNAME15778(G15778,G14740);
  not GNAME15779(G15779,G14742);
  not GNAME15780(G15780,G14781);
  not GNAME15781(G15781,G14808);
  not GNAME15782(G15782,G15108);
  not GNAME15783(G15783,G15109);
  not GNAME15784(G15784,G14756);
  not GNAME15785(G15785,G14766);
  not GNAME15786(G15786,G14821);
  not GNAME15787(G15787,G14824);
  not GNAME15788(G15788,G14823);
  not GNAME15789(G15789,G14825);
  not GNAME15790(G15790,G14822);
  not GNAME15791(G15791,G14904);
  not GNAME15792(G15792,G14937);
  not GNAME15793(G15793,G14830);
  not GNAME15794(G15794,G14799);
  not GNAME15795(G15795,G14787);
  not GNAME15796(G15796,G14810);
  nand GNAME15797(G15797,G14907,G14830);
  not GNAME15798(G15798,G14916);
  not GNAME15799(G15799,G14817);
  not GNAME15800(G15800,G14884);
  not GNAME15801(G15801,G14797);
  not GNAME15802(G15802,G14850);
  not GNAME15803(G15803,G14936);
  nand GNAME15804(G15804,G15235,G14793,G23088);
  or GNAME15805(G15805,G59842,G59843,G60207,G19982);
  nand GNAME15806(G15806,G14894,G15973,G59877);
  nand GNAME15807(G15807,G1589,G14836);
  nand GNAME15808(G15808,G14830,G14748,G14784);
  nand GNAME15809(G15809,G59874,G59877,G14799);
  nand GNAME15810(G15810,G60244,G14905);
  nand GNAME15811(G15811,G14814,G14809);
  not GNAME15812(G15812,G14891);
  nand GNAME15813(G15813,G59992,G14752);
  nand GNAME15814(G15814,G59984,G14755);
  nand GNAME15815(G15815,G59976,G14757);
  nand GNAME15816(G15816,G59968,G14761);
  nand GNAME15817(G15817,G59960,G14762);
  nand GNAME15818(G15818,G59952,G14763);
  nand GNAME15819(G15819,G59944,G14764);
  nand GNAME15820(G15820,G59936,G14767);
  nand GNAME15821(G15821,G59928,G14768);
  nand GNAME15822(G15822,G59920,G14769);
  nand GNAME15823(G15823,G59912,G14770);
  nand GNAME15824(G15824,G59904,G14772);
  nand GNAME15825(G15825,G59896,G14773);
  nand GNAME15826(G15826,G59888,G14774);
  nand GNAME15827(G15827,G59880,G14775);
  nand GNAME15828(G15828,G14776,G60000);
  not GNAME15829(G15829,G14777);
  nand GNAME15830(G15830,G14776,G60004);
  nand GNAME15831(G15831,G14752,G59996);
  nand GNAME15832(G15832,G14755,G59988);
  nand GNAME15833(G15833,G14757,G59980);
  nand GNAME15834(G15834,G14761,G59972);
  nand GNAME15835(G15835,G14762,G59964);
  nand GNAME15836(G15836,G14763,G59956);
  nand GNAME15837(G15837,G14764,G59948);
  nand GNAME15838(G15838,G14767,G59940);
  nand GNAME15839(G15839,G14768,G59932);
  nand GNAME15840(G15840,G14769,G59924);
  nand GNAME15841(G15841,G14770,G59916);
  nand GNAME15842(G15842,G14772,G59908);
  nand GNAME15843(G15843,G14773,G59900);
  nand GNAME15844(G15844,G14774,G59892);
  nand GNAME15845(G15845,G14775,G59884);
  not GNAME15846(G15846,G14793);
  nand GNAME15847(G15847,G14776,G60005);
  nand GNAME15848(G15848,G14752,G59997);
  nand GNAME15849(G15849,G14755,G59989);
  nand GNAME15850(G15850,G14757,G59981);
  nand GNAME15851(G15851,G14761,G59973);
  nand GNAME15852(G15852,G14762,G59965);
  nand GNAME15853(G15853,G14763,G59957);
  nand GNAME15854(G15854,G14764,G59949);
  nand GNAME15855(G15855,G14767,G59941);
  nand GNAME15856(G15856,G14768,G59933);
  nand GNAME15857(G15857,G14769,G59925);
  nand GNAME15858(G15858,G14770,G59917);
  nand GNAME15859(G15859,G14772,G59909);
  nand GNAME15860(G15860,G14773,G59901);
  nand GNAME15861(G15861,G14774,G59893);
  nand GNAME15862(G15862,G14775,G59885);
  not GNAME15863(G15863,G14789);
  nand GNAME15864(G15864,G14776,G60003);
  nand GNAME15865(G15865,G14752,G59995);
  nand GNAME15866(G15866,G14755,G59987);
  nand GNAME15867(G15867,G14757,G59979);
  nand GNAME15868(G15868,G14761,G59971);
  nand GNAME15869(G15869,G14762,G59963);
  nand GNAME15870(G15870,G14763,G59955);
  nand GNAME15871(G15871,G14764,G59947);
  nand GNAME15872(G15872,G14767,G59939);
  nand GNAME15873(G15873,G14768,G59931);
  nand GNAME15874(G15874,G14769,G59923);
  nand GNAME15875(G15875,G14770,G59915);
  nand GNAME15876(G15876,G14772,G59907);
  nand GNAME15877(G15877,G14773,G59899);
  nand GNAME15878(G15878,G14774,G59891);
  nand GNAME15879(G15879,G14775,G59883);
  not GNAME15880(G15880,G14778);
  nand GNAME15881(G15881,G14752,G59993);
  nand GNAME15882(G15882,G14755,G59985);
  nand GNAME15883(G15883,G14757,G59977);
  nand GNAME15884(G15884,G14761,G59969);
  nand GNAME15885(G15885,G14762,G59961);
  nand GNAME15886(G15886,G14763,G59953);
  nand GNAME15887(G15887,G14764,G59945);
  nand GNAME15888(G15888,G14767,G59937);
  nand GNAME15889(G15889,G14768,G59929);
  nand GNAME15890(G15890,G14769,G59921);
  nand GNAME15891(G15891,G14770,G59913);
  nand GNAME15892(G15892,G14772,G59905);
  nand GNAME15893(G15893,G14773,G59897);
  nand GNAME15894(G15894,G14774,G59889);
  nand GNAME15895(G15895,G14775,G59881);
  nand GNAME15896(G15896,G14776,G60001);
  not GNAME15897(G15897,G14780);
  nand GNAME15898(G15898,G14752,G59991);
  nand GNAME15899(G15899,G14755,G59983);
  nand GNAME15900(G15900,G14757,G59975);
  nand GNAME15901(G15901,G14761,G59967);
  nand GNAME15902(G15902,G14762,G59959);
  nand GNAME15903(G15903,G14763,G59951);
  nand GNAME15904(G15904,G14764,G59943);
  nand GNAME15905(G15905,G14767,G59935);
  nand GNAME15906(G15906,G14768,G59927);
  nand GNAME15907(G15907,G14769,G59919);
  nand GNAME15908(G15908,G14770,G59911);
  nand GNAME15909(G15909,G14772,G59903);
  nand GNAME15910(G15910,G14773,G59895);
  nand GNAME15911(G15911,G14774,G59887);
  nand GNAME15912(G15912,G14775,G59879);
  nand GNAME15913(G15913,G14776,G59999);
  not GNAME15914(G15914,G14779);
  nand GNAME15915(G15915,G14752,G59990);
  nand GNAME15916(G15916,G14755,G59982);
  nand GNAME15917(G15917,G14757,G59974);
  nand GNAME15918(G15918,G14761,G59966);
  nand GNAME15919(G15919,G14762,G59958);
  nand GNAME15920(G15920,G14763,G59950);
  nand GNAME15921(G15921,G14764,G59942);
  nand GNAME15922(G15922,G14767,G59934);
  nand GNAME15923(G15923,G14768,G59926);
  nand GNAME15924(G15924,G14769,G59918);
  nand GNAME15925(G15925,G14770,G59910);
  nand GNAME15926(G15926,G14772,G59902);
  nand GNAME15927(G15927,G14773,G59894);
  nand GNAME15928(G15928,G14774,G59886);
  nand GNAME15929(G15929,G14775,G59878);
  nand GNAME15930(G15930,G14776,G59998);
  not GNAME15931(G15931,G14849);
  nand GNAME15932(G15932,G14752,G59994);
  nand GNAME15933(G15933,G14755,G59986);
  nand GNAME15934(G15934,G14757,G59978);
  nand GNAME15935(G15935,G14761,G59970);
  nand GNAME15936(G15936,G14762,G59962);
  nand GNAME15937(G15937,G14763,G59954);
  nand GNAME15938(G15938,G14764,G59946);
  nand GNAME15939(G15939,G14767,G59938);
  nand GNAME15940(G15940,G14768,G59930);
  nand GNAME15941(G15941,G14769,G59922);
  nand GNAME15942(G15942,G14770,G59914);
  nand GNAME15943(G15943,G14772,G59906);
  nand GNAME15944(G15944,G14773,G59898);
  nand GNAME15945(G15945,G14774,G59890);
  nand GNAME15946(G15946,G14775,G59882);
  nand GNAME15947(G15947,G14776,G60002);
  not GNAME15948(G15948,G14743);
  not GNAME15949(G15949,G14783);
  not GNAME15950(G15950,G14785);
  nand GNAME15951(G15951,G14792,G59875,G19983);
  not GNAME15952(G15952,G14796);
  nand GNAME15953(G15953,G15951,G14874);
  nand GNAME15954(G15954,G15953,G23088);
  nand GNAME15955(G15955,G59875,G15863);
  or GNAME15956(G15956,G14748,G14740,G14782);
  nor GNAME15957(G15957,G14802,G14803);
  not GNAME15958(G15958,G14804);
  nand GNAME15959(G15959,G59841,G60251);
  nand GNAME15960(G15960,G14790,G15948,G15863);
  nand GNAME15961(G15961,G15960,G14778);
  nand GNAME15962(G15962,G14786,G14793);
  nand GNAME15963(G15963,G14781,G15962,G15829);
  nand GNAME15964(G15964,G14798,G19843);
  nand GNAME15965(G15965,G15963,G15880);
  nand GNAME15966(G15966,G14797,G14806);
  nand GNAME15967(G15967,G15966,G60250);
  nand GNAME15968(G15968,G59877,G14807);
  or GNAME15969(G15969,G1589,G14812);
  nand GNAME15970(G15970,G59875,G59877);
  nand GNAME15971(G15971,G15970,G14813);
  nand GNAME15972(G15972,G14801,G59839);
  nand GNAME15973(G15973,G15972,G14802);
  not GNAME15974(G15974,G14815);
  nand GNAME15975(G15975,G14815,G15863);
  nand GNAME15976(G15976,G14793,G15975);
  nand GNAME15977(G15977,G15974,G60246);
  nand GNAME15978(G15978,G15976,G15977);
  nand GNAME15979(G15979,G15978,G59875);
  nand GNAME15980(G15980,G15863,G14817);
  nand GNAME15981(G15981,G15979,G15980);
  nand GNAME15982(G15982,G14746,G15981);
  nand GNAME15983(G15983,G15982,G59877);
  and GNAME15984(G15984,G15794,G15983);
  nand GNAME15985(G15985,G14815,G19844);
  nand GNAME15986(G15986,G14746,G15985);
  or GNAME15987(G15987,G15101,G15801);
  not GNAME15988(G15988,G14861);
  nand GNAME15989(G15989,G15988,G15776);
  nand GNAME15990(G15990,G15989,G14787);
  nand GNAME15991(G15991,G15990,G15951,G14874);
  nand GNAME15992(G15992,G14819,G59875,G14792);
  nand GNAME15993(G15993,G14785,G14787);
  nand GNAME15994(G15994,G15992,G15993);
  nand GNAME15995(G15995,G14786,G15994);
  nand GNAME15996(G15996,G14798,G15991);
  and GNAME15997(G15997,G15995,G15996);
  or GNAME15998(G15998,G15101,G15997);
  nand GNAME15999(G15999,G15987,G60245);
  nand GNAME16000(G16000,G59875,G23753,G14792,G14819);
  nand GNAME16001(G16001,G15987,G60244);
  and GNAME16002(G16002,G59843,G59842);
  nand GNAME16003(G16003,G19982,G60241);
  and GNAME16004(G16004,G59842,G60207);
  or GNAME16005(G16005,G16004,G14828);
  or GNAME16006(G16006,G14827,G14829);
  nand GNAME16007(G16007,G19982,G60240);
  nand GNAME16008(G16008,G19982,G60239);
  not GNAME16009(G16009,G14839);
  not GNAME16010(G16010,G14832);
  nand GNAME16011(G16011,G14833,G14824,G14832);
  nand GNAME16012(G16012,G23190,G14839,G59876);
  nand GNAME16013(G16013,G16010,G14824,G14833,G15279);
  or GNAME16014(G16014,G14811,G23190,G16009);
  nand GNAME16015(G16015,G16013,G16014);
  nand GNAME16016(G16016,G15974,G14832);
  nand GNAME16017(G16017,G14824,G14835,G16010);
  nand GNAME16018(G16018,G16016,G14794);
  nand GNAME16019(G16019,G16017,G16018);
  nand GNAME16020(G16020,G14834,G60206);
  nand GNAME16021(G16021,G16015,G23190);
  nand GNAME16022(G16022,G60079,G14837);
  nand GNAME16023(G16023,G14840,G23488);
  nand GNAME16024(G16024,G23901,G14838);
  nand GNAME16025(G16025,G16009,G60238);
  nand GNAME16026(G16026,G14834,G60205);
  nand GNAME16027(G16027,G16015,G23122);
  nand GNAME16028(G16028,G14837,G60078);
  nand GNAME16029(G16029,G14840,G23427);
  nand GNAME16030(G16030,G14838,G23902);
  nand GNAME16031(G16031,G16009,G60237);
  nand GNAME16032(G16032,G14834,G60204);
  nand GNAME16033(G16033,G16015,G23176);
  nand GNAME16034(G16034,G14837,G60077);
  nand GNAME16035(G16035,G14840,G23475);
  nand GNAME16036(G16036,G14838,G23940);
  nand GNAME16037(G16037,G16009,G60236);
  nand GNAME16038(G16038,G14834,G60203);
  nand GNAME16039(G16039,G16015,G23177);
  nand GNAME16040(G16040,G14837,G60076);
  nand GNAME16041(G16041,G14840,G23476);
  nand GNAME16042(G16042,G14838,G23941);
  nand GNAME16043(G16043,G16009,G60235);
  nand GNAME16044(G16044,G14834,G60202);
  nand GNAME16045(G16045,G16015,G23178);
  nand GNAME16046(G16046,G14837,G60075);
  nand GNAME16047(G16047,G14840,G23477);
  nand GNAME16048(G16048,G14838,G23942);
  nand GNAME16049(G16049,G16009,G60234);
  nand GNAME16050(G16050,G14834,G60201);
  nand GNAME16051(G16051,G16015,G23179);
  nand GNAME16052(G16052,G14837,G60074);
  nand GNAME16053(G16053,G14840,G23478);
  nand GNAME16054(G16054,G14838,G23943);
  nand GNAME16055(G16055,G16009,G60233);
  nand GNAME16056(G16056,G14834,G60200);
  nand GNAME16057(G16057,G16015,G23180);
  nand GNAME16058(G16058,G14837,G60073);
  nand GNAME16059(G16059,G14840,G23479);
  nand GNAME16060(G16060,G14838,G23944);
  nand GNAME16061(G16061,G16009,G60232);
  nand GNAME16062(G16062,G14834,G60199);
  nand GNAME16063(G16063,G16015,G23181);
  nand GNAME16064(G16064,G14837,G60072);
  nand GNAME16065(G16065,G14840,G23517);
  nand GNAME16066(G16066,G14838,G23945);
  nand GNAME16067(G16067,G16009,G60231);
  nand GNAME16068(G16068,G14834,G60198);
  nand GNAME16069(G16069,G16015,G23182);
  nand GNAME16070(G16070,G14837,G60071);
  nand GNAME16071(G16071,G14840,G23520);
  nand GNAME16072(G16072,G14838,G23946);
  nand GNAME16073(G16073,G16009,G60230);
  nand GNAME16074(G16074,G14834,G60197);
  nand GNAME16075(G16075,G16015,G23183);
  nand GNAME16076(G16076,G14837,G60070);
  nand GNAME16077(G16077,G14840,G23523);
  nand GNAME16078(G16078,G14838,G23947);
  nand GNAME16079(G16079,G16009,G60229);
  nand GNAME16080(G16080,G14834,G60196);
  nand GNAME16081(G16081,G16015,G23184);
  nand GNAME16082(G16082,G14837,G60069);
  nand GNAME16083(G16083,G14840,G23526);
  nand GNAME16084(G16084,G14838,G23948);
  nand GNAME16085(G16085,G16009,G60228);
  nand GNAME16086(G16086,G14834,G60195);
  nand GNAME16087(G16087,G16015,G23185);
  nand GNAME16088(G16088,G14837,G60068);
  nand GNAME16089(G16089,G14840,G23529);
  nand GNAME16090(G16090,G14838,G23949);
  nand GNAME16091(G16091,G16009,G60227);
  nand GNAME16092(G16092,G14839,G14784,G14811);
  nand GNAME16093(G16093,G14834,G60194);
  nand GNAME16094(G16094,G16015,G23186);
  nand GNAME16095(G16095,G14837,G60067);
  nand GNAME16096(G16096,G14840,G23535);
  nand GNAME16097(G16097,G14838,G23953);
  nand GNAME16098(G16098,G16009,G60226);
  nand GNAME16099(G16099,G14834,G60193);
  nand GNAME16100(G16100,G16015,G23187);
  nand GNAME16101(G16101,G14837,G60066);
  nand GNAME16102(G16102,G14840,G23538);
  nand GNAME16103(G16103,G14838,G23954);
  nand GNAME16104(G16104,G16009,G60225);
  nand GNAME16105(G16105,G14834,G60192);
  nand GNAME16106(G16106,G16015,G23188);
  nand GNAME16107(G16107,G14837,G60065);
  nand GNAME16108(G16108,G14840,G23541);
  nand GNAME16109(G16109,G14838,G23955);
  nand GNAME16110(G16110,G16009,G60224);
  nand GNAME16111(G16111,G14834,G60191);
  nand GNAME16112(G16112,G16015,G23216);
  nand GNAME16113(G16113,G14837,G60064);
  nand GNAME16114(G16114,G14840,G23480);
  nand GNAME16115(G16115,G14838,G23956);
  nand GNAME16116(G16116,G16009,G60223);
  nand GNAME16117(G16117,G14834,G60190);
  nand GNAME16118(G16118,G16015,G23219);
  nand GNAME16119(G16119,G14837,G60063);
  nand GNAME16120(G16120,G14840,G23481);
  nand GNAME16121(G16121,G14838,G23957);
  nand GNAME16122(G16122,G16009,G60222);
  nand GNAME16123(G16123,G14834,G60189);
  nand GNAME16124(G16124,G16015,G23191);
  nand GNAME16125(G16125,G14837,G60062);
  nand GNAME16126(G16126,G14840,G23425);
  nand GNAME16127(G16127,G14838,G23903);
  nand GNAME16128(G16128,G16009,G60221);
  nand GNAME16129(G16129,G14834,G60188);
  nand GNAME16130(G16130,G16015,G23223);
  nand GNAME16131(G16131,G14837,G60061);
  nand GNAME16132(G16132,G14840,G23482);
  nand GNAME16133(G16133,G14838,G23958);
  nand GNAME16134(G16134,G16009,G60220);
  nand GNAME16135(G16135,G14834,G60187);
  nand GNAME16136(G16136,G16015,G23226);
  nand GNAME16137(G16137,G14837,G60060);
  nand GNAME16138(G16138,G14840,G23483);
  nand GNAME16139(G16139,G14838,G23959);
  nand GNAME16140(G16140,G16009,G60219);
  nand GNAME16141(G16141,G14834,G60186);
  nand GNAME16142(G16142,G16015,G23192);
  nand GNAME16143(G16143,G14837,G60059);
  nand GNAME16144(G16144,G14840,G23484);
  nand GNAME16145(G16145,G14838,G23839);
  nand GNAME16146(G16146,G16009,G60218);
  nand GNAME16147(G16147,G14834,G60185);
  nand GNAME16148(G16148,G16015,G23120);
  nand GNAME16149(G16149,G14837,G60058);
  nand GNAME16150(G16150,G14840,G23424);
  nand GNAME16151(G16151,G14838,G23838);
  nand GNAME16152(G16152,G16009,G60217);
  nand GNAME16153(G16153,G14834,G60184);
  nand GNAME16154(G16154,G16015,G23199);
  nand GNAME16155(G16155,G14837,G60057);
  nand GNAME16156(G16156,G14840,G23461);
  nand GNAME16157(G16157,G14838,G23930);
  nand GNAME16158(G16158,G16009,G60216);
  nand GNAME16159(G16159,G14834,G60183);
  nand GNAME16160(G16160,G16015,G23156);
  nand GNAME16161(G16161,G14837,G60056);
  nand GNAME16162(G16162,G14840,G23496);
  nand GNAME16163(G16163,G14838,G23931);
  nand GNAME16164(G16164,G16009,G60215);
  nand GNAME16165(G16165,G14834,G60182);
  nand GNAME16166(G16166,G16015,G23157);
  nand GNAME16167(G16167,G14837,G60055);
  nand GNAME16168(G16168,G14840,G23486);
  nand GNAME16169(G16169,G14838,G23899);
  nand GNAME16170(G16170,G16009,G60214);
  nand GNAME16171(G16171,G14834,G60181);
  nand GNAME16172(G16172,G16015,G23123);
  nand GNAME16173(G16173,G14837,G60054);
  nand GNAME16174(G16174,G14840,G23428);
  nand GNAME16175(G16175,G14838,G23841);
  nand GNAME16176(G16176,G16009,G60213);
  and GNAME16177(G16177,G14833,G14793,G14779);
  or GNAME16178(G16178,G16177,G14840);
  and GNAME16179(G16179,G14817,G14779,G14839);
  or GNAME16180(G16180,G16179,G14838);
  nand GNAME16181(G16181,G14834,G60180);
  nand GNAME16182(G16182,G16015,G23158);
  nand GNAME16183(G16183,G16180,G23935);
  nand GNAME16184(G16184,G14837,G60053);
  nand GNAME16185(G16185,G16178,G23500);
  nand GNAME16186(G16186,G16009,G60212);
  nand GNAME16187(G16187,G14834,G60179);
  nand GNAME16188(G16188,G16015,G23159);
  nand GNAME16189(G16189,G16180,G23938);
  nand GNAME16190(G16190,G14837,G60052);
  nand GNAME16191(G16191,G16178,G23503);
  nand GNAME16192(G16192,G16009,G60211);
  nand GNAME16193(G16193,G14834,G60178);
  nand GNAME16194(G16194,G16015,G23160);
  nand GNAME16195(G16195,G16180,G23900);
  nand GNAME16196(G16196,G14837,G60051);
  nand GNAME16197(G16197,G16009,G60210);
  nand GNAME16198(G16198,G16178,G23487);
  nand GNAME16199(G16199,G14834,G60177);
  nand GNAME16200(G16200,G16015,G23121);
  nand GNAME16201(G16201,G16180,G23840);
  nand GNAME16202(G16202,G14837,G60050);
  nand GNAME16203(G16203,G16009,G60209);
  nand GNAME16204(G16204,G16178,G23426);
  nand GNAME16205(G16205,G14834,G60176);
  nand GNAME16206(G16206,G16015,G23213);
  nand GNAME16207(G16207,G16180,G23952);
  nand GNAME16208(G16208,G14837,G60049);
  nand GNAME16209(G16209,G16178,G23532);
  nand GNAME16210(G16210,G60208,G16009);
  nand GNAME16211(G16211,G14834,G60175);
  nand GNAME16212(G16212,G16015,G23189);
  nand GNAME16213(G16213,G16180,G23898);
  nand GNAME16214(G16214,G14837,G60048);
  nand GNAME16215(G16215,G16178,G23485);
  nand GNAME16216(G16216,G60207,G16009);
  not GNAME16217(G16217,G14852);
  nand GNAME16218(G16218,G59877,G16217);
  nand GNAME16219(G16219,G23088,G14853);
  nand GNAME16220(G16220,G16218,G16219);
  nand GNAME16221(G16221,G14854,G60206);
  nand GNAME16222(G16222,G23190,G14855);
  nand GNAME16223(G16223,G14854,G60205);
  nand GNAME16224(G16224,G23427,G14856);
  nand GNAME16225(G16225,G23122,G14855);
  nand GNAME16226(G16226,G14854,G60204);
  nand GNAME16227(G16227,G23475,G14856);
  nand GNAME16228(G16228,G23176,G14855);
  nand GNAME16229(G16229,G14854,G60203);
  nand GNAME16230(G16230,G23476,G14856);
  nand GNAME16231(G16231,G23177,G14855);
  nand GNAME16232(G16232,G14854,G60202);
  nand GNAME16233(G16233,G23477,G14856);
  nand GNAME16234(G16234,G23178,G14855);
  nand GNAME16235(G16235,G14854,G60201);
  nand GNAME16236(G16236,G23478,G14856);
  nand GNAME16237(G16237,G23179,G14855);
  nand GNAME16238(G16238,G14854,G60200);
  nand GNAME16239(G16239,G23479,G14856);
  nand GNAME16240(G16240,G23180,G14855);
  nand GNAME16241(G16241,G14854,G60199);
  nand GNAME16242(G16242,G23517,G14856);
  nand GNAME16243(G16243,G23181,G14855);
  nand GNAME16244(G16244,G14854,G60198);
  nand GNAME16245(G16245,G23520,G14856);
  nand GNAME16246(G16246,G23182,G14855);
  nand GNAME16247(G16247,G14854,G60197);
  nand GNAME16248(G16248,G23523,G14856);
  nand GNAME16249(G16249,G23183,G14855);
  nand GNAME16250(G16250,G14854,G60196);
  nand GNAME16251(G16251,G23526,G14856);
  nand GNAME16252(G16252,G23184,G14855);
  nand GNAME16253(G16253,G14854,G60195);
  nand GNAME16254(G16254,G23529,G14856);
  nand GNAME16255(G16255,G23185,G14855);
  nand GNAME16256(G16256,G14854,G60194);
  nand GNAME16257(G16257,G23535,G14856);
  nand GNAME16258(G16258,G23186,G14855);
  nand GNAME16259(G16259,G14854,G60193);
  nand GNAME16260(G16260,G23538,G14856);
  nand GNAME16261(G16261,G23187,G14855);
  nand GNAME16262(G16262,G14854,G60192);
  nand GNAME16263(G16263,G23541,G14856);
  nand GNAME16264(G16264,G23188,G14855);
  nand GNAME16265(G16265,G14854,G60191);
  nand GNAME16266(G16266,G23480,G14856);
  nand GNAME16267(G16267,G23216,G14855);
  nand GNAME16268(G16268,G14854,G60190);
  nand GNAME16269(G16269,G23481,G14856);
  nand GNAME16270(G16270,G23219,G14855);
  nand GNAME16271(G16271,G14854,G60189);
  nand GNAME16272(G16272,G23425,G14856);
  nand GNAME16273(G16273,G23191,G14855);
  nand GNAME16274(G16274,G14854,G60188);
  nand GNAME16275(G16275,G23482,G14856);
  nand GNAME16276(G16276,G23223,G14855);
  nand GNAME16277(G16277,G14854,G60187);
  nand GNAME16278(G16278,G23483,G14856);
  nand GNAME16279(G16279,G23226,G14855);
  nand GNAME16280(G16280,G14854,G60186);
  nand GNAME16281(G16281,G23484,G14856);
  nand GNAME16282(G16282,G23192,G14855);
  nand GNAME16283(G16283,G14854,G60185);
  nand GNAME16284(G16284,G23424,G14856);
  nand GNAME16285(G16285,G23120,G14855);
  nand GNAME16286(G16286,G14854,G60184);
  nand GNAME16287(G16287,G23461,G14856);
  nand GNAME16288(G16288,G23199,G14855);
  nand GNAME16289(G16289,G14854,G60183);
  nand GNAME16290(G16290,G23496,G14856);
  nand GNAME16291(G16291,G23156,G14855);
  nand GNAME16292(G16292,G14854,G60182);
  nand GNAME16293(G16293,G23486,G14856);
  nand GNAME16294(G16294,G23157,G14855);
  nand GNAME16295(G16295,G14854,G60181);
  nand GNAME16296(G16296,G23428,G14856);
  nand GNAME16297(G16297,G23123,G14855);
  nand GNAME16298(G16298,G14854,G60180);
  nand GNAME16299(G16299,G23500,G14856);
  nand GNAME16300(G16300,G23158,G14855);
  nand GNAME16301(G16301,G14854,G60179);
  nand GNAME16302(G16302,G23503,G14856);
  nand GNAME16303(G16303,G23159,G14855);
  nand GNAME16304(G16304,G14854,G60178);
  nand GNAME16305(G16305,G23160,G14855);
  nand GNAME16306(G16306,G23487,G14856);
  nand GNAME16307(G16307,G14854,G60177);
  nand GNAME16308(G16308,G23121,G14855);
  nand GNAME16309(G16309,G23426,G14856);
  nand GNAME16310(G16310,G14854,G60176);
  nand GNAME16311(G16311,G23532,G14856);
  nand GNAME16312(G16312,G23213,G14855);
  nand GNAME16313(G16313,G14854,G60175);
  nand GNAME16314(G16314,G23189,G14855);
  nand GNAME16315(G16315,G23485,G14856);
  not GNAME16316(G16316,G14858);
  not GNAME16317(G16317,G15241);
  not GNAME16318(G16318,G14859);
  or GNAME16319(G16319,G14798,G14860);
  nand GNAME16320(G16320,G14785,G23753);
  nand GNAME16321(G16321,G16319,G16320);
  nand GNAME16322(G16322,G14746,G16321);
  nand GNAME16323(G16323,G23088,G14861);
  nand GNAME16324(G16324,G16323,G16317,G16322);
  nand GNAME16325(G16325,G14862,G60174);
  nand GNAME16326(G16326,G23190,G14863);
  nand GNAME16327(G16327,G14864,G1667);
  nand GNAME16328(G16328,G1686,G14865);
  nand GNAME16329(G16329,G14862,G60173);
  nand GNAME16330(G16330,G23122,G14863);
  nand GNAME16331(G16331,G23902,G14866);
  nand GNAME16332(G16332,G14864,G1668);
  nand GNAME16333(G16333,G14865,G1687);
  nand GNAME16334(G16334,G14862,G60172);
  nand GNAME16335(G16335,G23176,G14863);
  nand GNAME16336(G16336,G23940,G14866);
  nand GNAME16337(G16337,G14864,G1670);
  nand GNAME16338(G16338,G14865,G1688);
  nand GNAME16339(G16339,G14862,G60171);
  nand GNAME16340(G16340,G23177,G14863);
  nand GNAME16341(G16341,G23941,G14866);
  nand GNAME16342(G16342,G14864,G1671);
  nand GNAME16343(G16343,G14865,G1689);
  nand GNAME16344(G16344,G14862,G60170);
  nand GNAME16345(G16345,G23178,G14863);
  nand GNAME16346(G16346,G23942,G14866);
  nand GNAME16347(G16347,G14864,G1672);
  nand GNAME16348(G16348,G14865,G1690);
  nand GNAME16349(G16349,G14862,G60169);
  nand GNAME16350(G16350,G23179,G14863);
  nand GNAME16351(G16351,G23943,G14866);
  nand GNAME16352(G16352,G14864,G1673);
  nand GNAME16353(G16353,G14865,G1660);
  nand GNAME16354(G16354,G14862,G60168);
  nand GNAME16355(G16355,G23180,G14863);
  nand GNAME16356(G16356,G23944,G14866);
  nand GNAME16357(G16357,G14864,G1674);
  nand GNAME16358(G16358,G14865,G1661);
  nand GNAME16359(G16359,G14862,G60167);
  nand GNAME16360(G16360,G23181,G14863);
  nand GNAME16361(G16361,G23945,G14866);
  nand GNAME16362(G16362,G14864,G1675);
  nand GNAME16363(G16363,G14862,G60166);
  nand GNAME16364(G16364,G23182,G14863);
  nand GNAME16365(G16365,G23946,G14866);
  nand GNAME16366(G16366,G14864,G1676);
  nand GNAME16367(G16367,G14865,G1662);
  nand GNAME16368(G16368,G14862,G60165);
  nand GNAME16369(G16369,G23183,G14863);
  nand GNAME16370(G16370,G23947,G14866);
  nand GNAME16371(G16371,G14864,G1677);
  nand GNAME16372(G16372,G14865,G1663);
  nand GNAME16373(G16373,G14862,G60164);
  nand GNAME16374(G16374,G23184,G14863);
  nand GNAME16375(G16375,G23948,G14866);
  nand GNAME16376(G16376,G14864,G1678);
  nand GNAME16377(G16377,G14865,G1664);
  nand GNAME16378(G16378,G14862,G60163);
  nand GNAME16379(G16379,G23185,G14863);
  nand GNAME16380(G16380,G23949,G14866);
  nand GNAME16381(G16381,G14864,G1679);
  nand GNAME16382(G16382,G14865,G1665);
  nand GNAME16383(G16383,G14862,G60162);
  nand GNAME16384(G16384,G23186,G14863);
  nand GNAME16385(G16385,G23953,G14866);
  nand GNAME16386(G16386,G14864,G1681);
  nand GNAME16387(G16387,G14865,G1666);
  nand GNAME16388(G16388,G14862,G60161);
  nand GNAME16389(G16389,G23187,G14863);
  nand GNAME16390(G16390,G23954,G14866);
  nand GNAME16391(G16391,G14864,G1682);
  nand GNAME16392(G16392,G14865,G1669);
  nand GNAME16393(G16393,G14862,G60160);
  nand GNAME16394(G16394,G23188,G14863);
  nand GNAME16395(G16395,G23955,G14866);
  nand GNAME16396(G16396,G14864,G1683);
  nand GNAME16397(G16397,G14865,G1680);
  nand GNAME16398(G16398,G14862,G60159);
  nand GNAME16399(G16399,G23216,G14863);
  nand GNAME16400(G16400,G23956,G14866);
  nand GNAME16401(G16401,G14864,G1684);
  nand GNAME16402(G16402,G14865,G1691);
  nand GNAME16403(G16403,G1685,G14867);
  nand GNAME16404(G16404,G14862,G60158);
  nand GNAME16405(G16405,G23219,G14863);
  nand GNAME16406(G16406,G23957,G14866);
  nand GNAME16407(G16407,G1686,G14867);
  nand GNAME16408(G16408,G14862,G60157);
  nand GNAME16409(G16409,G23191,G14863);
  nand GNAME16410(G16410,G23903,G14866);
  nand GNAME16411(G16411,G1687,G14867);
  nand GNAME16412(G16412,G14862,G60156);
  nand GNAME16413(G16413,G23223,G14863);
  nand GNAME16414(G16414,G23958,G14866);
  nand GNAME16415(G16415,G1688,G14867);
  nand GNAME16416(G16416,G14862,G60155);
  nand GNAME16417(G16417,G23226,G14863);
  nand GNAME16418(G16418,G23959,G14866);
  nand GNAME16419(G16419,G1689,G14867);
  nand GNAME16420(G16420,G14862,G60154);
  nand GNAME16421(G16421,G23192,G14863);
  nand GNAME16422(G16422,G23839,G14866);
  nand GNAME16423(G16423,G1690,G14867);
  nand GNAME16424(G16424,G14862,G60153);
  nand GNAME16425(G16425,G23120,G14863);
  nand GNAME16426(G16426,G23838,G14866);
  nand GNAME16427(G16427,G1660,G14867);
  nand GNAME16428(G16428,G14862,G60152);
  nand GNAME16429(G16429,G23199,G14863);
  nand GNAME16430(G16430,G23930,G14866);
  nand GNAME16431(G16431,G1661,G14867);
  nand GNAME16432(G16432,G14862,G60151);
  nand GNAME16433(G16433,G23156,G14863);
  nand GNAME16434(G16434,G23931,G14866);
  nand GNAME16435(G16435,G14862,G60150);
  nand GNAME16436(G16436,G23157,G14863);
  nand GNAME16437(G16437,G23899,G14866);
  nand GNAME16438(G16438,G1662,G14867);
  nand GNAME16439(G16439,G14862,G60149);
  nand GNAME16440(G16440,G23123,G14863);
  nand GNAME16441(G16441,G23841,G14866);
  nand GNAME16442(G16442,G1663,G14867);
  nand GNAME16443(G16443,G14862,G60148);
  nand GNAME16444(G16444,G23158,G14863);
  nand GNAME16445(G16445,G23935,G14866);
  nand GNAME16446(G16446,G1664,G14867);
  nand GNAME16447(G16447,G14862,G60147);
  nand GNAME16448(G16448,G23159,G14863);
  nand GNAME16449(G16449,G23938,G14866);
  nand GNAME16450(G16450,G1665,G14867);
  nand GNAME16451(G16451,G14862,G60146);
  nand GNAME16452(G16452,G23900,G14866);
  nand GNAME16453(G16453,G23160,G14863);
  nand GNAME16454(G16454,G1666,G14867);
  nand GNAME16455(G16455,G14862,G60145);
  nand GNAME16456(G16456,G23840,G14866);
  nand GNAME16457(G16457,G23121,G14863);
  nand GNAME16458(G16458,G1669,G14867);
  nand GNAME16459(G16459,G14862,G60144);
  nand GNAME16460(G16460,G23952,G14866);
  nand GNAME16461(G16461,G23213,G14863);
  nand GNAME16462(G16462,G1680,G14867);
  nand GNAME16463(G16463,G14862,G60143);
  nand GNAME16464(G16464,G23898,G14866);
  nand GNAME16465(G16465,G23189,G14863);
  nand GNAME16466(G16466,G1691,G14867);
  not GNAME16467(G16467,G14868);
  nand GNAME16468(G16468,G14868,G59877,G15974);
  or GNAME16469(G16469,G59841,G14869);
  nand GNAME16470(G16470,G16468,G16469);
  nand GNAME16471(G16471,G23088,G16470,G14787);
  nand GNAME16472(G16472,G14870,G60141);
  nand GNAME16473(G16473,G60096,G14871);
  nand GNAME16474(G16474,G60173,G14873);
  nand GNAME16475(G16475,G14870,G60140);
  nand GNAME16476(G16476,G14871,G60097);
  nand GNAME16477(G16477,G60172,G14873);
  nand GNAME16478(G16478,G14870,G60139);
  nand GNAME16479(G16479,G14871,G60098);
  nand GNAME16480(G16480,G60171,G14873);
  nand GNAME16481(G16481,G14870,G60138);
  nand GNAME16482(G16482,G14871,G60099);
  nand GNAME16483(G16483,G60170,G14873);
  nand GNAME16484(G16484,G14870,G60137);
  nand GNAME16485(G16485,G14871,G60100);
  nand GNAME16486(G16486,G60169,G14873);
  nand GNAME16487(G16487,G14870,G60136);
  nand GNAME16488(G16488,G14871,G60101);
  nand GNAME16489(G16489,G60168,G14873);
  nand GNAME16490(G16490,G14870,G60135);
  nand GNAME16491(G16491,G14871,G60102);
  nand GNAME16492(G16492,G60167,G14873);
  nand GNAME16493(G16493,G14870,G60134);
  nand GNAME16494(G16494,G14871,G60103);
  nand GNAME16495(G16495,G60166,G14873);
  nand GNAME16496(G16496,G14870,G60133);
  nand GNAME16497(G16497,G14871,G60104);
  nand GNAME16498(G16498,G60165,G14873);
  nand GNAME16499(G16499,G14870,G60132);
  nand GNAME16500(G16500,G14871,G60105);
  nand GNAME16501(G16501,G60164,G14873);
  nand GNAME16502(G16502,G14870,G60131);
  nand GNAME16503(G16503,G14871,G60106);
  nand GNAME16504(G16504,G60163,G14873);
  nand GNAME16505(G16505,G14870,G60130);
  nand GNAME16506(G16506,G14871,G60107);
  nand GNAME16507(G16507,G60162,G14873);
  nand GNAME16508(G16508,G14870,G60129);
  nand GNAME16509(G16509,G14871,G60108);
  nand GNAME16510(G16510,G60161,G14873);
  nand GNAME16511(G16511,G14870,G60128);
  nand GNAME16512(G16512,G14871,G60109);
  nand GNAME16513(G16513,G60160,G14873);
  nand GNAME16514(G16514,G14870,G60127);
  nand GNAME16515(G16515,G14871,G60110);
  nand GNAME16516(G16516,G60159,G14873);
  nand GNAME16517(G16517,G14870,G60126);
  nand GNAME16518(G16518,G14871,G60080);
  nand GNAME16519(G16519,G60158,G14872);
  nand GNAME16520(G16520,G14870,G60125);
  nand GNAME16521(G16521,G14871,G60081);
  nand GNAME16522(G16522,G60157,G14872);
  nand GNAME16523(G16523,G14870,G60124);
  nand GNAME16524(G16524,G14871,G60082);
  nand GNAME16525(G16525,G60156,G14872);
  nand GNAME16526(G16526,G14870,G60123);
  nand GNAME16527(G16527,G14871,G60083);
  nand GNAME16528(G16528,G60155,G14872);
  nand GNAME16529(G16529,G14870,G60122);
  nand GNAME16530(G16530,G14871,G60084);
  nand GNAME16531(G16531,G60154,G14872);
  nand GNAME16532(G16532,G14870,G60121);
  nand GNAME16533(G16533,G14871,G60085);
  nand GNAME16534(G16534,G60153,G14872);
  nand GNAME16535(G16535,G14870,G60120);
  nand GNAME16536(G16536,G14871,G60086);
  nand GNAME16537(G16537,G60152,G14872);
  nand GNAME16538(G16538,G14870,G60119);
  nand GNAME16539(G16539,G14871,G60087);
  nand GNAME16540(G16540,G60151,G14872);
  nand GNAME16541(G16541,G14870,G60118);
  nand GNAME16542(G16542,G14871,G60088);
  nand GNAME16543(G16543,G60150,G14872);
  nand GNAME16544(G16544,G14870,G60117);
  nand GNAME16545(G16545,G14871,G60089);
  nand GNAME16546(G16546,G60149,G14872);
  nand GNAME16547(G16547,G14870,G60116);
  nand GNAME16548(G16548,G14871,G60090);
  nand GNAME16549(G16549,G60148,G14872);
  nand GNAME16550(G16550,G14870,G60115);
  nand GNAME16551(G16551,G14871,G60091);
  nand GNAME16552(G16552,G60147,G14872);
  nand GNAME16553(G16553,G14870,G60114);
  nand GNAME16554(G16554,G14871,G60092);
  nand GNAME16555(G16555,G60146,G14872);
  nand GNAME16556(G16556,G14870,G60113);
  nand GNAME16557(G16557,G14871,G60093);
  nand GNAME16558(G16558,G60145,G14872);
  nand GNAME16559(G16559,G14870,G60112);
  nand GNAME16560(G16560,G14871,G60094);
  nand GNAME16561(G16561,G60144,G14872);
  nand GNAME16562(G16562,G14870,G60111);
  nand GNAME16563(G16563,G14871,G60095);
  nand GNAME16564(G16564,G60143,G14872);
  or GNAME16565(G16565,G14798,G14874);
  or GNAME16566(G16566,G1589,G14875);
  nand GNAME16567(G16567,G60110,G14876);
  nand GNAME16568(G16568,G60159,G14877);
  nand GNAME16569(G16569,G60109,G14876);
  nand GNAME16570(G16570,G60160,G14877);
  nand GNAME16571(G16571,G60108,G14876);
  nand GNAME16572(G16572,G60161,G14877);
  nand GNAME16573(G16573,G60107,G14876);
  nand GNAME16574(G16574,G60162,G14877);
  nand GNAME16575(G16575,G60106,G14876);
  nand GNAME16576(G16576,G60163,G14877);
  nand GNAME16577(G16577,G60105,G14876);
  nand GNAME16578(G16578,G60164,G14877);
  nand GNAME16579(G16579,G60104,G14876);
  nand GNAME16580(G16580,G60165,G14877);
  nand GNAME16581(G16581,G60103,G14876);
  nand GNAME16582(G16582,G60166,G14877);
  nand GNAME16583(G16583,G60102,G14876);
  nand GNAME16584(G16584,G60167,G14877);
  nand GNAME16585(G16585,G60101,G14876);
  nand GNAME16586(G16586,G60168,G14877);
  nand GNAME16587(G16587,G60100,G14876);
  nand GNAME16588(G16588,G60169,G14877);
  nand GNAME16589(G16589,G60099,G14876);
  nand GNAME16590(G16590,G60170,G14877);
  nand GNAME16591(G16591,G60098,G14876);
  nand GNAME16592(G16592,G60171,G14877);
  nand GNAME16593(G16593,G60097,G14876);
  nand GNAME16594(G16594,G60172,G14877);
  nand GNAME16595(G16595,G60096,G14876);
  nand GNAME16596(G16596,G60173,G14877);
  nand GNAME16597(G16597,G60095,G14876);
  nand GNAME16598(G16598,G60143,G14877);
  nand GNAME16599(G16599,G1691,G14878);
  nand GNAME16600(G16600,G60094,G14876);
  nand GNAME16601(G16601,G60144,G14877);
  nand GNAME16602(G16602,G1680,G14878);
  nand GNAME16603(G16603,G60093,G14876);
  nand GNAME16604(G16604,G60145,G14877);
  nand GNAME16605(G16605,G1669,G14878);
  nand GNAME16606(G16606,G60092,G14876);
  nand GNAME16607(G16607,G60146,G14877);
  nand GNAME16608(G16608,G1666,G14878);
  nand GNAME16609(G16609,G60091,G14876);
  nand GNAME16610(G16610,G60147,G14877);
  nand GNAME16611(G16611,G1665,G14878);
  nand GNAME16612(G16612,G60090,G14876);
  nand GNAME16613(G16613,G60148,G14877);
  nand GNAME16614(G16614,G1664,G14878);
  nand GNAME16615(G16615,G60089,G14876);
  nand GNAME16616(G16616,G60149,G14877);
  nand GNAME16617(G16617,G1663,G14878);
  nand GNAME16618(G16618,G60088,G14876);
  nand GNAME16619(G16619,G60150,G14877);
  nand GNAME16620(G16620,G1662,G14878);
  nand GNAME16621(G16621,G1661,G14878);
  nand GNAME16622(G16622,G60087,G14876);
  nand GNAME16623(G16623,G60151,G14877);
  nand GNAME16624(G16624,G1660,G14878);
  nand GNAME16625(G16625,G60086,G14876);
  nand GNAME16626(G16626,G60152,G14877);
  nand GNAME16627(G16627,G1690,G14878);
  nand GNAME16628(G16628,G60085,G14876);
  nand GNAME16629(G16629,G60153,G14877);
  nand GNAME16630(G16630,G1689,G14878);
  nand GNAME16631(G16631,G60084,G14876);
  nand GNAME16632(G16632,G60154,G14877);
  nand GNAME16633(G16633,G1688,G14878);
  nand GNAME16634(G16634,G60083,G14876);
  nand GNAME16635(G16635,G60155,G14877);
  nand GNAME16636(G16636,G1687,G14878);
  nand GNAME16637(G16637,G60082,G14876);
  nand GNAME16638(G16638,G60156,G14877);
  nand GNAME16639(G16639,G1686,G14878);
  nand GNAME16640(G16640,G60081,G14876);
  nand GNAME16641(G16641,G60157,G14877);
  nand GNAME16642(G16642,G60080,G14876);
  nand GNAME16643(G16643,G1685,G14878);
  nand GNAME16644(G16644,G60158,G14877);
  nand GNAME16645(G16645,G14784,G14813);
  nand GNAME16646(G16646,G60079,G14879);
  nand GNAME16647(G16647,G23488,G14880);
  nand GNAME16648(G16648,G23190,G14881);
  nand GNAME16649(G16649,G23901,G14882);
  nand GNAME16650(G16650,G60238,G14883);
  nand GNAME16651(G16651,G60078,G14879);
  nand GNAME16652(G16652,G23427,G14880);
  nand GNAME16653(G16653,G23122,G14881);
  nand GNAME16654(G16654,G23902,G14882);
  nand GNAME16655(G16655,G60237,G14883);
  nand GNAME16656(G16656,G60077,G14879);
  nand GNAME16657(G16657,G23475,G14880);
  nand GNAME16658(G16658,G23176,G14881);
  nand GNAME16659(G16659,G23940,G14882);
  nand GNAME16660(G16660,G60236,G14883);
  nand GNAME16661(G16661,G60076,G14879);
  nand GNAME16662(G16662,G23476,G14880);
  nand GNAME16663(G16663,G23177,G14881);
  nand GNAME16664(G16664,G23941,G14882);
  nand GNAME16665(G16665,G60235,G14883);
  nand GNAME16666(G16666,G60075,G14879);
  nand GNAME16667(G16667,G23477,G14880);
  nand GNAME16668(G16668,G23178,G14881);
  nand GNAME16669(G16669,G23942,G14882);
  nand GNAME16670(G16670,G60234,G14883);
  nand GNAME16671(G16671,G60074,G14879);
  nand GNAME16672(G16672,G23478,G14880);
  nand GNAME16673(G16673,G23179,G14881);
  nand GNAME16674(G16674,G23943,G14882);
  nand GNAME16675(G16675,G60233,G14883);
  nand GNAME16676(G16676,G60073,G14879);
  nand GNAME16677(G16677,G23479,G14880);
  nand GNAME16678(G16678,G23180,G14881);
  nand GNAME16679(G16679,G23944,G14882);
  nand GNAME16680(G16680,G60232,G14883);
  nand GNAME16681(G16681,G60072,G14879);
  nand GNAME16682(G16682,G23517,G14880);
  nand GNAME16683(G16683,G23181,G14881);
  nand GNAME16684(G16684,G23945,G14882);
  nand GNAME16685(G16685,G60231,G14883);
  nand GNAME16686(G16686,G60071,G14879);
  nand GNAME16687(G16687,G23520,G14880);
  nand GNAME16688(G16688,G23182,G14881);
  nand GNAME16689(G16689,G23946,G14882);
  nand GNAME16690(G16690,G60230,G14883);
  nand GNAME16691(G16691,G60070,G14879);
  nand GNAME16692(G16692,G23523,G14880);
  nand GNAME16693(G16693,G23183,G14881);
  nand GNAME16694(G16694,G23947,G14882);
  nand GNAME16695(G16695,G60229,G14883);
  nand GNAME16696(G16696,G60069,G14879);
  nand GNAME16697(G16697,G23526,G14880);
  nand GNAME16698(G16698,G23184,G14881);
  nand GNAME16699(G16699,G23948,G14882);
  nand GNAME16700(G16700,G60228,G14883);
  nand GNAME16701(G16701,G60068,G14879);
  nand GNAME16702(G16702,G23529,G14880);
  nand GNAME16703(G16703,G23185,G14881);
  nand GNAME16704(G16704,G23949,G14882);
  nand GNAME16705(G16705,G60227,G14883);
  nand GNAME16706(G16706,G60067,G14879);
  nand GNAME16707(G16707,G23535,G14880);
  nand GNAME16708(G16708,G23186,G14881);
  nand GNAME16709(G16709,G23953,G14882);
  nand GNAME16710(G16710,G60226,G14883);
  nand GNAME16711(G16711,G60066,G14879);
  nand GNAME16712(G16712,G23538,G14880);
  nand GNAME16713(G16713,G23187,G14881);
  nand GNAME16714(G16714,G23954,G14882);
  nand GNAME16715(G16715,G60225,G14883);
  nand GNAME16716(G16716,G60065,G14879);
  nand GNAME16717(G16717,G23541,G14880);
  nand GNAME16718(G16718,G23188,G14881);
  nand GNAME16719(G16719,G23955,G14882);
  nand GNAME16720(G16720,G60224,G14883);
  nand GNAME16721(G16721,G60064,G14879);
  nand GNAME16722(G16722,G23480,G14880);
  nand GNAME16723(G16723,G23216,G14881);
  nand GNAME16724(G16724,G23956,G14882);
  nand GNAME16725(G16725,G60223,G14883);
  nand GNAME16726(G16726,G60063,G14879);
  nand GNAME16727(G16727,G23481,G14880);
  nand GNAME16728(G16728,G23219,G14881);
  nand GNAME16729(G16729,G23957,G14882);
  nand GNAME16730(G16730,G60222,G14883);
  nand GNAME16731(G16731,G60062,G14879);
  nand GNAME16732(G16732,G23425,G14880);
  nand GNAME16733(G16733,G23191,G14881);
  nand GNAME16734(G16734,G23903,G14882);
  nand GNAME16735(G16735,G60221,G14883);
  nand GNAME16736(G16736,G60061,G14879);
  nand GNAME16737(G16737,G23482,G14880);
  nand GNAME16738(G16738,G23223,G14881);
  nand GNAME16739(G16739,G23958,G14882);
  nand GNAME16740(G16740,G60220,G14883);
  nand GNAME16741(G16741,G60060,G14879);
  nand GNAME16742(G16742,G23483,G14880);
  nand GNAME16743(G16743,G23226,G14881);
  nand GNAME16744(G16744,G23959,G14882);
  nand GNAME16745(G16745,G60219,G14883);
  nand GNAME16746(G16746,G60059,G14879);
  nand GNAME16747(G16747,G23484,G14880);
  nand GNAME16748(G16748,G23192,G14881);
  nand GNAME16749(G16749,G23839,G14882);
  nand GNAME16750(G16750,G60218,G14883);
  nand GNAME16751(G16751,G60058,G14879);
  nand GNAME16752(G16752,G23424,G14880);
  nand GNAME16753(G16753,G23120,G14881);
  nand GNAME16754(G16754,G23838,G14882);
  nand GNAME16755(G16755,G60217,G14883);
  nand GNAME16756(G16756,G60057,G14879);
  nand GNAME16757(G16757,G23461,G14880);
  nand GNAME16758(G16758,G23199,G14881);
  nand GNAME16759(G16759,G23930,G14882);
  nand GNAME16760(G16760,G60216,G14883);
  nand GNAME16761(G16761,G60056,G14879);
  nand GNAME16762(G16762,G23496,G14880);
  nand GNAME16763(G16763,G23156,G14881);
  nand GNAME16764(G16764,G23931,G14882);
  nand GNAME16765(G16765,G60215,G14883);
  nand GNAME16766(G16766,G60055,G14879);
  nand GNAME16767(G16767,G23486,G14880);
  nand GNAME16768(G16768,G23157,G14881);
  nand GNAME16769(G16769,G23899,G14882);
  nand GNAME16770(G16770,G60214,G14883);
  nand GNAME16771(G16771,G60054,G14879);
  nand GNAME16772(G16772,G23428,G14880);
  nand GNAME16773(G16773,G23123,G14881);
  nand GNAME16774(G16774,G23841,G14882);
  nand GNAME16775(G16775,G60213,G14883);
  nand GNAME16776(G16776,G60053,G14879);
  nand GNAME16777(G16777,G23500,G14880);
  nand GNAME16778(G16778,G23158,G14881);
  nand GNAME16779(G16779,G23935,G14882);
  nand GNAME16780(G16780,G60212,G14883);
  nand GNAME16781(G16781,G60052,G14879);
  nand GNAME16782(G16782,G23503,G14880);
  nand GNAME16783(G16783,G23159,G14881);
  nand GNAME16784(G16784,G23938,G14882);
  nand GNAME16785(G16785,G60211,G14883);
  nand GNAME16786(G16786,G60051,G14879);
  nand GNAME16787(G16787,G23900,G14882);
  nand GNAME16788(G16788,G60210,G14883);
  nand GNAME16789(G16789,G23160,G14881);
  nand GNAME16790(G16790,G23487,G14880);
  nand GNAME16791(G16791,G60050,G14879);
  nand GNAME16792(G16792,G23840,G14882);
  nand GNAME16793(G16793,G60209,G14883);
  nand GNAME16794(G16794,G23121,G14881);
  nand GNAME16795(G16795,G23426,G14880);
  nand GNAME16796(G16796,G60049,G14879);
  nand GNAME16797(G16797,G23952,G14882);
  nand GNAME16798(G16798,G23532,G14880);
  nand GNAME16799(G16799,G23213,G14881);
  nand GNAME16800(G16800,G60208,G14883);
  nand GNAME16801(G16801,G60048,G14879);
  nand GNAME16802(G16802,G23898,G14882);
  nand GNAME16803(G16803,G23189,G14881);
  nand GNAME16804(G16804,G60207,G14883);
  nand GNAME16805(G16805,G23485,G14880);
  nand GNAME16806(G16806,G14777,G14781);
  nand GNAME16807(G16807,G15846,G14823);
  nand GNAME16808(G16808,G14780,G15846);
  nand GNAME16809(G16809,G16808,G14884);
  nand GNAME16810(G16810,G14780,G14779);
  nand GNAME16811(G16811,G15780,G15829);
  nand GNAME16812(G16812,G15897,G14746,G14793);
  nand GNAME16813(G16813,G16812,G15914);
  nand GNAME16814(G16814,G15829,G15974);
  nand GNAME16815(G16815,G16814,G15880);
  nand GNAME16816(G16816,G16815,G15846);
  nand GNAME16817(G16817,G14778,G15974);
  nand GNAME16818(G16818,G16816,G16817);
  nand GNAME16819(G16819,G14746,G16818);
  nand GNAME16820(G16820,G16819,G15897);
  nand GNAME16821(G16821,G23753,G16813,G15880);
  nand GNAME16822(G16822,G16820,G23088);
  nand GNAME16823(G16823,G14885,G16821,G16822);
  nand GNAME16824(G16824,G16823,G14797);
  nand GNAME16825(G16825,G14784,G14807);
  or GNAME16826(G16826,G14825,G14819,G14783,G16316);
  nand GNAME16827(G16827,G14888,G14780,G14794);
  or GNAME16828(G16828,G15897,G14747);
  nand GNAME16829(G16829,G16318,G16827,G16828,G14899);
  nand GNAME16830(G16830,G15246,G15931);
  nand GNAME16831(G16831,G14778,G14743);
  nand GNAME16832(G16832,G15897,G15778,G15948);
  nand GNAME16833(G16833,G16832,G15931);
  nand GNAME16834(G16834,G14778,G14820);
  nand GNAME16835(G16835,G15802,G14857);
  or GNAME16836(G16836,G14747,G14780);
  nand GNAME16837(G16837,G19967,G14850);
  nand GNAME16838(G16838,G16837,G15786);
  nand GNAME16839(G16839,G14789,G14893);
  nand GNAME16840(G16840,G15931,G14894);
  nand GNAME16841(G16841,G14896,G14897);
  nand GNAME16842(G16842,G8108,G14887);
  nand GNAME16843(G16843,G23488,G14898);
  nand GNAME16844(G16844,G23190,G14900);
  nand GNAME16845(G16845,G23901,G14901);
  nand GNAME16846(G16846,G60238,G14902);
  nand GNAME16847(G16847,G14903,G60047);
  nand GNAME16848(G16848,G14903,G60046);
  nand GNAME16849(G16849,G14887,G8107);
  nand GNAME16850(G16850,G23427,G14898);
  nand GNAME16851(G16851,G23122,G14900);
  nand GNAME16852(G16852,G23902,G14901);
  nand GNAME16853(G16853,G60237,G14902);
  nand GNAME16854(G16854,G14903,G60045);
  nand GNAME16855(G16855,G14887,G14029);
  nand GNAME16856(G16856,G23475,G14898);
  nand GNAME16857(G16857,G23176,G14900);
  nand GNAME16858(G16858,G23940,G14901);
  nand GNAME16859(G16859,G60236,G14902);
  nand GNAME16860(G16860,G14903,G60044);
  nand GNAME16861(G16861,G14887,G14030);
  nand GNAME16862(G16862,G23476,G14898);
  nand GNAME16863(G16863,G23177,G14900);
  nand GNAME16864(G16864,G23941,G14901);
  nand GNAME16865(G16865,G60235,G14902);
  nand GNAME16866(G16866,G14903,G60043);
  nand GNAME16867(G16867,G14887,G8105);
  nand GNAME16868(G16868,G23477,G14898);
  nand GNAME16869(G16869,G23178,G14900);
  nand GNAME16870(G16870,G23942,G14901);
  nand GNAME16871(G16871,G60234,G14902);
  nand GNAME16872(G16872,G14903,G60042);
  nand GNAME16873(G16873,G14887,G14031);
  nand GNAME16874(G16874,G23478,G14898);
  nand GNAME16875(G16875,G23179,G14900);
  nand GNAME16876(G16876,G23943,G14901);
  nand GNAME16877(G16877,G60233,G14902);
  nand GNAME16878(G16878,G14903,G60041);
  nand GNAME16879(G16879,G14887,G14032);
  nand GNAME16880(G16880,G23479,G14898);
  nand GNAME16881(G16881,G23180,G14900);
  nand GNAME16882(G16882,G23944,G14901);
  nand GNAME16883(G16883,G60232,G14902);
  nand GNAME16884(G16884,G14903,G60040);
  nand GNAME16885(G16885,G14887,G8081);
  nand GNAME16886(G16886,G23517,G14898);
  nand GNAME16887(G16887,G23181,G14900);
  nand GNAME16888(G16888,G23945,G14901);
  nand GNAME16889(G16889,G60231,G14902);
  nand GNAME16890(G16890,G14903,G60039);
  nand GNAME16891(G16891,G14887,G8080);
  nand GNAME16892(G16892,G23520,G14898);
  nand GNAME16893(G16893,G23182,G14900);
  nand GNAME16894(G16894,G23946,G14901);
  nand GNAME16895(G16895,G60230,G14902);
  nand GNAME16896(G16896,G14887,G8079);
  nand GNAME16897(G16897,G23523,G14898);
  nand GNAME16898(G16898,G23183,G14900);
  nand GNAME16899(G16899,G23947,G14901);
  nand GNAME16900(G16900,G60229,G14902);
  nand GNAME16901(G16901,G14903,G60038);
  nand GNAME16902(G16902,G14887,G8078);
  nand GNAME16903(G16903,G23526,G14898);
  nand GNAME16904(G16904,G23184,G14900);
  nand GNAME16905(G16905,G23948,G14901);
  nand GNAME16906(G16906,G60228,G14902);
  nand GNAME16907(G16907,G14903,G60037);
  nand GNAME16908(G16908,G14887,G8077);
  nand GNAME16909(G16909,G23529,G14898);
  nand GNAME16910(G16910,G23185,G14900);
  nand GNAME16911(G16911,G23949,G14901);
  nand GNAME16912(G16912,G60227,G14902);
  nand GNAME16913(G16913,G14903,G60036);
  nand GNAME16914(G16914,G14887,G8075);
  nand GNAME16915(G16915,G23535,G14898);
  nand GNAME16916(G16916,G23186,G14900);
  nand GNAME16917(G16917,G23953,G14901);
  nand GNAME16918(G16918,G60226,G14902);
  nand GNAME16919(G16919,G14903,G60035);
  nand GNAME16920(G16920,G14887,G8074);
  nand GNAME16921(G16921,G23538,G14898);
  nand GNAME16922(G16922,G23187,G14900);
  nand GNAME16923(G16923,G23954,G14901);
  nand GNAME16924(G16924,G60225,G14902);
  nand GNAME16925(G16925,G14903,G60034);
  nand GNAME16926(G16926,G14887,G8073);
  nand GNAME16927(G16927,G23541,G14898);
  nand GNAME16928(G16928,G23188,G14900);
  nand GNAME16929(G16929,G23955,G14901);
  nand GNAME16930(G16930,G60224,G14902);
  nand GNAME16931(G16931,G14903,G60033);
  nand GNAME16932(G16932,G14887,G8103);
  nand GNAME16933(G16933,G23480,G14898);
  nand GNAME16934(G16934,G23216,G14900);
  nand GNAME16935(G16935,G23956,G14901);
  nand GNAME16936(G16936,G60223,G14902);
  nand GNAME16937(G16937,G14903,G60032);
  nand GNAME16938(G16938,G14887,G8102);
  nand GNAME16939(G16939,G23481,G14898);
  nand GNAME16940(G16940,G23219,G14900);
  nand GNAME16941(G16941,G23957,G14901);
  nand GNAME16942(G16942,G60222,G14902);
  nand GNAME16943(G16943,G14903,G60031);
  nand GNAME16944(G16944,G14887,G8101);
  nand GNAME16945(G16945,G23425,G14898);
  nand GNAME16946(G16946,G23191,G14900);
  nand GNAME16947(G16947,G23903,G14901);
  nand GNAME16948(G16948,G60221,G14902);
  nand GNAME16949(G16949,G14903,G60030);
  nand GNAME16950(G16950,G14887,G8100);
  nand GNAME16951(G16951,G23482,G14898);
  nand GNAME16952(G16952,G23223,G14900);
  nand GNAME16953(G16953,G23958,G14901);
  nand GNAME16954(G16954,G60220,G14902);
  nand GNAME16955(G16955,G14903,G60029);
  nand GNAME16956(G16956,G14887,G8099);
  nand GNAME16957(G16957,G23483,G14898);
  nand GNAME16958(G16958,G23226,G14900);
  nand GNAME16959(G16959,G23959,G14901);
  nand GNAME16960(G16960,G60219,G14902);
  nand GNAME16961(G16961,G14903,G60028);
  nand GNAME16962(G16962,G14887,G8098);
  nand GNAME16963(G16963,G23484,G14898);
  nand GNAME16964(G16964,G23192,G14900);
  nand GNAME16965(G16965,G23839,G14901);
  nand GNAME16966(G16966,G60218,G14902);
  nand GNAME16967(G16967,G14903,G60027);
  nand GNAME16968(G16968,G14887,G8097);
  nand GNAME16969(G16969,G23424,G14898);
  nand GNAME16970(G16970,G23120,G14900);
  nand GNAME16971(G16971,G23838,G14901);
  nand GNAME16972(G16972,G60217,G14902);
  nand GNAME16973(G16973,G14903,G60026);
  nand GNAME16974(G16974,G14887,G13988);
  nand GNAME16975(G16975,G23461,G14898);
  nand GNAME16976(G16976,G23199,G14900);
  nand GNAME16977(G16977,G23930,G14901);
  nand GNAME16978(G16978,G60216,G14902);
  nand GNAME16979(G16979,G14903,G60025);
  nand GNAME16980(G16980,G14887,G8114);
  nand GNAME16981(G16981,G23496,G14898);
  nand GNAME16982(G16982,G23156,G14900);
  nand GNAME16983(G16983,G23931,G14901);
  nand GNAME16984(G16984,G60215,G14902);
  nand GNAME16985(G16985,G14903,G60024);
  nand GNAME16986(G16986,G14887,G8113);
  nand GNAME16987(G16987,G23486,G14898);
  nand GNAME16988(G16988,G23157,G14900);
  nand GNAME16989(G16989,G23899,G14901);
  nand GNAME16990(G16990,G60214,G14902);
  nand GNAME16991(G16991,G14903,G60023);
  nand GNAME16992(G16992,G14887,G8112);
  nand GNAME16993(G16993,G23428,G14898);
  nand GNAME16994(G16994,G23123,G14900);
  nand GNAME16995(G16995,G23841,G14901);
  nand GNAME16996(G16996,G60213,G14902);
  nand GNAME16997(G16997,G14903,G60022);
  nand GNAME16998(G16998,G14887,G8111);
  nand GNAME16999(G16999,G23500,G14898);
  nand GNAME17000(G17000,G23158,G14900);
  nand GNAME17001(G17001,G23935,G14901);
  nand GNAME17002(G17002,G60212,G14902);
  nand GNAME17003(G17003,G14903,G60021);
  nand GNAME17004(G17004,G14887,G8110);
  nand GNAME17005(G17005,G23503,G14898);
  nand GNAME17006(G17006,G23159,G14900);
  nand GNAME17007(G17007,G23938,G14901);
  nand GNAME17008(G17008,G60211,G14902);
  nand GNAME17009(G17009,G14903,G60020);
  nand GNAME17010(G17010,G14887,G8109);
  nand GNAME17011(G17011,G23900,G14901);
  nand GNAME17012(G17012,G60210,G14902);
  nand GNAME17013(G17013,G23160,G14900);
  nand GNAME17014(G17014,G23487,G14898);
  nand GNAME17015(G17015,G14903,G60019);
  nand GNAME17016(G17016,G14887,G8106);
  nand GNAME17017(G17017,G23840,G14901);
  nand GNAME17018(G17018,G60209,G14902);
  nand GNAME17019(G17019,G23121,G14900);
  nand GNAME17020(G17020,G23426,G14898);
  nand GNAME17021(G17021,G14903,G60018);
  nand GNAME17022(G17022,G14887,G8104);
  nand GNAME17023(G17023,G23952,G14901);
  nand GNAME17024(G17024,G23532,G14898);
  nand GNAME17025(G17025,G60208,G14902);
  nand GNAME17026(G17026,G23213,G14900);
  nand GNAME17027(G17027,G14903,G60017);
  nand GNAME17028(G17028,G14887,G8096);
  nand GNAME17029(G17029,G23898,G14901);
  nand GNAME17030(G17030,G60207,G14902);
  nand GNAME17031(G17031,G23485,G14898);
  nand GNAME17032(G17032,G23189,G14900);
  nand GNAME17033(G17033,G14903,G60016);
  or GNAME17034(G17034,G14798,G14906);
  not GNAME17035(G17035,G14907);
  or GNAME17036(G17036,G23088,G19981);
  not GNAME17037(G17037,G14914);
  nand GNAME17038(G17038,G60010,G14792);
  nor GNAME17039(G17039,G14782,G59876);
  nand GNAME17040(G17040,G14909,G14910);
  not GNAME17041(G17041,G14911);
  nand GNAME17042(G17042,G14748,G15793);
  nand GNAME17043(G17043,G17042,G15796);
  nand GNAME17044(G17044,G17041,G14912);
  nand GNAME17045(G17045,G23189,G14913);
  nand GNAME17046(G17046,G14904,G19864,G19865);
  nand GNAME17047(G17047,G14742,G14792);
  not GNAME17048(G17048,G14917);
  nand GNAME17049(G17049,G14748,G14949);
  nand GNAME17050(G17050,G60009,G14792);
  nand GNAME17051(G17051,G14810,G60014);
  not GNAME17052(G17052,G14918);
  nand GNAME17053(G17053,G15247,G14912);
  nand GNAME17054(G17054,G23213,G14913);
  nand GNAME17055(G17055,G17037,G60014);
  nand GNAME17056(G17056,G14748,G15248);
  nand GNAME17057(G17057,G60008,G14792);
  nand GNAME17058(G17058,G14810,G60013);
  nand GNAME17059(G17059,G14918,G15798);
  nand GNAME17060(G17060,G17059,G17048);
  nand GNAME17061(G17061,G14916,G17052);
  nand GNAME17062(G17062,G14922,G14921);
  not GNAME17063(G17063,G14923);
  nand GNAME17064(G17064,G14912,G17063);
  nand GNAME17065(G17065,G23121,G14913);
  nand GNAME17066(G17066,G17037,G60013);
  nor GNAME17067(G17067,G14920,G14925);
  nand GNAME17068(G17068,G14748,G14950);
  nand GNAME17069(G17069,G60007,G14792);
  nand GNAME17070(G17070,G14810,G60012);
  nand GNAME17071(G17071,G14912,G19876);
  nand GNAME17072(G17072,G23160,G14913);
  nand GNAME17073(G17073,G17037,G60012);
  nand GNAME17074(G17074,G16467,G14796);
  nand GNAME17075(G17075,G17074,G15974);
  nand GNAME17076(G17076,G17075,G16318);
  nand GNAME17077(G17077,G17076,G23088);
  nand GNAME17078(G17078,G14783,G23753);
  nand GNAME17079(G17079,G17077,G17078);
  nand GNAME17080(G17080,G14746,G17079);
  or GNAME17081(G17081,G15102,G14798);
  nand GNAME17082(G17082,G15775,G14797);
  nand GNAME17083(G17083,G15973,G14891);
  nand GNAME17084(G17084,G17083,G19452);
  nand GNAME17085(G17085,G14789,G59875);
  nand GNAME17086(G17086,G17085,G15772,G15799);
  not GNAME17087(G17087,G14927);
  nand GNAME17088(G17088,G14789,G17087);
  nand GNAME17089(G17089,G17088,G59875);
  nand GNAME17090(G17090,G14911,G14927);
  not GNAME17091(G17091,G14930);
  nand GNAME17092(G17092,G15863,G14927,G59875);
  not GNAME17093(G17093,G14928);
  nand GNAME17094(G17094,G14794,G14888);
  nand GNAME17095(G17095,G17094,G14747);
  nand GNAME17096(G17096,G14780,G17095);
  nand GNAME17097(G17097,G15863,G14893);
  nand GNAME17098(G17098,G14858,G16318,G17096,G17097);
  nand GNAME17099(G17099,G14793,G14818);
  nand GNAME17100(G17100,G17099,G14897);
  nand GNAME17101(G17101,G15949,G14895);
  nand GNAME17102(G17102,G14852,G16467);
  or GNAME17103(G17103,G60010,G15102);
  nand GNAME17104(G17104,G17102,G17093);
  nand GNAME17105(G17105,G17101,G17041);
  nand GNAME17106(G17106,G17100,G23189);
  nand GNAME17107(G17107,G17098,G23485);
  nand GNAME17108(G17108,G17106,G17107,G17105,G17103,G17104);
  nand GNAME17109(G17109,G14911,G19861);
  nand GNAME17110(G17110,G23485,G14926);
  nand GNAME17111(G17111,G17109,G59876);
  nand GNAME17112(G17112,G17108,G14787);
  nand GNAME17113(G17113,G17112,G17110,G17111);
  nand GNAME17114(G17114,G17086,G60009);
  nand GNAME17115(G17115,G14748,G15247);
  not GNAME17116(G17116,G14931);
  not GNAME17117(G17117,G15184);
  nand GNAME17118(G17118,G60010,G15863);
  not GNAME17119(G17119,G15158);
  or GNAME17120(G17120,G14751,G17119);
  nand GNAME17121(G17121,G17120,G14822);
  nand GNAME17122(G17122,G17102,G19883);
  nand GNAME17123(G17123,G17101,G15247);
  nand GNAME17124(G17124,G17100,G23213);
  nand GNAME17125(G17125,G17098,G23532);
  nand GNAME17126(G17126,G15184,G14825);
  nand GNAME17127(G17127,G15398,G17123,G17125,G17122);
  nand GNAME17128(G17128,G15247,G14929);
  nand GNAME17129(G17129,G23532,G14926);
  nand GNAME17130(G17130,G17127,G14787);
  nand GNAME17131(G17131,G17130,G17128,G17129);
  nand GNAME17132(G17132,G14931,G17091);
  nand GNAME17133(G17133,G15772,G17132);
  nand GNAME17134(G17134,G14930,G17116);
  not GNAME17135(G17135,G14933);
  nand GNAME17136(G17136,G17086,G60008);
  nand GNAME17137(G17137,G14748,G17063);
  not GNAME17138(G17138,G14932);
  nand GNAME17139(G17139,G15784,G15252);
  not GNAME17140(G17140,G14934);
  not GNAME17141(G17141,G15773);
  nand GNAME17142(G17142,G17102,G19889);
  nand GNAME17143(G17143,G17101,G17063);
  nand GNAME17144(G17144,G17100,G23121);
  nand GNAME17145(G17145,G17098,G23426);
  nand GNAME17146(G17146,G14822,G19895);
  nand GNAME17147(G17147,G14825,G17140);
  nand GNAME17148(G17148,G15399,G17144,G17142,G17145);
  nand GNAME17149(G17149,G17063,G14929);
  nand GNAME17150(G17150,G23426,G14926);
  nand GNAME17151(G17151,G17148,G14787);
  nand GNAME17152(G17152,G17151,G17149,G17150);
  nand GNAME17153(G17153,G17086,G60007);
  nand GNAME17154(G17154,G17153,G17159);
  nand GNAME17155(G17155,G17160,G17135);
  nand GNAME17156(G17156,G17157,G17154,G17155);
  nand GNAME17157(G17157,G14932,G14817);
  nand GNAME17158(G17158,G14933,G17157);
  nand GNAME17159(G17159,G14748,G19876);
  nand GNAME17160(G17160,G15799,G17138);
  nand GNAME17161(G17161,G17153,G17158,G17159,G17160);
  not GNAME17162(G17162,G14938);
  nand GNAME17163(G17163,G17141,G14750);
  nand GNAME17164(G17164,G14758,G17141);
  nand GNAME17165(G17165,G17164,G60007);
  and GNAME17166(G17166,G14765,G15863);
  or GNAME17167(G17167,G17166,G14750);
  nand GNAME17168(G17168,G14789,G14771);
  not GNAME17169(G17169,G14935);
  nand GNAME17170(G17170,G17102,G14938);
  nand GNAME17171(G17171,G17101,G19876);
  nand GNAME17172(G17172,G17100,G23160);
  nand GNAME17173(G17173,G17098,G23487);
  nand GNAME17174(G17174,G14825,G17169);
  nand GNAME17175(G17175,G14822,G15803);
  nand GNAME17176(G17176,G15400,G17172,G17170,G17173);
  nand GNAME17177(G17177,G23487,G14926);
  nand GNAME17178(G17178,G17176,G14787);
  nand GNAME17179(G17179,G17177,G17178);
  nand GNAME17180(G17180,G14789,G14959);
  nand GNAME17181(G17181,G59875,G14956);
  nand GNAME17182(G17182,G17180,G17181);
  not GNAME17183(G17183,G14944);
  nand GNAME17184(G17184,G14830,G14953);
  nand GNAME17185(G17185,G59875,G17183);
  nand GNAME17186(G17186,G17184,G17185);
  nand GNAME17187(G17187,G14944,G14945);
  and GNAME17188(G17188,G17187,G15797);
  nand GNAME17189(G17189,G14953,G14944,G14945);
  nand GNAME17190(G17190,G14954,G14955);
  nand GNAME17191(G17191,G17189,G17190);
  and GNAME17192(G17192,G14944,G59875);
  nor GNAME17193(G17193,G17192,G14799,G14955);
  or GNAME17194(G17194,G14954,G17193);
  nand GNAME17195(G17195,G17194,G14907);
  nand GNAME17196(G17196,G1684,G14946);
  nand GNAME17197(G17197,G17195,G60005);
  nand GNAME17198(G17198,G17191,G1691);
  nand GNAME17199(G17199,G17186,G14956);
  nand GNAME17200(G17200,G14957,G14958);
  nand GNAME17201(G17201,G17182,G14954);
  nand GNAME17202(G17202,G14793,G14959);
  nand GNAME17203(G17203,G59875,G14960);
  nand GNAME17204(G17204,G17202,G17203);
  nand GNAME17205(G17205,G1683,G14946);
  nand GNAME17206(G17206,G17195,G60004);
  nand GNAME17207(G17207,G17191,G1680);
  nand GNAME17208(G17208,G17186,G14960);
  nand GNAME17209(G17209,G14957,G14961);
  nand GNAME17210(G17210,G17204,G14954);
  nand GNAME17211(G17211,G14778,G14959);
  nand GNAME17212(G17212,G59875,G14962);
  nand GNAME17213(G17213,G17211,G17212);
  nand GNAME17214(G17214,G1682,G14946);
  nand GNAME17215(G17215,G17195,G60003);
  nand GNAME17216(G17216,G17191,G1669);
  nand GNAME17217(G17217,G17186,G14962);
  nand GNAME17218(G17218,G14957,G14963);
  nand GNAME17219(G17219,G17213,G14954);
  nand GNAME17220(G17220,G14743,G14959);
  nand GNAME17221(G17221,G59875,G14964);
  nand GNAME17222(G17222,G17220,G17221);
  nand GNAME17223(G17223,G1681,G14946);
  nand GNAME17224(G17224,G17195,G60002);
  nand GNAME17225(G17225,G17191,G1666);
  nand GNAME17226(G17226,G17186,G14964);
  nand GNAME17227(G17227,G14957,G14965);
  nand GNAME17228(G17228,G17222,G14954);
  nand GNAME17229(G17229,G14780,G14959);
  nand GNAME17230(G17230,G59875,G14966);
  nand GNAME17231(G17231,G17229,G17230);
  nand GNAME17232(G17232,G1679,G14946);
  nand GNAME17233(G17233,G17195,G60001);
  nand GNAME17234(G17234,G17191,G1665);
  nand GNAME17235(G17235,G17186,G14966);
  nand GNAME17236(G17236,G14957,G14967);
  nand GNAME17237(G17237,G17231,G14954);
  nand GNAME17238(G17238,G14777,G14959);
  nand GNAME17239(G17239,G59875,G14968);
  nand GNAME17240(G17240,G17238,G17239);
  nand GNAME17241(G17241,G1678,G14946);
  nand GNAME17242(G17242,G17195,G60000);
  nand GNAME17243(G17243,G17191,G1664);
  nand GNAME17244(G17244,G17186,G14968);
  nand GNAME17245(G17245,G14957,G14969);
  nand GNAME17246(G17246,G17240,G14954);
  nand GNAME17247(G17247,G14779,G14959);
  nand GNAME17248(G17248,G59875,G14970);
  nand GNAME17249(G17249,G17247,G17248);
  nand GNAME17250(G17250,G1677,G14946);
  nand GNAME17251(G17251,G17195,G59999);
  nand GNAME17252(G17252,G17191,G1663);
  nand GNAME17253(G17253,G17186,G14970);
  nand GNAME17254(G17254,G14957,G14971);
  nand GNAME17255(G17255,G17249,G14954);
  nand GNAME17256(G17256,G14849,G14959);
  nand GNAME17257(G17257,G59875,G14972);
  nand GNAME17258(G17258,G17256,G17257);
  nand GNAME17259(G17259,G1676,G14946);
  nand GNAME17260(G17260,G17195,G59998);
  nand GNAME17261(G17261,G17191,G1662);
  nand GNAME17262(G17262,G17186,G14972);
  nand GNAME17263(G17263,G14957,G14973);
  nand GNAME17264(G17264,G17258,G14954);
  not GNAME17265(G17265,G14976);
  nand GNAME17266(G17266,G14830,G14981);
  nand GNAME17267(G17267,G59875,G17265);
  nand GNAME17268(G17268,G17266,G17267);
  nand GNAME17269(G17269,G14976,G14977);
  and GNAME17270(G17270,G17269,G15797);
  nand GNAME17271(G17271,G14981,G14976,G14977);
  nand GNAME17272(G17272,G14982,G14983);
  nand GNAME17273(G17273,G17271,G17272);
  and GNAME17274(G17274,G14976,G59875);
  nor GNAME17275(G17275,G17274,G14799,G14983);
  or GNAME17276(G17276,G14982,G17275);
  nand GNAME17277(G17277,G17276,G14907);
  nand GNAME17278(G17278,G1684,G14978);
  nand GNAME17279(G17279,G17277,G59997);
  nand GNAME17280(G17280,G17273,G1691);
  nand GNAME17281(G17281,G17268,G14956);
  nand GNAME17282(G17282,G14958,G14984);
  nand GNAME17283(G17283,G17182,G14982);
  nand GNAME17284(G17284,G1683,G14978);
  nand GNAME17285(G17285,G17277,G59996);
  nand GNAME17286(G17286,G17273,G1680);
  nand GNAME17287(G17287,G17268,G14960);
  nand GNAME17288(G17288,G14961,G14984);
  nand GNAME17289(G17289,G17204,G14982);
  nand GNAME17290(G17290,G1682,G14978);
  nand GNAME17291(G17291,G17277,G59995);
  nand GNAME17292(G17292,G17273,G1669);
  nand GNAME17293(G17293,G17268,G14962);
  nand GNAME17294(G17294,G14963,G14984);
  nand GNAME17295(G17295,G17213,G14982);
  nand GNAME17296(G17296,G1681,G14978);
  nand GNAME17297(G17297,G17277,G59994);
  nand GNAME17298(G17298,G17273,G1666);
  nand GNAME17299(G17299,G17268,G14964);
  nand GNAME17300(G17300,G14965,G14984);
  nand GNAME17301(G17301,G17222,G14982);
  nand GNAME17302(G17302,G1679,G14978);
  nand GNAME17303(G17303,G17277,G59993);
  nand GNAME17304(G17304,G17273,G1665);
  nand GNAME17305(G17305,G17268,G14966);
  nand GNAME17306(G17306,G14967,G14984);
  nand GNAME17307(G17307,G17231,G14982);
  nand GNAME17308(G17308,G1678,G14978);
  nand GNAME17309(G17309,G17277,G59992);
  nand GNAME17310(G17310,G17273,G1664);
  nand GNAME17311(G17311,G17268,G14968);
  nand GNAME17312(G17312,G14969,G14984);
  nand GNAME17313(G17313,G17240,G14982);
  nand GNAME17314(G17314,G1677,G14978);
  nand GNAME17315(G17315,G17277,G59991);
  nand GNAME17316(G17316,G17273,G1663);
  nand GNAME17317(G17317,G17268,G14970);
  nand GNAME17318(G17318,G14971,G14984);
  nand GNAME17319(G17319,G17249,G14982);
  nand GNAME17320(G17320,G1676,G14978);
  nand GNAME17321(G17321,G17277,G59990);
  nand GNAME17322(G17322,G17273,G1662);
  nand GNAME17323(G17323,G17268,G14972);
  nand GNAME17324(G17324,G14973,G14984);
  nand GNAME17325(G17325,G17258,G14982);
  not GNAME17326(G17326,G14987);
  nand GNAME17327(G17327,G14830,G14992);
  nand GNAME17328(G17328,G59875,G17326);
  nand GNAME17329(G17329,G17327,G17328);
  nand GNAME17330(G17330,G14987,G14988);
  and GNAME17331(G17331,G17330,G15797);
  nand GNAME17332(G17332,G14992,G14987,G14988);
  nand GNAME17333(G17333,G14993,G14994);
  nand GNAME17334(G17334,G17332,G17333);
  and GNAME17335(G17335,G14987,G59875);
  nor GNAME17336(G17336,G17335,G14799,G14994);
  or GNAME17337(G17337,G14993,G17336);
  nand GNAME17338(G17338,G17337,G14907);
  nand GNAME17339(G17339,G1684,G14989);
  nand GNAME17340(G17340,G17338,G59989);
  nand GNAME17341(G17341,G17334,G1691);
  nand GNAME17342(G17342,G17329,G14956);
  nand GNAME17343(G17343,G14958,G14995);
  nand GNAME17344(G17344,G17182,G14993);
  nand GNAME17345(G17345,G1683,G14989);
  nand GNAME17346(G17346,G17338,G59988);
  nand GNAME17347(G17347,G17334,G1680);
  nand GNAME17348(G17348,G17329,G14960);
  nand GNAME17349(G17349,G14961,G14995);
  nand GNAME17350(G17350,G17204,G14993);
  nand GNAME17351(G17351,G1682,G14989);
  nand GNAME17352(G17352,G17338,G59987);
  nand GNAME17353(G17353,G17334,G1669);
  nand GNAME17354(G17354,G17329,G14962);
  nand GNAME17355(G17355,G14963,G14995);
  nand GNAME17356(G17356,G17213,G14993);
  nand GNAME17357(G17357,G1681,G14989);
  nand GNAME17358(G17358,G17338,G59986);
  nand GNAME17359(G17359,G17334,G1666);
  nand GNAME17360(G17360,G17329,G14964);
  nand GNAME17361(G17361,G14965,G14995);
  nand GNAME17362(G17362,G17222,G14993);
  nand GNAME17363(G17363,G1679,G14989);
  nand GNAME17364(G17364,G17338,G59985);
  nand GNAME17365(G17365,G17334,G1665);
  nand GNAME17366(G17366,G17329,G14966);
  nand GNAME17367(G17367,G14967,G14995);
  nand GNAME17368(G17368,G17231,G14993);
  nand GNAME17369(G17369,G1678,G14989);
  nand GNAME17370(G17370,G17338,G59984);
  nand GNAME17371(G17371,G17334,G1664);
  nand GNAME17372(G17372,G17329,G14968);
  nand GNAME17373(G17373,G14969,G14995);
  nand GNAME17374(G17374,G17240,G14993);
  nand GNAME17375(G17375,G1677,G14989);
  nand GNAME17376(G17376,G17338,G59983);
  nand GNAME17377(G17377,G17334,G1663);
  nand GNAME17378(G17378,G17329,G14970);
  nand GNAME17379(G17379,G14971,G14995);
  nand GNAME17380(G17380,G17249,G14993);
  nand GNAME17381(G17381,G1676,G14989);
  nand GNAME17382(G17382,G17338,G59982);
  nand GNAME17383(G17383,G17334,G1662);
  nand GNAME17384(G17384,G17329,G14972);
  nand GNAME17385(G17385,G14973,G14995);
  nand GNAME17386(G17386,G17258,G14993);
  not GNAME17387(G17387,G14996);
  nand GNAME17388(G17388,G14830,G15000);
  nand GNAME17389(G17389,G59875,G17387);
  nand GNAME17390(G17390,G17388,G17389);
  nand GNAME17391(G17391,G14996,G14997);
  and GNAME17392(G17392,G17391,G15797);
  nand GNAME17393(G17393,G14997,G15000);
  nand GNAME17394(G17394,G15001,G15002);
  nand GNAME17395(G17395,G17393,G17394);
  and GNAME17396(G17396,G14996,G59875);
  nor GNAME17397(G17397,G17396,G14799,G15002);
  or GNAME17398(G17398,G15001,G17397);
  nand GNAME17399(G17399,G17398,G14907);
  nand GNAME17400(G17400,G1684,G14998);
  nand GNAME17401(G17401,G17399,G59981);
  nand GNAME17402(G17402,G17395,G1691);
  nand GNAME17403(G17403,G17390,G14956);
  nand GNAME17404(G17404,G14958,G15003);
  nand GNAME17405(G17405,G17182,G15001);
  nand GNAME17406(G17406,G1683,G14998);
  nand GNAME17407(G17407,G17399,G59980);
  nand GNAME17408(G17408,G17395,G1680);
  nand GNAME17409(G17409,G17390,G14960);
  nand GNAME17410(G17410,G14961,G15003);
  nand GNAME17411(G17411,G17204,G15001);
  nand GNAME17412(G17412,G1682,G14998);
  nand GNAME17413(G17413,G17399,G59979);
  nand GNAME17414(G17414,G17395,G1669);
  nand GNAME17415(G17415,G17390,G14962);
  nand GNAME17416(G17416,G14963,G15003);
  nand GNAME17417(G17417,G17213,G15001);
  nand GNAME17418(G17418,G1681,G14998);
  nand GNAME17419(G17419,G17399,G59978);
  nand GNAME17420(G17420,G17395,G1666);
  nand GNAME17421(G17421,G17390,G14964);
  nand GNAME17422(G17422,G14965,G15003);
  nand GNAME17423(G17423,G17222,G15001);
  nand GNAME17424(G17424,G1679,G14998);
  nand GNAME17425(G17425,G17399,G59977);
  nand GNAME17426(G17426,G17395,G1665);
  nand GNAME17427(G17427,G17390,G14966);
  nand GNAME17428(G17428,G14967,G15003);
  nand GNAME17429(G17429,G17231,G15001);
  nand GNAME17430(G17430,G1678,G14998);
  nand GNAME17431(G17431,G17399,G59976);
  nand GNAME17432(G17432,G17395,G1664);
  nand GNAME17433(G17433,G17390,G14968);
  nand GNAME17434(G17434,G14969,G15003);
  nand GNAME17435(G17435,G17240,G15001);
  nand GNAME17436(G17436,G1677,G14998);
  nand GNAME17437(G17437,G17399,G59975);
  nand GNAME17438(G17438,G17395,G1663);
  nand GNAME17439(G17439,G17390,G14970);
  nand GNAME17440(G17440,G14971,G15003);
  nand GNAME17441(G17441,G17249,G15001);
  nand GNAME17442(G17442,G1676,G14998);
  nand GNAME17443(G17443,G17399,G59974);
  nand GNAME17444(G17444,G17395,G1662);
  nand GNAME17445(G17445,G17390,G14972);
  nand GNAME17446(G17446,G14973,G15003);
  nand GNAME17447(G17447,G17258,G15001);
  not GNAME17448(G17448,G15006);
  nand GNAME17449(G17449,G14830,G15010);
  nand GNAME17450(G17450,G59875,G17448);
  nand GNAME17451(G17451,G17449,G17450);
  nand GNAME17452(G17452,G15006,G15007);
  and GNAME17453(G17453,G17452,G15797);
  nand GNAME17454(G17454,G15010,G15006,G15007);
  nand GNAME17455(G17455,G15011,G15012);
  nand GNAME17456(G17456,G17454,G17455);
  and GNAME17457(G17457,G15006,G59875);
  nor GNAME17458(G17458,G17457,G14799,G15012);
  or GNAME17459(G17459,G15011,G17458);
  nand GNAME17460(G17460,G17459,G14907);
  nand GNAME17461(G17461,G1684,G15008);
  nand GNAME17462(G17462,G17460,G59973);
  nand GNAME17463(G17463,G17456,G1691);
  nand GNAME17464(G17464,G17451,G14956);
  nand GNAME17465(G17465,G14958,G15013);
  nand GNAME17466(G17466,G17182,G15011);
  nand GNAME17467(G17467,G1683,G15008);
  nand GNAME17468(G17468,G17460,G59972);
  nand GNAME17469(G17469,G17456,G1680);
  nand GNAME17470(G17470,G17451,G14960);
  nand GNAME17471(G17471,G14961,G15013);
  nand GNAME17472(G17472,G17204,G15011);
  nand GNAME17473(G17473,G1682,G15008);
  nand GNAME17474(G17474,G17460,G59971);
  nand GNAME17475(G17475,G17456,G1669);
  nand GNAME17476(G17476,G17451,G14962);
  nand GNAME17477(G17477,G14963,G15013);
  nand GNAME17478(G17478,G17213,G15011);
  nand GNAME17479(G17479,G1681,G15008);
  nand GNAME17480(G17480,G17460,G59970);
  nand GNAME17481(G17481,G17456,G1666);
  nand GNAME17482(G17482,G17451,G14964);
  nand GNAME17483(G17483,G14965,G15013);
  nand GNAME17484(G17484,G17222,G15011);
  nand GNAME17485(G17485,G1679,G15008);
  nand GNAME17486(G17486,G17460,G59969);
  nand GNAME17487(G17487,G17456,G1665);
  nand GNAME17488(G17488,G17451,G14966);
  nand GNAME17489(G17489,G14967,G15013);
  nand GNAME17490(G17490,G17231,G15011);
  nand GNAME17491(G17491,G1678,G15008);
  nand GNAME17492(G17492,G17460,G59968);
  nand GNAME17493(G17493,G17456,G1664);
  nand GNAME17494(G17494,G17451,G14968);
  nand GNAME17495(G17495,G14969,G15013);
  nand GNAME17496(G17496,G17240,G15011);
  nand GNAME17497(G17497,G1677,G15008);
  nand GNAME17498(G17498,G17460,G59967);
  nand GNAME17499(G17499,G17456,G1663);
  nand GNAME17500(G17500,G17451,G14970);
  nand GNAME17501(G17501,G14971,G15013);
  nand GNAME17502(G17502,G17249,G15011);
  nand GNAME17503(G17503,G1676,G15008);
  nand GNAME17504(G17504,G17460,G59966);
  nand GNAME17505(G17505,G17456,G1662);
  nand GNAME17506(G17506,G17451,G14972);
  nand GNAME17507(G17507,G14973,G15013);
  nand GNAME17508(G17508,G17258,G15011);
  not GNAME17509(G17509,G15016);
  nand GNAME17510(G17510,G14830,G15019);
  nand GNAME17511(G17511,G59875,G17509);
  nand GNAME17512(G17512,G17510,G17511);
  nand GNAME17513(G17513,G15016,G15017);
  and GNAME17514(G17514,G17513,G15797);
  nand GNAME17515(G17515,G15017,G15019);
  nand GNAME17516(G17516,G15020,G15021);
  nand GNAME17517(G17517,G17515,G17516);
  and GNAME17518(G17518,G15016,G59875);
  nor GNAME17519(G17519,G17518,G14799,G15021);
  or GNAME17520(G17520,G15020,G17519);
  nand GNAME17521(G17521,G17520,G14907);
  nand GNAME17522(G17522,G1684,G15018);
  nand GNAME17523(G17523,G17521,G59965);
  nand GNAME17524(G17524,G17517,G1691);
  nand GNAME17525(G17525,G17512,G14956);
  nand GNAME17526(G17526,G14958,G15022);
  nand GNAME17527(G17527,G17182,G15020);
  nand GNAME17528(G17528,G1683,G15018);
  nand GNAME17529(G17529,G17521,G59964);
  nand GNAME17530(G17530,G17517,G1680);
  nand GNAME17531(G17531,G17512,G14960);
  nand GNAME17532(G17532,G14961,G15022);
  nand GNAME17533(G17533,G17204,G15020);
  nand GNAME17534(G17534,G1682,G15018);
  nand GNAME17535(G17535,G17521,G59963);
  nand GNAME17536(G17536,G17517,G1669);
  nand GNAME17537(G17537,G17512,G14962);
  nand GNAME17538(G17538,G14963,G15022);
  nand GNAME17539(G17539,G17213,G15020);
  nand GNAME17540(G17540,G1681,G15018);
  nand GNAME17541(G17541,G17521,G59962);
  nand GNAME17542(G17542,G17517,G1666);
  nand GNAME17543(G17543,G17512,G14964);
  nand GNAME17544(G17544,G14965,G15022);
  nand GNAME17545(G17545,G17222,G15020);
  nand GNAME17546(G17546,G1679,G15018);
  nand GNAME17547(G17547,G17521,G59961);
  nand GNAME17548(G17548,G17517,G1665);
  nand GNAME17549(G17549,G17512,G14966);
  nand GNAME17550(G17550,G14967,G15022);
  nand GNAME17551(G17551,G17231,G15020);
  nand GNAME17552(G17552,G1678,G15018);
  nand GNAME17553(G17553,G17521,G59960);
  nand GNAME17554(G17554,G17517,G1664);
  nand GNAME17555(G17555,G17512,G14968);
  nand GNAME17556(G17556,G14969,G15022);
  nand GNAME17557(G17557,G17240,G15020);
  nand GNAME17558(G17558,G1677,G15018);
  nand GNAME17559(G17559,G17521,G59959);
  nand GNAME17560(G17560,G17517,G1663);
  nand GNAME17561(G17561,G17512,G14970);
  nand GNAME17562(G17562,G14971,G15022);
  nand GNAME17563(G17563,G17249,G15020);
  nand GNAME17564(G17564,G1676,G15018);
  nand GNAME17565(G17565,G17521,G59958);
  nand GNAME17566(G17566,G17517,G1662);
  nand GNAME17567(G17567,G17512,G14972);
  nand GNAME17568(G17568,G14973,G15022);
  nand GNAME17569(G17569,G17258,G15020);
  not GNAME17570(G17570,G15023);
  nand GNAME17571(G17571,G14830,G15026);
  nand GNAME17572(G17572,G59875,G17570);
  nand GNAME17573(G17573,G17571,G17572);
  nand GNAME17574(G17574,G15023,G15024);
  and GNAME17575(G17575,G17574,G15797);
  nand GNAME17576(G17576,G15026,G15023,G15024);
  nand GNAME17577(G17577,G15027,G15028);
  nand GNAME17578(G17578,G17576,G17577);
  and GNAME17579(G17579,G15023,G59875);
  nor GNAME17580(G17580,G17579,G14799,G15028);
  or GNAME17581(G17581,G15027,G17580);
  nand GNAME17582(G17582,G17581,G14907);
  nand GNAME17583(G17583,G1684,G15025);
  nand GNAME17584(G17584,G17582,G59957);
  nand GNAME17585(G17585,G17578,G1691);
  nand GNAME17586(G17586,G17573,G14956);
  nand GNAME17587(G17587,G14958,G15029);
  nand GNAME17588(G17588,G17182,G15027);
  nand GNAME17589(G17589,G1683,G15025);
  nand GNAME17590(G17590,G17582,G59956);
  nand GNAME17591(G17591,G17578,G1680);
  nand GNAME17592(G17592,G17573,G14960);
  nand GNAME17593(G17593,G14961,G15029);
  nand GNAME17594(G17594,G17204,G15027);
  nand GNAME17595(G17595,G1682,G15025);
  nand GNAME17596(G17596,G17582,G59955);
  nand GNAME17597(G17597,G17578,G1669);
  nand GNAME17598(G17598,G17573,G14962);
  nand GNAME17599(G17599,G14963,G15029);
  nand GNAME17600(G17600,G17213,G15027);
  nand GNAME17601(G17601,G1681,G15025);
  nand GNAME17602(G17602,G17582,G59954);
  nand GNAME17603(G17603,G17578,G1666);
  nand GNAME17604(G17604,G17573,G14964);
  nand GNAME17605(G17605,G14965,G15029);
  nand GNAME17606(G17606,G17222,G15027);
  nand GNAME17607(G17607,G1679,G15025);
  nand GNAME17608(G17608,G17582,G59953);
  nand GNAME17609(G17609,G17578,G1665);
  nand GNAME17610(G17610,G17573,G14966);
  nand GNAME17611(G17611,G14967,G15029);
  nand GNAME17612(G17612,G17231,G15027);
  nand GNAME17613(G17613,G1678,G15025);
  nand GNAME17614(G17614,G17582,G59952);
  nand GNAME17615(G17615,G17578,G1664);
  nand GNAME17616(G17616,G17573,G14968);
  nand GNAME17617(G17617,G14969,G15029);
  nand GNAME17618(G17618,G17240,G15027);
  nand GNAME17619(G17619,G1677,G15025);
  nand GNAME17620(G17620,G17582,G59951);
  nand GNAME17621(G17621,G17578,G1663);
  nand GNAME17622(G17622,G17573,G14970);
  nand GNAME17623(G17623,G14971,G15029);
  nand GNAME17624(G17624,G17249,G15027);
  nand GNAME17625(G17625,G1676,G15025);
  nand GNAME17626(G17626,G17582,G59950);
  nand GNAME17627(G17627,G17578,G1662);
  nand GNAME17628(G17628,G17573,G14972);
  nand GNAME17629(G17629,G14973,G15029);
  nand GNAME17630(G17630,G17258,G15027);
  not GNAME17631(G17631,G15030);
  nand GNAME17632(G17632,G14830,G15033);
  nand GNAME17633(G17633,G59875,G17631);
  nand GNAME17634(G17634,G17632,G17633);
  nand GNAME17635(G17635,G15030,G15031);
  and GNAME17636(G17636,G17635,G15797);
  nand GNAME17637(G17637,G15031,G15033);
  nand GNAME17638(G17638,G15034,G15035);
  nand GNAME17639(G17639,G17637,G17638);
  and GNAME17640(G17640,G15030,G59875);
  nor GNAME17641(G17641,G17640,G14799,G15034);
  or GNAME17642(G17642,G15035,G17641);
  nand GNAME17643(G17643,G17642,G14907);
  nand GNAME17644(G17644,G1684,G15032);
  nand GNAME17645(G17645,G17643,G59949);
  nand GNAME17646(G17646,G17639,G1691);
  nand GNAME17647(G17647,G17634,G14956);
  nand GNAME17648(G17648,G14958,G15036);
  nand GNAME17649(G17649,G17182,G15035);
  nand GNAME17650(G17650,G1683,G15032);
  nand GNAME17651(G17651,G17643,G59948);
  nand GNAME17652(G17652,G17639,G1680);
  nand GNAME17653(G17653,G17634,G14960);
  nand GNAME17654(G17654,G14961,G15036);
  nand GNAME17655(G17655,G17204,G15035);
  nand GNAME17656(G17656,G1682,G15032);
  nand GNAME17657(G17657,G17643,G59947);
  nand GNAME17658(G17658,G17639,G1669);
  nand GNAME17659(G17659,G17634,G14962);
  nand GNAME17660(G17660,G14963,G15036);
  nand GNAME17661(G17661,G17213,G15035);
  nand GNAME17662(G17662,G1681,G15032);
  nand GNAME17663(G17663,G17643,G59946);
  nand GNAME17664(G17664,G17639,G1666);
  nand GNAME17665(G17665,G17634,G14964);
  nand GNAME17666(G17666,G14965,G15036);
  nand GNAME17667(G17667,G17222,G15035);
  nand GNAME17668(G17668,G1679,G15032);
  nand GNAME17669(G17669,G17643,G59945);
  nand GNAME17670(G17670,G17639,G1665);
  nand GNAME17671(G17671,G17634,G14966);
  nand GNAME17672(G17672,G14967,G15036);
  nand GNAME17673(G17673,G17231,G15035);
  nand GNAME17674(G17674,G1678,G15032);
  nand GNAME17675(G17675,G17643,G59944);
  nand GNAME17676(G17676,G17639,G1664);
  nand GNAME17677(G17677,G17634,G14968);
  nand GNAME17678(G17678,G14969,G15036);
  nand GNAME17679(G17679,G17240,G15035);
  nand GNAME17680(G17680,G1677,G15032);
  nand GNAME17681(G17681,G17643,G59943);
  nand GNAME17682(G17682,G17639,G1663);
  nand GNAME17683(G17683,G17634,G14970);
  nand GNAME17684(G17684,G14971,G15036);
  nand GNAME17685(G17685,G17249,G15035);
  nand GNAME17686(G17686,G1676,G15032);
  nand GNAME17687(G17687,G17643,G59942);
  nand GNAME17688(G17688,G17639,G1662);
  nand GNAME17689(G17689,G17634,G14972);
  nand GNAME17690(G17690,G14973,G15036);
  nand GNAME17691(G17691,G17258,G15035);
  not GNAME17692(G17692,G15039);
  nand GNAME17693(G17693,G59875,G17692);
  nand GNAME17694(G17694,G14830,G15044);
  nand GNAME17695(G17695,G17693,G17694);
  nand GNAME17696(G17696,G15039,G15040);
  and GNAME17697(G17697,G17696,G15797);
  nand GNAME17698(G17698,G15044,G15039,G15040);
  nand GNAME17699(G17699,G15045,G15046);
  nand GNAME17700(G17700,G17698,G17699);
  and GNAME17701(G17701,G15039,G59875);
  nor GNAME17702(G17702,G17701,G14799,G15046);
  or GNAME17703(G17703,G15045,G17702);
  nand GNAME17704(G17704,G17703,G14907);
  nand GNAME17705(G17705,G1684,G15041);
  nand GNAME17706(G17706,G17704,G59941);
  nand GNAME17707(G17707,G17700,G1691);
  nand GNAME17708(G17708,G17695,G14956);
  nand GNAME17709(G17709,G14958,G15047);
  nand GNAME17710(G17710,G17182,G15045);
  nand GNAME17711(G17711,G1683,G15041);
  nand GNAME17712(G17712,G17704,G59940);
  nand GNAME17713(G17713,G17700,G1680);
  nand GNAME17714(G17714,G17695,G14960);
  nand GNAME17715(G17715,G14961,G15047);
  nand GNAME17716(G17716,G17204,G15045);
  nand GNAME17717(G17717,G1682,G15041);
  nand GNAME17718(G17718,G17704,G59939);
  nand GNAME17719(G17719,G17700,G1669);
  nand GNAME17720(G17720,G17695,G14962);
  nand GNAME17721(G17721,G14963,G15047);
  nand GNAME17722(G17722,G17213,G15045);
  nand GNAME17723(G17723,G1681,G15041);
  nand GNAME17724(G17724,G17704,G59938);
  nand GNAME17725(G17725,G17700,G1666);
  nand GNAME17726(G17726,G17695,G14964);
  nand GNAME17727(G17727,G14965,G15047);
  nand GNAME17728(G17728,G17222,G15045);
  nand GNAME17729(G17729,G1679,G15041);
  nand GNAME17730(G17730,G17704,G59937);
  nand GNAME17731(G17731,G17700,G1665);
  nand GNAME17732(G17732,G17695,G14966);
  nand GNAME17733(G17733,G14967,G15047);
  nand GNAME17734(G17734,G17231,G15045);
  nand GNAME17735(G17735,G1678,G15041);
  nand GNAME17736(G17736,G17704,G59936);
  nand GNAME17737(G17737,G17700,G1664);
  nand GNAME17738(G17738,G17695,G14968);
  nand GNAME17739(G17739,G14969,G15047);
  nand GNAME17740(G17740,G17240,G15045);
  nand GNAME17741(G17741,G1677,G15041);
  nand GNAME17742(G17742,G17704,G59935);
  nand GNAME17743(G17743,G17700,G1663);
  nand GNAME17744(G17744,G17695,G14970);
  nand GNAME17745(G17745,G14971,G15047);
  nand GNAME17746(G17746,G17249,G15045);
  nand GNAME17747(G17747,G1676,G15041);
  nand GNAME17748(G17748,G17704,G59934);
  nand GNAME17749(G17749,G17700,G1662);
  nand GNAME17750(G17750,G17695,G14972);
  nand GNAME17751(G17751,G14973,G15047);
  nand GNAME17752(G17752,G17258,G15045);
  not GNAME17753(G17753,G15048);
  nand GNAME17754(G17754,G59875,G17753);
  nand GNAME17755(G17755,G14830,G15051);
  nand GNAME17756(G17756,G17754,G17755);
  nand GNAME17757(G17757,G15048,G15049);
  and GNAME17758(G17758,G17757,G15797);
  nand GNAME17759(G17759,G15051,G15048,G15049);
  nand GNAME17760(G17760,G15052,G15053);
  nand GNAME17761(G17761,G17759,G17760);
  and GNAME17762(G17762,G15048,G59875);
  nor GNAME17763(G17763,G17762,G14799,G15053);
  or GNAME17764(G17764,G15052,G17763);
  nand GNAME17765(G17765,G17764,G14907);
  nand GNAME17766(G17766,G1684,G15050);
  nand GNAME17767(G17767,G17765,G59933);
  nand GNAME17768(G17768,G17761,G1691);
  nand GNAME17769(G17769,G17756,G14956);
  nand GNAME17770(G17770,G14958,G15054);
  nand GNAME17771(G17771,G17182,G15052);
  nand GNAME17772(G17772,G1683,G15050);
  nand GNAME17773(G17773,G17765,G59932);
  nand GNAME17774(G17774,G17761,G1680);
  nand GNAME17775(G17775,G17756,G14960);
  nand GNAME17776(G17776,G14961,G15054);
  nand GNAME17777(G17777,G17204,G15052);
  nand GNAME17778(G17778,G1682,G15050);
  nand GNAME17779(G17779,G17765,G59931);
  nand GNAME17780(G17780,G17761,G1669);
  nand GNAME17781(G17781,G17756,G14962);
  nand GNAME17782(G17782,G14963,G15054);
  nand GNAME17783(G17783,G17213,G15052);
  nand GNAME17784(G17784,G1681,G15050);
  nand GNAME17785(G17785,G17765,G59930);
  nand GNAME17786(G17786,G17761,G1666);
  nand GNAME17787(G17787,G17756,G14964);
  nand GNAME17788(G17788,G14965,G15054);
  nand GNAME17789(G17789,G17222,G15052);
  nand GNAME17790(G17790,G1679,G15050);
  nand GNAME17791(G17791,G17765,G59929);
  nand GNAME17792(G17792,G17761,G1665);
  nand GNAME17793(G17793,G17756,G14966);
  nand GNAME17794(G17794,G14967,G15054);
  nand GNAME17795(G17795,G17231,G15052);
  nand GNAME17796(G17796,G1678,G15050);
  nand GNAME17797(G17797,G17765,G59928);
  nand GNAME17798(G17798,G17761,G1664);
  nand GNAME17799(G17799,G17756,G14968);
  nand GNAME17800(G17800,G14969,G15054);
  nand GNAME17801(G17801,G17240,G15052);
  nand GNAME17802(G17802,G1677,G15050);
  nand GNAME17803(G17803,G17765,G59927);
  nand GNAME17804(G17804,G17761,G1663);
  nand GNAME17805(G17805,G17756,G14970);
  nand GNAME17806(G17806,G14971,G15054);
  nand GNAME17807(G17807,G17249,G15052);
  nand GNAME17808(G17808,G1676,G15050);
  nand GNAME17809(G17809,G17765,G59926);
  nand GNAME17810(G17810,G17761,G1662);
  nand GNAME17811(G17811,G17756,G14972);
  nand GNAME17812(G17812,G14973,G15054);
  nand GNAME17813(G17813,G17258,G15052);
  not GNAME17814(G17814,G15057);
  nand GNAME17815(G17815,G59875,G17814);
  nand GNAME17816(G17816,G14830,G15060);
  nand GNAME17817(G17817,G17815,G17816);
  nand GNAME17818(G17818,G15057,G15058);
  and GNAME17819(G17819,G17818,G15797);
  nand GNAME17820(G17820,G15060,G15057,G15058);
  nand GNAME17821(G17821,G15061,G15062);
  nand GNAME17822(G17822,G17820,G17821);
  and GNAME17823(G17823,G15057,G59875);
  nor GNAME17824(G17824,G17823,G14799,G15062);
  or GNAME17825(G17825,G15061,G17824);
  nand GNAME17826(G17826,G17825,G14907);
  nand GNAME17827(G17827,G1684,G15059);
  nand GNAME17828(G17828,G17826,G59925);
  nand GNAME17829(G17829,G17822,G1691);
  nand GNAME17830(G17830,G17817,G14956);
  nand GNAME17831(G17831,G14958,G15063);
  nand GNAME17832(G17832,G17182,G15061);
  nand GNAME17833(G17833,G1683,G15059);
  nand GNAME17834(G17834,G17826,G59924);
  nand GNAME17835(G17835,G17822,G1680);
  nand GNAME17836(G17836,G17817,G14960);
  nand GNAME17837(G17837,G14961,G15063);
  nand GNAME17838(G17838,G17204,G15061);
  nand GNAME17839(G17839,G1682,G15059);
  nand GNAME17840(G17840,G17826,G59923);
  nand GNAME17841(G17841,G17822,G1669);
  nand GNAME17842(G17842,G17817,G14962);
  nand GNAME17843(G17843,G14963,G15063);
  nand GNAME17844(G17844,G17213,G15061);
  nand GNAME17845(G17845,G1681,G15059);
  nand GNAME17846(G17846,G17826,G59922);
  nand GNAME17847(G17847,G17822,G1666);
  nand GNAME17848(G17848,G17817,G14964);
  nand GNAME17849(G17849,G14965,G15063);
  nand GNAME17850(G17850,G17222,G15061);
  nand GNAME17851(G17851,G1679,G15059);
  nand GNAME17852(G17852,G17826,G59921);
  nand GNAME17853(G17853,G17822,G1665);
  nand GNAME17854(G17854,G17817,G14966);
  nand GNAME17855(G17855,G14967,G15063);
  nand GNAME17856(G17856,G17231,G15061);
  nand GNAME17857(G17857,G1678,G15059);
  nand GNAME17858(G17858,G17826,G59920);
  nand GNAME17859(G17859,G17822,G1664);
  nand GNAME17860(G17860,G17817,G14968);
  nand GNAME17861(G17861,G14969,G15063);
  nand GNAME17862(G17862,G17240,G15061);
  nand GNAME17863(G17863,G1677,G15059);
  nand GNAME17864(G17864,G17826,G59919);
  nand GNAME17865(G17865,G17822,G1663);
  nand GNAME17866(G17866,G17817,G14970);
  nand GNAME17867(G17867,G14971,G15063);
  nand GNAME17868(G17868,G17249,G15061);
  nand GNAME17869(G17869,G1676,G15059);
  nand GNAME17870(G17870,G17826,G59918);
  nand GNAME17871(G17871,G17822,G1662);
  nand GNAME17872(G17872,G17817,G14972);
  nand GNAME17873(G17873,G14973,G15063);
  nand GNAME17874(G17874,G17258,G15061);
  not GNAME17875(G17875,G15064);
  nand GNAME17876(G17876,G59875,G17875);
  nand GNAME17877(G17877,G14830,G15067);
  nand GNAME17878(G17878,G17876,G17877);
  nand GNAME17879(G17879,G15064,G15065);
  and GNAME17880(G17880,G17879,G15797);
  nand GNAME17881(G17881,G15065,G15067);
  nand GNAME17882(G17882,G15068,G15069);
  nand GNAME17883(G17883,G17881,G17882);
  and GNAME17884(G17884,G15064,G59875);
  nor GNAME17885(G17885,G17884,G14799,G15069);
  or GNAME17886(G17886,G15068,G17885);
  nand GNAME17887(G17887,G17886,G14907);
  nand GNAME17888(G17888,G1684,G15066);
  nand GNAME17889(G17889,G17887,G59917);
  nand GNAME17890(G17890,G17883,G1691);
  nand GNAME17891(G17891,G17878,G14956);
  nand GNAME17892(G17892,G14958,G15070);
  nand GNAME17893(G17893,G17182,G15068);
  nand GNAME17894(G17894,G1683,G15066);
  nand GNAME17895(G17895,G17887,G59916);
  nand GNAME17896(G17896,G17883,G1680);
  nand GNAME17897(G17897,G17878,G14960);
  nand GNAME17898(G17898,G14961,G15070);
  nand GNAME17899(G17899,G17204,G15068);
  nand GNAME17900(G17900,G1682,G15066);
  nand GNAME17901(G17901,G17887,G59915);
  nand GNAME17902(G17902,G17883,G1669);
  nand GNAME17903(G17903,G17878,G14962);
  nand GNAME17904(G17904,G14963,G15070);
  nand GNAME17905(G17905,G17213,G15068);
  nand GNAME17906(G17906,G1681,G15066);
  nand GNAME17907(G17907,G17887,G59914);
  nand GNAME17908(G17908,G17883,G1666);
  nand GNAME17909(G17909,G17878,G14964);
  nand GNAME17910(G17910,G14965,G15070);
  nand GNAME17911(G17911,G17222,G15068);
  nand GNAME17912(G17912,G1679,G15066);
  nand GNAME17913(G17913,G17887,G59913);
  nand GNAME17914(G17914,G17883,G1665);
  nand GNAME17915(G17915,G17878,G14966);
  nand GNAME17916(G17916,G14967,G15070);
  nand GNAME17917(G17917,G17231,G15068);
  nand GNAME17918(G17918,G1678,G15066);
  nand GNAME17919(G17919,G17887,G59912);
  nand GNAME17920(G17920,G17883,G1664);
  nand GNAME17921(G17921,G17878,G14968);
  nand GNAME17922(G17922,G14969,G15070);
  nand GNAME17923(G17923,G17240,G15068);
  nand GNAME17924(G17924,G1677,G15066);
  nand GNAME17925(G17925,G17887,G59911);
  nand GNAME17926(G17926,G17883,G1663);
  nand GNAME17927(G17927,G17878,G14970);
  nand GNAME17928(G17928,G14971,G15070);
  nand GNAME17929(G17929,G17249,G15068);
  nand GNAME17930(G17930,G1676,G15066);
  nand GNAME17931(G17931,G17887,G59910);
  nand GNAME17932(G17932,G17883,G1662);
  nand GNAME17933(G17933,G17878,G14972);
  nand GNAME17934(G17934,G14973,G15070);
  nand GNAME17935(G17935,G17258,G15068);
  not GNAME17936(G17936,G15071);
  nand GNAME17937(G17937,G59875,G17936);
  nand GNAME17938(G17938,G14830,G15076);
  nand GNAME17939(G17939,G17937,G17938);
  nand GNAME17940(G17940,G15071,G15072);
  and GNAME17941(G17941,G17940,G15797);
  nand GNAME17942(G17942,G15076,G15071,G15072);
  nand GNAME17943(G17943,G15077,G15078);
  nand GNAME17944(G17944,G17942,G17943);
  and GNAME17945(G17945,G15071,G59875);
  nor GNAME17946(G17946,G17945,G14799,G15078);
  or GNAME17947(G17947,G15077,G17946);
  nand GNAME17948(G17948,G17947,G14907);
  nand GNAME17949(G17949,G1684,G15073);
  nand GNAME17950(G17950,G17948,G59909);
  nand GNAME17951(G17951,G17944,G1691);
  nand GNAME17952(G17952,G17939,G14956);
  nand GNAME17953(G17953,G14958,G15079);
  nand GNAME17954(G17954,G17182,G15077);
  nand GNAME17955(G17955,G1683,G15073);
  nand GNAME17956(G17956,G17948,G59908);
  nand GNAME17957(G17957,G17944,G1680);
  nand GNAME17958(G17958,G17939,G14960);
  nand GNAME17959(G17959,G14961,G15079);
  nand GNAME17960(G17960,G17204,G15077);
  nand GNAME17961(G17961,G1682,G15073);
  nand GNAME17962(G17962,G17948,G59907);
  nand GNAME17963(G17963,G17944,G1669);
  nand GNAME17964(G17964,G17939,G14962);
  nand GNAME17965(G17965,G14963,G15079);
  nand GNAME17966(G17966,G17213,G15077);
  nand GNAME17967(G17967,G1681,G15073);
  nand GNAME17968(G17968,G17948,G59906);
  nand GNAME17969(G17969,G17944,G1666);
  nand GNAME17970(G17970,G17939,G14964);
  nand GNAME17971(G17971,G14965,G15079);
  nand GNAME17972(G17972,G17222,G15077);
  nand GNAME17973(G17973,G1679,G15073);
  nand GNAME17974(G17974,G17948,G59905);
  nand GNAME17975(G17975,G17944,G1665);
  nand GNAME17976(G17976,G17939,G14966);
  nand GNAME17977(G17977,G14967,G15079);
  nand GNAME17978(G17978,G17231,G15077);
  nand GNAME17979(G17979,G1678,G15073);
  nand GNAME17980(G17980,G17948,G59904);
  nand GNAME17981(G17981,G17944,G1664);
  nand GNAME17982(G17982,G17939,G14968);
  nand GNAME17983(G17983,G14969,G15079);
  nand GNAME17984(G17984,G17240,G15077);
  nand GNAME17985(G17985,G1677,G15073);
  nand GNAME17986(G17986,G17948,G59903);
  nand GNAME17987(G17987,G17944,G1663);
  nand GNAME17988(G17988,G17939,G14970);
  nand GNAME17989(G17989,G14971,G15079);
  nand GNAME17990(G17990,G17249,G15077);
  nand GNAME17991(G17991,G1676,G15073);
  nand GNAME17992(G17992,G17948,G59902);
  nand GNAME17993(G17993,G17944,G1662);
  nand GNAME17994(G17994,G17939,G14972);
  nand GNAME17995(G17995,G14973,G15079);
  nand GNAME17996(G17996,G17258,G15077);
  not GNAME17997(G17997,G15080);
  nand GNAME17998(G17998,G59875,G17997);
  nand GNAME17999(G17999,G14830,G15083);
  nand GNAME18000(G18000,G17998,G17999);
  nand GNAME18001(G18001,G15080,G15081);
  and GNAME18002(G18002,G18001,G15797);
  nand GNAME18003(G18003,G15083,G15080,G15081);
  nand GNAME18004(G18004,G15084,G15085);
  nand GNAME18005(G18005,G18003,G18004);
  and GNAME18006(G18006,G15080,G59875);
  nor GNAME18007(G18007,G18006,G14799,G15085);
  or GNAME18008(G18008,G15084,G18007);
  nand GNAME18009(G18009,G18008,G14907);
  nand GNAME18010(G18010,G1684,G15082);
  nand GNAME18011(G18011,G18009,G59901);
  nand GNAME18012(G18012,G18005,G1691);
  nand GNAME18013(G18013,G18000,G14956);
  nand GNAME18014(G18014,G14958,G15086);
  nand GNAME18015(G18015,G17182,G15084);
  nand GNAME18016(G18016,G1683,G15082);
  nand GNAME18017(G18017,G18009,G59900);
  nand GNAME18018(G18018,G18005,G1680);
  nand GNAME18019(G18019,G18000,G14960);
  nand GNAME18020(G18020,G14961,G15086);
  nand GNAME18021(G18021,G17204,G15084);
  nand GNAME18022(G18022,G1682,G15082);
  nand GNAME18023(G18023,G18009,G59899);
  nand GNAME18024(G18024,G18005,G1669);
  nand GNAME18025(G18025,G18000,G14962);
  nand GNAME18026(G18026,G14963,G15086);
  nand GNAME18027(G18027,G17213,G15084);
  nand GNAME18028(G18028,G1681,G15082);
  nand GNAME18029(G18029,G18009,G59898);
  nand GNAME18030(G18030,G18005,G1666);
  nand GNAME18031(G18031,G18000,G14964);
  nand GNAME18032(G18032,G14965,G15086);
  nand GNAME18033(G18033,G17222,G15084);
  nand GNAME18034(G18034,G1679,G15082);
  nand GNAME18035(G18035,G18009,G59897);
  nand GNAME18036(G18036,G18005,G1665);
  nand GNAME18037(G18037,G18000,G14966);
  nand GNAME18038(G18038,G14967,G15086);
  nand GNAME18039(G18039,G17231,G15084);
  nand GNAME18040(G18040,G1678,G15082);
  nand GNAME18041(G18041,G18009,G59896);
  nand GNAME18042(G18042,G18005,G1664);
  nand GNAME18043(G18043,G18000,G14968);
  nand GNAME18044(G18044,G14969,G15086);
  nand GNAME18045(G18045,G17240,G15084);
  nand GNAME18046(G18046,G1677,G15082);
  nand GNAME18047(G18047,G18009,G59895);
  nand GNAME18048(G18048,G18005,G1663);
  nand GNAME18049(G18049,G18000,G14970);
  nand GNAME18050(G18050,G14971,G15086);
  nand GNAME18051(G18051,G17249,G15084);
  nand GNAME18052(G18052,G1676,G15082);
  nand GNAME18053(G18053,G18009,G59894);
  nand GNAME18054(G18054,G18005,G1662);
  nand GNAME18055(G18055,G18000,G14972);
  nand GNAME18056(G18056,G14973,G15086);
  nand GNAME18057(G18057,G17258,G15084);
  not GNAME18058(G18058,G15087);
  nand GNAME18059(G18059,G59875,G18058);
  nand GNAME18060(G18060,G14830,G15090);
  nand GNAME18061(G18061,G18059,G18060);
  nand GNAME18062(G18062,G15087,G15088);
  and GNAME18063(G18063,G18062,G15797);
  nand GNAME18064(G18064,G15090,G15087,G15088);
  nand GNAME18065(G18065,G15091,G15092);
  nand GNAME18066(G18066,G18064,G18065);
  and GNAME18067(G18067,G15087,G59875);
  nor GNAME18068(G18068,G18067,G14799,G15092);
  or GNAME18069(G18069,G15091,G18068);
  nand GNAME18070(G18070,G18069,G14907);
  nand GNAME18071(G18071,G1684,G15089);
  nand GNAME18072(G18072,G18070,G59893);
  nand GNAME18073(G18073,G18066,G1691);
  nand GNAME18074(G18074,G18061,G14956);
  nand GNAME18075(G18075,G14958,G15093);
  nand GNAME18076(G18076,G17182,G15091);
  nand GNAME18077(G18077,G1683,G15089);
  nand GNAME18078(G18078,G18070,G59892);
  nand GNAME18079(G18079,G18066,G1680);
  nand GNAME18080(G18080,G18061,G14960);
  nand GNAME18081(G18081,G14961,G15093);
  nand GNAME18082(G18082,G17204,G15091);
  nand GNAME18083(G18083,G1682,G15089);
  nand GNAME18084(G18084,G18070,G59891);
  nand GNAME18085(G18085,G18066,G1669);
  nand GNAME18086(G18086,G18061,G14962);
  nand GNAME18087(G18087,G14963,G15093);
  nand GNAME18088(G18088,G17213,G15091);
  nand GNAME18089(G18089,G1681,G15089);
  nand GNAME18090(G18090,G18070,G59890);
  nand GNAME18091(G18091,G18066,G1666);
  nand GNAME18092(G18092,G18061,G14964);
  nand GNAME18093(G18093,G14965,G15093);
  nand GNAME18094(G18094,G17222,G15091);
  nand GNAME18095(G18095,G1679,G15089);
  nand GNAME18096(G18096,G18070,G59889);
  nand GNAME18097(G18097,G18066,G1665);
  nand GNAME18098(G18098,G18061,G14966);
  nand GNAME18099(G18099,G14967,G15093);
  nand GNAME18100(G18100,G17231,G15091);
  nand GNAME18101(G18101,G1678,G15089);
  nand GNAME18102(G18102,G18070,G59888);
  nand GNAME18103(G18103,G18066,G1664);
  nand GNAME18104(G18104,G18061,G14968);
  nand GNAME18105(G18105,G14969,G15093);
  nand GNAME18106(G18106,G17240,G15091);
  nand GNAME18107(G18107,G1677,G15089);
  nand GNAME18108(G18108,G18070,G59887);
  nand GNAME18109(G18109,G18066,G1663);
  nand GNAME18110(G18110,G18061,G14970);
  nand GNAME18111(G18111,G14971,G15093);
  nand GNAME18112(G18112,G17249,G15091);
  nand GNAME18113(G18113,G1676,G15089);
  nand GNAME18114(G18114,G18070,G59886);
  nand GNAME18115(G18115,G18066,G1662);
  nand GNAME18116(G18116,G18061,G14972);
  nand GNAME18117(G18117,G14973,G15093);
  nand GNAME18118(G18118,G17258,G15091);
  not GNAME18119(G18119,G15094);
  nand GNAME18120(G18120,G59875,G18119);
  nand GNAME18121(G18121,G14830,G15097);
  nand GNAME18122(G18122,G18120,G18121);
  nand GNAME18123(G18123,G15094,G15095);
  and GNAME18124(G18124,G18123,G15797);
  nand GNAME18125(G18125,G15095,G15097);
  nand GNAME18126(G18126,G15098,G15099);
  nand GNAME18127(G18127,G18125,G18126);
  and GNAME18128(G18128,G15094,G59875);
  nor GNAME18129(G18129,G18128,G14799,G15098);
  or GNAME18130(G18130,G15099,G18129);
  nand GNAME18131(G18131,G18130,G14907);
  nand GNAME18132(G18132,G1684,G15096);
  nand GNAME18133(G18133,G18131,G59885);
  nand GNAME18134(G18134,G18127,G1691);
  nand GNAME18135(G18135,G18122,G14956);
  nand GNAME18136(G18136,G17182,G15099);
  nand GNAME18137(G18137,G14958,G15100);
  nand GNAME18138(G18138,G1683,G15096);
  nand GNAME18139(G18139,G18131,G59884);
  nand GNAME18140(G18140,G18127,G1680);
  nand GNAME18141(G18141,G18122,G14960);
  nand GNAME18142(G18142,G17204,G15099);
  nand GNAME18143(G18143,G14961,G15100);
  nand GNAME18144(G18144,G1682,G15096);
  nand GNAME18145(G18145,G18131,G59883);
  nand GNAME18146(G18146,G18127,G1669);
  nand GNAME18147(G18147,G18122,G14962);
  nand GNAME18148(G18148,G17213,G15099);
  nand GNAME18149(G18149,G14963,G15100);
  nand GNAME18150(G18150,G1681,G15096);
  nand GNAME18151(G18151,G18131,G59882);
  nand GNAME18152(G18152,G18127,G1666);
  nand GNAME18153(G18153,G18122,G14964);
  nand GNAME18154(G18154,G17222,G15099);
  nand GNAME18155(G18155,G14965,G15100);
  nand GNAME18156(G18156,G1679,G15096);
  nand GNAME18157(G18157,G18131,G59881);
  nand GNAME18158(G18158,G18127,G1665);
  nand GNAME18159(G18159,G18122,G14966);
  nand GNAME18160(G18160,G17231,G15099);
  nand GNAME18161(G18161,G14967,G15100);
  nand GNAME18162(G18162,G1678,G15096);
  nand GNAME18163(G18163,G18131,G59880);
  nand GNAME18164(G18164,G18127,G1664);
  nand GNAME18165(G18165,G18122,G14968);
  nand GNAME18166(G18166,G17240,G15099);
  nand GNAME18167(G18167,G14969,G15100);
  nand GNAME18168(G18168,G1677,G15096);
  nand GNAME18169(G18169,G18131,G59879);
  nand GNAME18170(G18170,G18127,G1663);
  nand GNAME18171(G18171,G18122,G14970);
  nand GNAME18172(G18172,G17249,G15099);
  nand GNAME18173(G18173,G14971,G15100);
  nand GNAME18174(G18174,G1676,G15096);
  nand GNAME18175(G18175,G18131,G59878);
  nand GNAME18176(G18176,G18127,G1662);
  nand GNAME18177(G18177,G18122,G14972);
  nand GNAME18178(G18178,G17258,G15099);
  nand GNAME18179(G18179,G14973,G15100);
  nand GNAME18180(G18180,G15102,G14791,G14796);
  or GNAME18181(G18181,G60244,G60245);
  nand GNAME18182(G18182,G14798,G18180);
  nand GNAME18183(G18183,G14786,G14783);
  nand GNAME18184(G18184,G14811,G15103);
  nand GNAME18185(G18185,G1589,G59876);
  nand GNAME18186(G18186,G14832,G15952,G15974);
  nand GNAME18187(G18187,G59874,G23088,G14799);
  nand GNAME18188(G18188,G14784,G18187);
  or GNAME18189(G18189,G15103,G15795);
  nand GNAME18190(G18190,G23088,G14904);
  nand GNAME18191(G18191,G18190,G18188,G18189);
  nand GNAME18192(G18192,G15105,G14746,G59877);
  nand GNAME18193(G18193,G18192,G15801);
  nand GNAME18194(G18194,G15807,G15104);
  nand GNAME18195(G18195,G18194,G59876);
  nand GNAME18196(G18196,G15104,G18193);
  nand GNAME18197(G18197,G14836,G14746,G59876);
  nand GNAME18198(G18198,G14784,G14937);
  or GNAME18199(G18199,G14831,G15104);
  or GNAME18200(G18200,G59839,G59841);
  nand GNAME18201(G18201,G18200,G15768);
  nand GNAME18202(G18202,G14745,G60247);
  nand GNAME18203(G18203,G14803,G34);
  nand GNAME18204(G18204,G60247,G15107,G18203);
  or GNAME18205(G18205,G14746,G14802);
  nand GNAME18206(G18206,G14746,G59839);
  or GNAME18207(G18207,G1589,G33);
  nand GNAME18208(G18208,G14809,G59839);
  nand GNAME18209(G18209,G14745,G18202);
  nand GNAME18210(G18210,G59841,G15106,G18209);
  nand GNAME18211(G18211,G18210,G14814);
  or GNAME18212(G18212,G15107,G14809,G14745);
  nand GNAME18213(G18213,G15781,G59838);
  nand GNAME18214(G18214,G60209,G15108);
  nand GNAME18215(G18215,G60208,G15109);
  nand GNAME18216(G18216,G15781,G59837);
  nand GNAME18217(G18217,G60209,G15109);
  nand GNAME18218(G18218,G60210,G15108);
  nand GNAME18219(G18219,G15781,G59836);
  nand GNAME18220(G18220,G60210,G15109);
  nand GNAME18221(G18221,G60211,G15108);
  nand GNAME18222(G18222,G15781,G59835);
  nand GNAME18223(G18223,G60211,G15109);
  nand GNAME18224(G18224,G60212,G15108);
  nand GNAME18225(G18225,G15781,G59834);
  nand GNAME18226(G18226,G60212,G15109);
  nand GNAME18227(G18227,G60213,G15108);
  nand GNAME18228(G18228,G15781,G59833);
  nand GNAME18229(G18229,G60213,G15109);
  nand GNAME18230(G18230,G60214,G15108);
  nand GNAME18231(G18231,G15781,G59832);
  nand GNAME18232(G18232,G60214,G15109);
  nand GNAME18233(G18233,G60215,G15108);
  nand GNAME18234(G18234,G15781,G59831);
  nand GNAME18235(G18235,G60215,G15109);
  nand GNAME18236(G18236,G60216,G15108);
  nand GNAME18237(G18237,G15781,G59830);
  nand GNAME18238(G18238,G60216,G15109);
  nand GNAME18239(G18239,G60217,G15108);
  nand GNAME18240(G18240,G15781,G59829);
  nand GNAME18241(G18241,G60217,G15109);
  nand GNAME18242(G18242,G60218,G15108);
  nand GNAME18243(G18243,G15781,G59828);
  nand GNAME18244(G18244,G60218,G15109);
  nand GNAME18245(G18245,G60219,G15108);
  nand GNAME18246(G18246,G15781,G59827);
  nand GNAME18247(G18247,G60219,G15109);
  nand GNAME18248(G18248,G60220,G15108);
  nand GNAME18249(G18249,G15781,G59826);
  nand GNAME18250(G18250,G60220,G15109);
  nand GNAME18251(G18251,G60221,G15108);
  nand GNAME18252(G18252,G15781,G59825);
  nand GNAME18253(G18253,G60221,G15109);
  nand GNAME18254(G18254,G60222,G15108);
  nand GNAME18255(G18255,G15781,G59824);
  nand GNAME18256(G18256,G60222,G15109);
  nand GNAME18257(G18257,G60223,G15108);
  nand GNAME18258(G18258,G15781,G59823);
  nand GNAME18259(G18259,G60223,G15109);
  nand GNAME18260(G18260,G60224,G15108);
  nand GNAME18261(G18261,G15781,G59822);
  nand GNAME18262(G18262,G60224,G15109);
  nand GNAME18263(G18263,G60225,G15108);
  nand GNAME18264(G18264,G15781,G59821);
  nand GNAME18265(G18265,G60225,G15109);
  nand GNAME18266(G18266,G60226,G15108);
  nand GNAME18267(G18267,G15781,G59820);
  nand GNAME18268(G18268,G60226,G15109);
  nand GNAME18269(G18269,G60227,G15108);
  nand GNAME18270(G18270,G15781,G59819);
  nand GNAME18271(G18271,G60227,G15109);
  nand GNAME18272(G18272,G60228,G15108);
  nand GNAME18273(G18273,G15781,G59818);
  nand GNAME18274(G18274,G60228,G15109);
  nand GNAME18275(G18275,G60229,G15108);
  nand GNAME18276(G18276,G15781,G59817);
  nand GNAME18277(G18277,G60229,G15109);
  nand GNAME18278(G18278,G60230,G15108);
  nand GNAME18279(G18279,G15781,G59816);
  nand GNAME18280(G18280,G60230,G15109);
  nand GNAME18281(G18281,G60231,G15108);
  nand GNAME18282(G18282,G15781,G59815);
  nand GNAME18283(G18283,G60231,G15109);
  nand GNAME18284(G18284,G60232,G15108);
  nand GNAME18285(G18285,G15781,G59814);
  nand GNAME18286(G18286,G60232,G15109);
  nand GNAME18287(G18287,G60233,G15108);
  nand GNAME18288(G18288,G15781,G59813);
  nand GNAME18289(G18289,G60233,G15109);
  nand GNAME18290(G18290,G60234,G15108);
  nand GNAME18291(G18291,G15781,G59812);
  nand GNAME18292(G18292,G60234,G15109);
  nand GNAME18293(G18293,G60235,G15108);
  nand GNAME18294(G18294,G15781,G59811);
  nand GNAME18295(G18295,G60235,G15109);
  nand GNAME18296(G18296,G60236,G15108);
  nand GNAME18297(G18297,G15781,G59810);
  nand GNAME18298(G18298,G60236,G15109);
  nand GNAME18299(G18299,G60237,G15108);
  nand GNAME18300(G18300,G15781,G59809);
  nand GNAME18301(G18301,G60237,G15109);
  nand GNAME18302(G18302,G60238,G15108);
  nand GNAME18303(G18303,G59990,G15112);
  nand GNAME18304(G18304,G59982,G15115);
  nand GNAME18305(G18305,G59974,G15116);
  nand GNAME18306(G18306,G59966,G15118);
  nand GNAME18307(G18307,G59958,G15119);
  nand GNAME18308(G18308,G59950,G15121);
  nand GNAME18309(G18309,G59942,G15122);
  nand GNAME18310(G18310,G59934,G15124);
  nand GNAME18311(G18311,G59926,G15126);
  nand GNAME18312(G18312,G59918,G15127);
  nand GNAME18313(G18313,G59910,G15128);
  nand GNAME18314(G18314,G59902,G15129);
  nand GNAME18315(G18315,G59894,G15130);
  nand GNAME18316(G18316,G59886,G15131);
  nand GNAME18317(G18317,G59878,G15132);
  nand GNAME18318(G18318,G59998,G15133);
  nand GNAME18319(G18319,G59991,G15112);
  nand GNAME18320(G18320,G59983,G15115);
  nand GNAME18321(G18321,G59975,G15116);
  nand GNAME18322(G18322,G59967,G15118);
  nand GNAME18323(G18323,G59959,G15119);
  nand GNAME18324(G18324,G59951,G15121);
  nand GNAME18325(G18325,G59943,G15122);
  nand GNAME18326(G18326,G59935,G15124);
  nand GNAME18327(G18327,G59927,G15126);
  nand GNAME18328(G18328,G59919,G15127);
  nand GNAME18329(G18329,G59911,G15128);
  nand GNAME18330(G18330,G59903,G15129);
  nand GNAME18331(G18331,G59895,G15130);
  nand GNAME18332(G18332,G59887,G15131);
  nand GNAME18333(G18333,G59879,G15132);
  nand GNAME18334(G18334,G59999,G15133);
  nand GNAME18335(G18335,G59992,G15112);
  nand GNAME18336(G18336,G59984,G15115);
  nand GNAME18337(G18337,G59976,G15116);
  nand GNAME18338(G18338,G59968,G15118);
  nand GNAME18339(G18339,G59960,G15119);
  nand GNAME18340(G18340,G59952,G15121);
  nand GNAME18341(G18341,G59944,G15122);
  nand GNAME18342(G18342,G59936,G15124);
  nand GNAME18343(G18343,G59928,G15126);
  nand GNAME18344(G18344,G59920,G15127);
  nand GNAME18345(G18345,G59912,G15128);
  nand GNAME18346(G18346,G59904,G15129);
  nand GNAME18347(G18347,G59896,G15130);
  nand GNAME18348(G18348,G59888,G15131);
  nand GNAME18349(G18349,G59880,G15132);
  nand GNAME18350(G18350,G60000,G15133);
  nand GNAME18351(G18351,G59993,G15112);
  nand GNAME18352(G18352,G59985,G15115);
  nand GNAME18353(G18353,G59977,G15116);
  nand GNAME18354(G18354,G59969,G15118);
  nand GNAME18355(G18355,G59961,G15119);
  nand GNAME18356(G18356,G59953,G15121);
  nand GNAME18357(G18357,G59945,G15122);
  nand GNAME18358(G18358,G59937,G15124);
  nand GNAME18359(G18359,G59929,G15126);
  nand GNAME18360(G18360,G59921,G15127);
  nand GNAME18361(G18361,G59913,G15128);
  nand GNAME18362(G18362,G59905,G15129);
  nand GNAME18363(G18363,G59897,G15130);
  nand GNAME18364(G18364,G59889,G15131);
  nand GNAME18365(G18365,G59881,G15132);
  nand GNAME18366(G18366,G60001,G15133);
  nand GNAME18367(G18367,G59994,G15112);
  nand GNAME18368(G18368,G59986,G15115);
  nand GNAME18369(G18369,G59978,G15116);
  nand GNAME18370(G18370,G59970,G15118);
  nand GNAME18371(G18371,G59962,G15119);
  nand GNAME18372(G18372,G59954,G15121);
  nand GNAME18373(G18373,G59946,G15122);
  nand GNAME18374(G18374,G59938,G15124);
  nand GNAME18375(G18375,G59930,G15126);
  nand GNAME18376(G18376,G59922,G15127);
  nand GNAME18377(G18377,G59914,G15128);
  nand GNAME18378(G18378,G59906,G15129);
  nand GNAME18379(G18379,G59898,G15130);
  nand GNAME18380(G18380,G59890,G15131);
  nand GNAME18381(G18381,G59882,G15132);
  nand GNAME18382(G18382,G60002,G15133);
  nand GNAME18383(G18383,G60003,G15133);
  nand GNAME18384(G18384,G59995,G15112);
  nand GNAME18385(G18385,G59987,G15115);
  nand GNAME18386(G18386,G59979,G15116);
  nand GNAME18387(G18387,G59971,G15118);
  nand GNAME18388(G18388,G59963,G15119);
  nand GNAME18389(G18389,G59955,G15121);
  nand GNAME18390(G18390,G59947,G15122);
  nand GNAME18391(G18391,G59939,G15124);
  nand GNAME18392(G18392,G59931,G15126);
  nand GNAME18393(G18393,G59923,G15127);
  nand GNAME18394(G18394,G59915,G15128);
  nand GNAME18395(G18395,G59907,G15129);
  nand GNAME18396(G18396,G59899,G15130);
  nand GNAME18397(G18397,G59891,G15131);
  nand GNAME18398(G18398,G59883,G15132);
  nand GNAME18399(G18399,G60004,G15133);
  nand GNAME18400(G18400,G59996,G15112);
  nand GNAME18401(G18401,G59988,G15115);
  nand GNAME18402(G18402,G59980,G15116);
  nand GNAME18403(G18403,G59972,G15118);
  nand GNAME18404(G18404,G59964,G15119);
  nand GNAME18405(G18405,G59956,G15121);
  nand GNAME18406(G18406,G59948,G15122);
  nand GNAME18407(G18407,G59940,G15124);
  nand GNAME18408(G18408,G59932,G15126);
  nand GNAME18409(G18409,G59924,G15127);
  nand GNAME18410(G18410,G59916,G15128);
  nand GNAME18411(G18411,G59908,G15129);
  nand GNAME18412(G18412,G59900,G15130);
  nand GNAME18413(G18413,G59892,G15131);
  nand GNAME18414(G18414,G59884,G15132);
  nand GNAME18415(G18415,G60005,G15133);
  nand GNAME18416(G18416,G59997,G15112);
  nand GNAME18417(G18417,G59989,G15115);
  nand GNAME18418(G18418,G59981,G15116);
  nand GNAME18419(G18419,G59973,G15118);
  nand GNAME18420(G18420,G59965,G15119);
  nand GNAME18421(G18421,G59957,G15121);
  nand GNAME18422(G18422,G59949,G15122);
  nand GNAME18423(G18423,G59941,G15124);
  nand GNAME18424(G18424,G59933,G15126);
  nand GNAME18425(G18425,G59925,G15127);
  nand GNAME18426(G18426,G59917,G15128);
  nand GNAME18427(G18427,G59909,G15129);
  nand GNAME18428(G18428,G59901,G15130);
  nand GNAME18429(G18429,G59893,G15131);
  nand GNAME18430(G18430,G59885,G15132);
  not GNAME18431(G18431,G15134);
  nand GNAME18432(G18432,G59990,G15136);
  nand GNAME18433(G18433,G59982,G15137);
  nand GNAME18434(G18434,G59974,G15138);
  nand GNAME18435(G18435,G59966,G15140);
  nand GNAME18436(G18436,G59958,G15141);
  nand GNAME18437(G18437,G59950,G15142);
  nand GNAME18438(G18438,G59942,G15143);
  nand GNAME18439(G18439,G59934,G15145);
  nand GNAME18440(G18440,G59926,G15146);
  nand GNAME18441(G18441,G59918,G15147);
  nand GNAME18442(G18442,G59910,G15148);
  nand GNAME18443(G18443,G59902,G15150);
  nand GNAME18444(G18444,G59894,G15151);
  nand GNAME18445(G18445,G59886,G15152);
  nand GNAME18446(G18446,G59878,G15153);
  nand GNAME18447(G18447,G59998,G15154);
  nand GNAME18448(G18448,G59991,G15136);
  nand GNAME18449(G18449,G59983,G15137);
  nand GNAME18450(G18450,G59975,G15138);
  nand GNAME18451(G18451,G59967,G15140);
  nand GNAME18452(G18452,G59959,G15141);
  nand GNAME18453(G18453,G59951,G15142);
  nand GNAME18454(G18454,G59943,G15143);
  nand GNAME18455(G18455,G59935,G15145);
  nand GNAME18456(G18456,G59927,G15146);
  nand GNAME18457(G18457,G59919,G15147);
  nand GNAME18458(G18458,G59911,G15148);
  nand GNAME18459(G18459,G59903,G15150);
  nand GNAME18460(G18460,G59895,G15151);
  nand GNAME18461(G18461,G59887,G15152);
  nand GNAME18462(G18462,G59879,G15153);
  nand GNAME18463(G18463,G59999,G15154);
  nand GNAME18464(G18464,G59992,G15136);
  nand GNAME18465(G18465,G59984,G15137);
  nand GNAME18466(G18466,G59976,G15138);
  nand GNAME18467(G18467,G59968,G15140);
  nand GNAME18468(G18468,G59960,G15141);
  nand GNAME18469(G18469,G59952,G15142);
  nand GNAME18470(G18470,G59944,G15143);
  nand GNAME18471(G18471,G59936,G15145);
  nand GNAME18472(G18472,G59928,G15146);
  nand GNAME18473(G18473,G59920,G15147);
  nand GNAME18474(G18474,G59912,G15148);
  nand GNAME18475(G18475,G59904,G15150);
  nand GNAME18476(G18476,G59896,G15151);
  nand GNAME18477(G18477,G59888,G15152);
  nand GNAME18478(G18478,G59880,G15153);
  nand GNAME18479(G18479,G60000,G15154);
  nand GNAME18480(G18480,G59993,G15136);
  nand GNAME18481(G18481,G59985,G15137);
  nand GNAME18482(G18482,G59977,G15138);
  nand GNAME18483(G18483,G59969,G15140);
  nand GNAME18484(G18484,G59961,G15141);
  nand GNAME18485(G18485,G59953,G15142);
  nand GNAME18486(G18486,G59945,G15143);
  nand GNAME18487(G18487,G59937,G15145);
  nand GNAME18488(G18488,G59929,G15146);
  nand GNAME18489(G18489,G59921,G15147);
  nand GNAME18490(G18490,G59913,G15148);
  nand GNAME18491(G18491,G59905,G15150);
  nand GNAME18492(G18492,G59897,G15151);
  nand GNAME18493(G18493,G59889,G15152);
  nand GNAME18494(G18494,G59881,G15153);
  nand GNAME18495(G18495,G60001,G15154);
  nand GNAME18496(G18496,G59994,G15136);
  nand GNAME18497(G18497,G59986,G15137);
  nand GNAME18498(G18498,G59978,G15138);
  nand GNAME18499(G18499,G59970,G15140);
  nand GNAME18500(G18500,G59962,G15141);
  nand GNAME18501(G18501,G59954,G15142);
  nand GNAME18502(G18502,G59946,G15143);
  nand GNAME18503(G18503,G59938,G15145);
  nand GNAME18504(G18504,G59930,G15146);
  nand GNAME18505(G18505,G59922,G15147);
  nand GNAME18506(G18506,G59914,G15148);
  nand GNAME18507(G18507,G59906,G15150);
  nand GNAME18508(G18508,G59898,G15151);
  nand GNAME18509(G18509,G59890,G15152);
  nand GNAME18510(G18510,G59882,G15153);
  nand GNAME18511(G18511,G60002,G15154);
  nand GNAME18512(G18512,G60003,G15154);
  nand GNAME18513(G18513,G59995,G15136);
  nand GNAME18514(G18514,G59987,G15137);
  nand GNAME18515(G18515,G59979,G15138);
  nand GNAME18516(G18516,G59971,G15140);
  nand GNAME18517(G18517,G59963,G15141);
  nand GNAME18518(G18518,G59955,G15142);
  nand GNAME18519(G18519,G59947,G15143);
  nand GNAME18520(G18520,G59939,G15145);
  nand GNAME18521(G18521,G59931,G15146);
  nand GNAME18522(G18522,G59923,G15147);
  nand GNAME18523(G18523,G59915,G15148);
  nand GNAME18524(G18524,G59907,G15150);
  nand GNAME18525(G18525,G59899,G15151);
  nand GNAME18526(G18526,G59891,G15152);
  nand GNAME18527(G18527,G59883,G15153);
  nand GNAME18528(G18528,G60004,G15154);
  nand GNAME18529(G18529,G59996,G15136);
  nand GNAME18530(G18530,G59988,G15137);
  nand GNAME18531(G18531,G59980,G15138);
  nand GNAME18532(G18532,G59972,G15140);
  nand GNAME18533(G18533,G59964,G15141);
  nand GNAME18534(G18534,G59956,G15142);
  nand GNAME18535(G18535,G59948,G15143);
  nand GNAME18536(G18536,G59940,G15145);
  nand GNAME18537(G18537,G59932,G15146);
  nand GNAME18538(G18538,G59924,G15147);
  nand GNAME18539(G18539,G59916,G15148);
  nand GNAME18540(G18540,G59908,G15150);
  nand GNAME18541(G18541,G59900,G15151);
  nand GNAME18542(G18542,G59892,G15152);
  nand GNAME18543(G18543,G59884,G15153);
  nand GNAME18544(G18544,G60005,G15154);
  nand GNAME18545(G18545,G59997,G15136);
  nand GNAME18546(G18546,G59989,G15137);
  nand GNAME18547(G18547,G59981,G15138);
  nand GNAME18548(G18548,G59973,G15140);
  nand GNAME18549(G18549,G59965,G15141);
  nand GNAME18550(G18550,G59957,G15142);
  nand GNAME18551(G18551,G59949,G15143);
  nand GNAME18552(G18552,G59941,G15145);
  nand GNAME18553(G18553,G59933,G15146);
  nand GNAME18554(G18554,G59925,G15147);
  nand GNAME18555(G18555,G59917,G15148);
  nand GNAME18556(G18556,G59909,G15150);
  nand GNAME18557(G18557,G59901,G15151);
  nand GNAME18558(G18558,G59893,G15152);
  nand GNAME18559(G18559,G59885,G15153);
  nand GNAME18560(G18560,G59990,G14984);
  nand GNAME18561(G18561,G59982,G14995);
  nand GNAME18562(G18562,G59974,G15003);
  nand GNAME18563(G18563,G59966,G15013);
  nand GNAME18564(G18564,G59958,G15022);
  nand GNAME18565(G18565,G59950,G15029);
  nand GNAME18566(G18566,G59942,G15036);
  nand GNAME18567(G18567,G59934,G15047);
  nand GNAME18568(G18568,G59926,G15054);
  nand GNAME18569(G18569,G59918,G15063);
  nand GNAME18570(G18570,G59910,G15070);
  nand GNAME18571(G18571,G59902,G15079);
  nand GNAME18572(G18572,G59894,G15086);
  nand GNAME18573(G18573,G59886,G15093);
  nand GNAME18574(G18574,G59878,G15100);
  nand GNAME18575(G18575,G59998,G14957);
  nand GNAME18576(G18576,G15594,G15595,G15596,G15597);
  nand GNAME18577(G18577,G59991,G14984);
  nand GNAME18578(G18578,G59983,G14995);
  nand GNAME18579(G18579,G59975,G15003);
  nand GNAME18580(G18580,G59967,G15013);
  nand GNAME18581(G18581,G59959,G15022);
  nand GNAME18582(G18582,G59951,G15029);
  nand GNAME18583(G18583,G59943,G15036);
  nand GNAME18584(G18584,G59935,G15047);
  nand GNAME18585(G18585,G59927,G15054);
  nand GNAME18586(G18586,G59919,G15063);
  nand GNAME18587(G18587,G59911,G15070);
  nand GNAME18588(G18588,G59903,G15079);
  nand GNAME18589(G18589,G59895,G15086);
  nand GNAME18590(G18590,G59887,G15093);
  nand GNAME18591(G18591,G59879,G15100);
  nand GNAME18592(G18592,G59999,G14957);
  nand GNAME18593(G18593,G15598,G15599,G15600,G15601);
  nand GNAME18594(G18594,G59992,G14984);
  nand GNAME18595(G18595,G59984,G14995);
  nand GNAME18596(G18596,G59976,G15003);
  nand GNAME18597(G18597,G59968,G15013);
  nand GNAME18598(G18598,G59960,G15022);
  nand GNAME18599(G18599,G59952,G15029);
  nand GNAME18600(G18600,G59944,G15036);
  nand GNAME18601(G18601,G59936,G15047);
  nand GNAME18602(G18602,G59928,G15054);
  nand GNAME18603(G18603,G59920,G15063);
  nand GNAME18604(G18604,G59912,G15070);
  nand GNAME18605(G18605,G59904,G15079);
  nand GNAME18606(G18606,G59896,G15086);
  nand GNAME18607(G18607,G59888,G15093);
  nand GNAME18608(G18608,G59880,G15100);
  nand GNAME18609(G18609,G60000,G14957);
  nand GNAME18610(G18610,G15602,G15603,G15604,G15605);
  nand GNAME18611(G18611,G59993,G14984);
  nand GNAME18612(G18612,G59985,G14995);
  nand GNAME18613(G18613,G59977,G15003);
  nand GNAME18614(G18614,G59969,G15013);
  nand GNAME18615(G18615,G59961,G15022);
  nand GNAME18616(G18616,G59953,G15029);
  nand GNAME18617(G18617,G59945,G15036);
  nand GNAME18618(G18618,G59937,G15047);
  nand GNAME18619(G18619,G59929,G15054);
  nand GNAME18620(G18620,G59921,G15063);
  nand GNAME18621(G18621,G59913,G15070);
  nand GNAME18622(G18622,G59905,G15079);
  nand GNAME18623(G18623,G59897,G15086);
  nand GNAME18624(G18624,G59889,G15093);
  nand GNAME18625(G18625,G59881,G15100);
  nand GNAME18626(G18626,G60001,G14957);
  nand GNAME18627(G18627,G15606,G15607,G15608,G15609);
  nand GNAME18628(G18628,G59994,G14984);
  nand GNAME18629(G18629,G59986,G14995);
  nand GNAME18630(G18630,G59978,G15003);
  nand GNAME18631(G18631,G59970,G15013);
  nand GNAME18632(G18632,G59962,G15022);
  nand GNAME18633(G18633,G59954,G15029);
  nand GNAME18634(G18634,G59946,G15036);
  nand GNAME18635(G18635,G59938,G15047);
  nand GNAME18636(G18636,G59930,G15054);
  nand GNAME18637(G18637,G59922,G15063);
  nand GNAME18638(G18638,G59914,G15070);
  nand GNAME18639(G18639,G59906,G15079);
  nand GNAME18640(G18640,G59898,G15086);
  nand GNAME18641(G18641,G59890,G15093);
  nand GNAME18642(G18642,G59882,G15100);
  nand GNAME18643(G18643,G60002,G14957);
  nand GNAME18644(G18644,G15610,G15611,G15612,G15613);
  nand GNAME18645(G18645,G60003,G14957);
  nand GNAME18646(G18646,G59995,G14984);
  nand GNAME18647(G18647,G59987,G14995);
  nand GNAME18648(G18648,G59979,G15003);
  nand GNAME18649(G18649,G59971,G15013);
  nand GNAME18650(G18650,G59963,G15022);
  nand GNAME18651(G18651,G59955,G15029);
  nand GNAME18652(G18652,G59947,G15036);
  nand GNAME18653(G18653,G59939,G15047);
  nand GNAME18654(G18654,G59931,G15054);
  nand GNAME18655(G18655,G59923,G15063);
  nand GNAME18656(G18656,G59915,G15070);
  nand GNAME18657(G18657,G59907,G15079);
  nand GNAME18658(G18658,G59899,G15086);
  nand GNAME18659(G18659,G59891,G15093);
  nand GNAME18660(G18660,G59883,G15100);
  nand GNAME18661(G18661,G15614,G15615,G15616,G15617);
  nand GNAME18662(G18662,G60004,G14957);
  nand GNAME18663(G18663,G59996,G14984);
  nand GNAME18664(G18664,G59988,G14995);
  nand GNAME18665(G18665,G59980,G15003);
  nand GNAME18666(G18666,G59972,G15013);
  nand GNAME18667(G18667,G59964,G15022);
  nand GNAME18668(G18668,G59956,G15029);
  nand GNAME18669(G18669,G59948,G15036);
  nand GNAME18670(G18670,G59940,G15047);
  nand GNAME18671(G18671,G59932,G15054);
  nand GNAME18672(G18672,G59924,G15063);
  nand GNAME18673(G18673,G59916,G15070);
  nand GNAME18674(G18674,G59908,G15079);
  nand GNAME18675(G18675,G59900,G15086);
  nand GNAME18676(G18676,G59892,G15093);
  nand GNAME18677(G18677,G59884,G15100);
  nand GNAME18678(G18678,G15618,G15619,G15620,G15621);
  nand GNAME18679(G18679,G60005,G14957);
  nand GNAME18680(G18680,G59997,G14984);
  nand GNAME18681(G18681,G59989,G14995);
  nand GNAME18682(G18682,G59981,G15003);
  nand GNAME18683(G18683,G59973,G15013);
  nand GNAME18684(G18684,G59965,G15022);
  nand GNAME18685(G18685,G59957,G15029);
  nand GNAME18686(G18686,G59949,G15036);
  nand GNAME18687(G18687,G59941,G15047);
  nand GNAME18688(G18688,G59933,G15054);
  nand GNAME18689(G18689,G59925,G15063);
  nand GNAME18690(G18690,G59917,G15070);
  nand GNAME18691(G18691,G59909,G15079);
  nand GNAME18692(G18692,G59901,G15086);
  nand GNAME18693(G18693,G59893,G15093);
  nand GNAME18694(G18694,G59885,G15100);
  nand GNAME18695(G18695,G15622,G15623,G15624,G15625);
  nand GNAME18696(G18696,G59990,G15157);
  nand GNAME18697(G18697,G59982,G15160);
  nand GNAME18698(G18698,G59974,G15162);
  nand GNAME18699(G18699,G59966,G15165);
  nand GNAME18700(G18700,G59958,G15166);
  nand GNAME18701(G18701,G59950,G15167);
  nand GNAME18702(G18702,G59942,G15168);
  nand GNAME18703(G18703,G59934,G15170);
  nand GNAME18704(G18704,G59926,G15171);
  nand GNAME18705(G18705,G59918,G15172);
  nand GNAME18706(G18706,G59910,G15173);
  nand GNAME18707(G18707,G59902,G15175);
  nand GNAME18708(G18708,G59894,G15176);
  nand GNAME18709(G18709,G59886,G15177);
  nand GNAME18710(G18710,G59878,G15178);
  nand GNAME18711(G18711,G59998,G15179);
  nand GNAME18712(G18712,G15626,G15627,G15628,G15629);
  nand GNAME18713(G18713,G59991,G15157);
  nand GNAME18714(G18714,G59983,G15160);
  nand GNAME18715(G18715,G59975,G15162);
  nand GNAME18716(G18716,G59967,G15165);
  nand GNAME18717(G18717,G59959,G15166);
  nand GNAME18718(G18718,G59951,G15167);
  nand GNAME18719(G18719,G59943,G15168);
  nand GNAME18720(G18720,G59935,G15170);
  nand GNAME18721(G18721,G59927,G15171);
  nand GNAME18722(G18722,G59919,G15172);
  nand GNAME18723(G18723,G59911,G15173);
  nand GNAME18724(G18724,G59903,G15175);
  nand GNAME18725(G18725,G59895,G15176);
  nand GNAME18726(G18726,G59887,G15177);
  nand GNAME18727(G18727,G59879,G15178);
  nand GNAME18728(G18728,G59999,G15179);
  nand GNAME18729(G18729,G15630,G15631,G15632,G15633);
  nand GNAME18730(G18730,G59992,G15157);
  nand GNAME18731(G18731,G59984,G15160);
  nand GNAME18732(G18732,G59976,G15162);
  nand GNAME18733(G18733,G59968,G15165);
  nand GNAME18734(G18734,G59960,G15166);
  nand GNAME18735(G18735,G59952,G15167);
  nand GNAME18736(G18736,G59944,G15168);
  nand GNAME18737(G18737,G59936,G15170);
  nand GNAME18738(G18738,G59928,G15171);
  nand GNAME18739(G18739,G59920,G15172);
  nand GNAME18740(G18740,G59912,G15173);
  nand GNAME18741(G18741,G59904,G15175);
  nand GNAME18742(G18742,G59896,G15176);
  nand GNAME18743(G18743,G59888,G15177);
  nand GNAME18744(G18744,G59880,G15178);
  nand GNAME18745(G18745,G60000,G15179);
  nand GNAME18746(G18746,G15634,G15635,G15636,G15637);
  nand GNAME18747(G18747,G59993,G15157);
  nand GNAME18748(G18748,G59985,G15160);
  nand GNAME18749(G18749,G59977,G15162);
  nand GNAME18750(G18750,G59969,G15165);
  nand GNAME18751(G18751,G59961,G15166);
  nand GNAME18752(G18752,G59953,G15167);
  nand GNAME18753(G18753,G59945,G15168);
  nand GNAME18754(G18754,G59937,G15170);
  nand GNAME18755(G18755,G59929,G15171);
  nand GNAME18756(G18756,G59921,G15172);
  nand GNAME18757(G18757,G59913,G15173);
  nand GNAME18758(G18758,G59905,G15175);
  nand GNAME18759(G18759,G59897,G15176);
  nand GNAME18760(G18760,G59889,G15177);
  nand GNAME18761(G18761,G59881,G15178);
  nand GNAME18762(G18762,G60001,G15179);
  nand GNAME18763(G18763,G15638,G15639,G15640,G15641);
  nand GNAME18764(G18764,G59994,G15157);
  nand GNAME18765(G18765,G59986,G15160);
  nand GNAME18766(G18766,G59978,G15162);
  nand GNAME18767(G18767,G59970,G15165);
  nand GNAME18768(G18768,G59962,G15166);
  nand GNAME18769(G18769,G59954,G15167);
  nand GNAME18770(G18770,G59946,G15168);
  nand GNAME18771(G18771,G59938,G15170);
  nand GNAME18772(G18772,G59930,G15171);
  nand GNAME18773(G18773,G59922,G15172);
  nand GNAME18774(G18774,G59914,G15173);
  nand GNAME18775(G18775,G59906,G15175);
  nand GNAME18776(G18776,G59898,G15176);
  nand GNAME18777(G18777,G59890,G15177);
  nand GNAME18778(G18778,G59882,G15178);
  nand GNAME18779(G18779,G60002,G15179);
  nand GNAME18780(G18780,G15642,G15643,G15644,G15645);
  nand GNAME18781(G18781,G60003,G15179);
  nand GNAME18782(G18782,G59995,G15157);
  nand GNAME18783(G18783,G59987,G15160);
  nand GNAME18784(G18784,G59979,G15162);
  nand GNAME18785(G18785,G59971,G15165);
  nand GNAME18786(G18786,G59963,G15166);
  nand GNAME18787(G18787,G59955,G15167);
  nand GNAME18788(G18788,G59947,G15168);
  nand GNAME18789(G18789,G59939,G15170);
  nand GNAME18790(G18790,G59931,G15171);
  nand GNAME18791(G18791,G59923,G15172);
  nand GNAME18792(G18792,G59915,G15173);
  nand GNAME18793(G18793,G59907,G15175);
  nand GNAME18794(G18794,G59899,G15176);
  nand GNAME18795(G18795,G59891,G15177);
  nand GNAME18796(G18796,G59883,G15178);
  nand GNAME18797(G18797,G15646,G15647,G15648,G15649);
  nand GNAME18798(G18798,G60004,G15179);
  nand GNAME18799(G18799,G59996,G15157);
  nand GNAME18800(G18800,G59988,G15160);
  nand GNAME18801(G18801,G59980,G15162);
  nand GNAME18802(G18802,G59972,G15165);
  nand GNAME18803(G18803,G59964,G15166);
  nand GNAME18804(G18804,G59956,G15167);
  nand GNAME18805(G18805,G59948,G15168);
  nand GNAME18806(G18806,G59940,G15170);
  nand GNAME18807(G18807,G59932,G15171);
  nand GNAME18808(G18808,G59924,G15172);
  nand GNAME18809(G18809,G59916,G15173);
  nand GNAME18810(G18810,G59908,G15175);
  nand GNAME18811(G18811,G59900,G15176);
  nand GNAME18812(G18812,G59892,G15177);
  nand GNAME18813(G18813,G59884,G15178);
  nand GNAME18814(G18814,G15650,G15651,G15652,G15653);
  nand GNAME18815(G18815,G60005,G15179);
  nand GNAME18816(G18816,G59997,G15157);
  nand GNAME18817(G18817,G59989,G15160);
  nand GNAME18818(G18818,G59981,G15162);
  nand GNAME18819(G18819,G59973,G15165);
  nand GNAME18820(G18820,G59965,G15166);
  nand GNAME18821(G18821,G59957,G15167);
  nand GNAME18822(G18822,G59949,G15168);
  nand GNAME18823(G18823,G59941,G15170);
  nand GNAME18824(G18824,G59933,G15171);
  nand GNAME18825(G18825,G59925,G15172);
  nand GNAME18826(G18826,G59917,G15173);
  nand GNAME18827(G18827,G59909,G15175);
  nand GNAME18828(G18828,G59901,G15176);
  nand GNAME18829(G18829,G59893,G15177);
  nand GNAME18830(G18830,G59885,G15178);
  nand GNAME18831(G18831,G15654,G15655,G15656,G15657);
  nand GNAME18832(G18832,G15802,G15779,G15788);
  or GNAME18833(G18833,G15233,G15234);
  nand GNAME18834(G18834,G14821,G20030);
  nand GNAME18835(G18835,G18833,G23461);
  nand GNAME18836(G18836,G18832,G60025);
  nand GNAME18837(G18837,G23199,G15181);
  nand GNAME18838(G18838,G60216,G15183);
  nand GNAME18839(G18839,G14821,G20029);
  nand GNAME18840(G18840,G18833,G23496);
  nand GNAME18841(G18841,G18832,G60024);
  nand GNAME18842(G18842,G23156,G15181);
  nand GNAME18843(G18843,G60215,G15183);
  nand GNAME18844(G18844,G14821,G23486);
  nand GNAME18845(G18845,G18833,G23486);
  nand GNAME18846(G18846,G18832,G60023);
  nand GNAME18847(G18847,G23157,G15181);
  nand GNAME18848(G18848,G60214,G15183);
  nand GNAME18849(G18849,G14821,G23428);
  nand GNAME18850(G18850,G18833,G23428);
  nand GNAME18851(G18851,G18832,G60022);
  nand GNAME18852(G18852,G23123,G15181);
  nand GNAME18853(G18853,G60213,G15183);
  nand GNAME18854(G18854,G14821,G23500);
  nand GNAME18855(G18855,G18833,G23500);
  nand GNAME18856(G18856,G18832,G60021);
  nand GNAME18857(G18857,G23158,G15181);
  nand GNAME18858(G18858,G60212,G15183);
  nand GNAME18859(G18859,G14821,G23503);
  nand GNAME18860(G18860,G18833,G23503);
  nand GNAME18861(G18861,G18832,G60020);
  nand GNAME18862(G18862,G23159,G15181);
  nand GNAME18863(G18863,G60211,G15183);
  nand GNAME18864(G18864,G18833,G23488);
  nand GNAME18865(G18865,G18832,G60047);
  nand GNAME18866(G18866,G23190,G15181);
  nand GNAME18867(G18867,G60238,G15183);
  nand GNAME18868(G18868,G14821,G20028);
  nand GNAME18869(G18869,G18833,G23427);
  nand GNAME18870(G18870,G18832,G60046);
  nand GNAME18871(G18871,G23122,G15181);
  nand GNAME18872(G18872,G60237,G15183);
  nand GNAME18873(G18873,G14821,G23487);
  nand GNAME18874(G18874,G18833,G23487);
  nand GNAME18875(G18875,G18832,G60019);
  nand GNAME18876(G18876,G60210,G15183);
  nand GNAME18877(G18877,G23160,G15181);
  nand GNAME18878(G18878,G14821,G20027);
  nand GNAME18879(G18879,G18833,G23475);
  nand GNAME18880(G18880,G18832,G60045);
  nand GNAME18881(G18881,G23176,G15181);
  nand GNAME18882(G18882,G60236,G15183);
  nand GNAME18883(G18883,G14821,G20026);
  nand GNAME18884(G18884,G18833,G23476);
  nand GNAME18885(G18885,G18832,G60044);
  nand GNAME18886(G18886,G23177,G15181);
  nand GNAME18887(G18887,G60235,G15183);
  nand GNAME18888(G18888,G14821,G20025);
  nand GNAME18889(G18889,G18833,G23477);
  nand GNAME18890(G18890,G18832,G60043);
  nand GNAME18891(G18891,G23178,G15181);
  nand GNAME18892(G18892,G60234,G15183);
  nand GNAME18893(G18893,G14821,G20024);
  nand GNAME18894(G18894,G18833,G23478);
  nand GNAME18895(G18895,G18832,G60042);
  nand GNAME18896(G18896,G23179,G15181);
  nand GNAME18897(G18897,G60233,G15183);
  nand GNAME18898(G18898,G14821,G20023);
  nand GNAME18899(G18899,G18833,G23479);
  nand GNAME18900(G18900,G18832,G60041);
  nand GNAME18901(G18901,G23180,G15181);
  nand GNAME18902(G18902,G60232,G15183);
  nand GNAME18903(G18903,G14821,G20022);
  nand GNAME18904(G18904,G18833,G23517);
  nand GNAME18905(G18905,G18832,G60040);
  nand GNAME18906(G18906,G23181,G15181);
  nand GNAME18907(G18907,G60231,G15183);
  nand GNAME18908(G18908,G14821,G20021);
  nand GNAME18909(G18909,G18833,G23520);
  nand GNAME18910(G18910,G18832,G60039);
  nand GNAME18911(G18911,G23182,G15181);
  nand GNAME18912(G18912,G60230,G15183);
  nand GNAME18913(G18913,G14821,G20020);
  nand GNAME18914(G18914,G18833,G23523);
  nand GNAME18915(G18915,G18832,G60038);
  nand GNAME18916(G18916,G23183,G15181);
  nand GNAME18917(G18917,G60229,G15183);
  nand GNAME18918(G18918,G14821,G20019);
  nand GNAME18919(G18919,G18833,G23526);
  nand GNAME18920(G18920,G18832,G60037);
  nand GNAME18921(G18921,G23184,G15181);
  nand GNAME18922(G18922,G60228,G15183);
  nand GNAME18923(G18923,G14821,G20018);
  nand GNAME18924(G18924,G18833,G23529);
  nand GNAME18925(G18925,G18832,G60036);
  nand GNAME18926(G18926,G23185,G15181);
  nand GNAME18927(G18927,G60227,G15183);
  nand GNAME18928(G18928,G14821,G23426);
  nand GNAME18929(G18929,G18833,G23426);
  nand GNAME18930(G18930,G18832,G60018);
  nand GNAME18931(G18931,G60209,G15183);
  nand GNAME18932(G18932,G23121,G15181);
  nand GNAME18933(G18933,G14821,G20017);
  nand GNAME18934(G18934,G18833,G23535);
  nand GNAME18935(G18935,G18832,G60035);
  nand GNAME18936(G18936,G23186,G15181);
  nand GNAME18937(G18937,G60226,G15183);
  nand GNAME18938(G18938,G14821,G20016);
  nand GNAME18939(G18939,G18833,G23538);
  nand GNAME18940(G18940,G18832,G60034);
  nand GNAME18941(G18941,G23187,G15181);
  nand GNAME18942(G18942,G60225,G15183);
  nand GNAME18943(G18943,G14821,G20015);
  nand GNAME18944(G18944,G18833,G23541);
  nand GNAME18945(G18945,G18832,G60033);
  nand GNAME18946(G18946,G23188,G15181);
  nand GNAME18947(G18947,G60224,G15183);
  nand GNAME18948(G18948,G14821,G20002);
  nand GNAME18949(G18949,G18833,G23480);
  nand GNAME18950(G18950,G18832,G60032);
  nand GNAME18951(G18951,G23216,G15181);
  nand GNAME18952(G18952,G60223,G15183);
  nand GNAME18953(G18953,G14821,G20065);
  nand GNAME18954(G18954,G18833,G23481);
  nand GNAME18955(G18955,G18832,G60031);
  nand GNAME18956(G18956,G23219,G15181);
  nand GNAME18957(G18957,G60222,G15183);
  nand GNAME18958(G18958,G14821,G20000);
  nand GNAME18959(G18959,G18833,G23425);
  nand GNAME18960(G18960,G18832,G60030);
  nand GNAME18961(G18961,G23191,G15181);
  nand GNAME18962(G18962,G60221,G15183);
  nand GNAME18963(G18963,G14821,G19999);
  nand GNAME18964(G18964,G18833,G23482);
  nand GNAME18965(G18965,G18832,G60029);
  nand GNAME18966(G18966,G23223,G15181);
  nand GNAME18967(G18967,G60220,G15183);
  nand GNAME18968(G18968,G14821,G19998);
  nand GNAME18969(G18969,G18833,G23483);
  nand GNAME18970(G18970,G18832,G60028);
  nand GNAME18971(G18971,G23226,G15181);
  nand GNAME18972(G18972,G60219,G15183);
  nand GNAME18973(G18973,G14821,G19997);
  nand GNAME18974(G18974,G18833,G23484);
  nand GNAME18975(G18975,G18832,G60027);
  nand GNAME18976(G18976,G23192,G15181);
  nand GNAME18977(G18977,G60218,G15183);
  nand GNAME18978(G18978,G14821,G19996);
  nand GNAME18979(G18979,G18833,G23424);
  nand GNAME18980(G18980,G18832,G60026);
  nand GNAME18981(G18981,G23120,G15181);
  nand GNAME18982(G18982,G60217,G15183);
  nand GNAME18983(G18983,G14821,G23532);
  nand GNAME18984(G18984,G18833,G23532);
  nand GNAME18985(G18985,G18832,G60017);
  nand GNAME18986(G18986,G23213,G15181);
  nand GNAME18987(G18987,G60208,G15183);
  nand GNAME18988(G18988,G14821,G23485);
  nand GNAME18989(G18989,G18833,G23485);
  nand GNAME18990(G18990,G18832,G60016);
  nand GNAME18991(G18991,G23189,G15181);
  nand GNAME18992(G18992,G60207,G15183);
  nand GNAME18993(G18993,G59990,G17265);
  nand GNAME18994(G18994,G59982,G17326);
  nand GNAME18995(G18995,G59974,G17387);
  nand GNAME18996(G18996,G59966,G17448);
  nand GNAME18997(G18997,G59958,G17509);
  nand GNAME18998(G18998,G59950,G17570);
  nand GNAME18999(G18999,G59942,G17631);
  nand GNAME19000(G19000,G59934,G17692);
  nand GNAME19001(G19001,G59926,G17753);
  nand GNAME19002(G19002,G59918,G17814);
  nand GNAME19003(G19003,G59910,G17875);
  nand GNAME19004(G19004,G59902,G17936);
  nand GNAME19005(G19005,G59894,G17997);
  nand GNAME19006(G19006,G59886,G18058);
  nand GNAME19007(G19007,G59878,G18119);
  nand GNAME19008(G19008,G59998,G17183);
  nand GNAME19009(G19009,G15667,G15668,G15669,G15670);
  nand GNAME19010(G19010,G59990,G15211);
  nand GNAME19011(G19011,G59982,G15213);
  nand GNAME19012(G19012,G59974,G15215);
  nand GNAME19013(G19013,G59966,G15218);
  nand GNAME19014(G19014,G59958,G15219);
  nand GNAME19015(G19015,G59950,G15220);
  nand GNAME19016(G19016,G59942,G15221);
  nand GNAME19017(G19017,G59934,G15223);
  nand GNAME19018(G19018,G59926,G15224);
  nand GNAME19019(G19019,G59918,G15225);
  nand GNAME19020(G19020,G59910,G15226);
  nand GNAME19021(G19021,G59902,G15228);
  nand GNAME19022(G19022,G59894,G15229);
  nand GNAME19023(G19023,G59886,G15230);
  nand GNAME19024(G19024,G59878,G15231);
  nand GNAME19025(G19025,G59998,G15232);
  nand GNAME19026(G19026,G15663,G15664,G15665,G15666);
  nand GNAME19027(G19027,G59990,G15187);
  nand GNAME19028(G19028,G59982,G15190);
  nand GNAME19029(G19029,G59974,G15191);
  nand GNAME19030(G19030,G59966,G15193);
  nand GNAME19031(G19031,G59958,G15195);
  nand GNAME19032(G19032,G59950,G15196);
  nand GNAME19033(G19033,G59942,G15197);
  nand GNAME19034(G19034,G59934,G15199);
  nand GNAME19035(G19035,G59926,G15200);
  nand GNAME19036(G19036,G59918,G15202);
  nand GNAME19037(G19037,G59910,G15203);
  nand GNAME19038(G19038,G59902,G15204);
  nand GNAME19039(G19039,G59894,G15205);
  nand GNAME19040(G19040,G59886,G15206);
  nand GNAME19041(G19041,G59878,G15207);
  nand GNAME19042(G19042,G59998,G15208);
  nand GNAME19043(G19043,G15659,G15660,G15661,G15662);
  nand GNAME19044(G19044,G15181,G23418);
  nand GNAME19045(G19045,G19043,G14821);
  nand GNAME19046(G19046,G19026,G15233);
  nand GNAME19047(G19047,G19009,G15234);
  nand GNAME19048(G19048,G59991,G17265);
  nand GNAME19049(G19049,G59983,G17326);
  nand GNAME19050(G19050,G59975,G17387);
  nand GNAME19051(G19051,G59967,G17448);
  nand GNAME19052(G19052,G59959,G17509);
  nand GNAME19053(G19053,G59951,G17570);
  nand GNAME19054(G19054,G59943,G17631);
  nand GNAME19055(G19055,G59935,G17692);
  nand GNAME19056(G19056,G59927,G17753);
  nand GNAME19057(G19057,G59919,G17814);
  nand GNAME19058(G19058,G59911,G17875);
  nand GNAME19059(G19059,G59903,G17936);
  nand GNAME19060(G19060,G59895,G17997);
  nand GNAME19061(G19061,G59887,G18058);
  nand GNAME19062(G19062,G59879,G18119);
  nand GNAME19063(G19063,G59999,G17183);
  nand GNAME19064(G19064,G15679,G15680,G15681,G15682);
  nand GNAME19065(G19065,G59991,G15211);
  nand GNAME19066(G19066,G59983,G15213);
  nand GNAME19067(G19067,G59975,G15215);
  nand GNAME19068(G19068,G59967,G15218);
  nand GNAME19069(G19069,G59959,G15219);
  nand GNAME19070(G19070,G59951,G15220);
  nand GNAME19071(G19071,G59943,G15221);
  nand GNAME19072(G19072,G59935,G15223);
  nand GNAME19073(G19073,G59927,G15224);
  nand GNAME19074(G19074,G59919,G15225);
  nand GNAME19075(G19075,G59911,G15226);
  nand GNAME19076(G19076,G59903,G15228);
  nand GNAME19077(G19077,G59895,G15229);
  nand GNAME19078(G19078,G59887,G15230);
  nand GNAME19079(G19079,G59879,G15231);
  nand GNAME19080(G19080,G59999,G15232);
  nand GNAME19081(G19081,G15675,G15676,G15677,G15678);
  nand GNAME19082(G19082,G59991,G15187);
  nand GNAME19083(G19083,G59983,G15190);
  nand GNAME19084(G19084,G59975,G15191);
  nand GNAME19085(G19085,G59967,G15193);
  nand GNAME19086(G19086,G59959,G15195);
  nand GNAME19087(G19087,G59951,G15196);
  nand GNAME19088(G19088,G59943,G15197);
  nand GNAME19089(G19089,G59935,G15199);
  nand GNAME19090(G19090,G59927,G15200);
  nand GNAME19091(G19091,G59919,G15202);
  nand GNAME19092(G19092,G59911,G15203);
  nand GNAME19093(G19093,G59903,G15204);
  nand GNAME19094(G19094,G59895,G15205);
  nand GNAME19095(G19095,G59887,G15206);
  nand GNAME19096(G19096,G59879,G15207);
  nand GNAME19097(G19097,G59999,G15208);
  nand GNAME19098(G19098,G15671,G15672,G15673,G15674);
  nand GNAME19099(G19099,G15181,G23416);
  nand GNAME19100(G19100,G19098,G14821);
  nand GNAME19101(G19101,G19081,G15233);
  nand GNAME19102(G19102,G19064,G15234);
  nand GNAME19103(G19103,G59992,G17265);
  nand GNAME19104(G19104,G59984,G17326);
  nand GNAME19105(G19105,G59976,G17387);
  nand GNAME19106(G19106,G59968,G17448);
  nand GNAME19107(G19107,G59960,G17509);
  nand GNAME19108(G19108,G59952,G17570);
  nand GNAME19109(G19109,G59944,G17631);
  nand GNAME19110(G19110,G59936,G17692);
  nand GNAME19111(G19111,G59928,G17753);
  nand GNAME19112(G19112,G59920,G17814);
  nand GNAME19113(G19113,G59912,G17875);
  nand GNAME19114(G19114,G59904,G17936);
  nand GNAME19115(G19115,G59896,G17997);
  nand GNAME19116(G19116,G59888,G18058);
  nand GNAME19117(G19117,G59880,G18119);
  nand GNAME19118(G19118,G60000,G17183);
  nand GNAME19119(G19119,G15691,G15692,G15693,G15694);
  nand GNAME19120(G19120,G59992,G15211);
  nand GNAME19121(G19121,G59984,G15213);
  nand GNAME19122(G19122,G59976,G15215);
  nand GNAME19123(G19123,G59968,G15218);
  nand GNAME19124(G19124,G59960,G15219);
  nand GNAME19125(G19125,G59952,G15220);
  nand GNAME19126(G19126,G59944,G15221);
  nand GNAME19127(G19127,G59936,G15223);
  nand GNAME19128(G19128,G59928,G15224);
  nand GNAME19129(G19129,G59920,G15225);
  nand GNAME19130(G19130,G59912,G15226);
  nand GNAME19131(G19131,G59904,G15228);
  nand GNAME19132(G19132,G59896,G15229);
  nand GNAME19133(G19133,G59888,G15230);
  nand GNAME19134(G19134,G59880,G15231);
  nand GNAME19135(G19135,G60000,G15232);
  nand GNAME19136(G19136,G15687,G15688,G15689,G15690);
  nand GNAME19137(G19137,G59992,G15187);
  nand GNAME19138(G19138,G59984,G15190);
  nand GNAME19139(G19139,G59976,G15191);
  nand GNAME19140(G19140,G59968,G15193);
  nand GNAME19141(G19141,G59960,G15195);
  nand GNAME19142(G19142,G59952,G15196);
  nand GNAME19143(G19143,G59944,G15197);
  nand GNAME19144(G19144,G59936,G15199);
  nand GNAME19145(G19145,G59928,G15200);
  nand GNAME19146(G19146,G59920,G15202);
  nand GNAME19147(G19147,G59912,G15203);
  nand GNAME19148(G19148,G59904,G15204);
  nand GNAME19149(G19149,G59896,G15205);
  nand GNAME19150(G19150,G59888,G15206);
  nand GNAME19151(G19151,G59880,G15207);
  nand GNAME19152(G19152,G60000,G15208);
  nand GNAME19153(G19153,G15683,G15684,G15685,G15686);
  nand GNAME19154(G19154,G15181,G23419);
  nand GNAME19155(G19155,G19153,G14821);
  nand GNAME19156(G19156,G19136,G15233);
  nand GNAME19157(G19157,G19119,G15234);
  nand GNAME19158(G19158,G59993,G15211);
  nand GNAME19159(G19159,G59985,G15213);
  nand GNAME19160(G19160,G59977,G15215);
  nand GNAME19161(G19161,G59969,G15218);
  nand GNAME19162(G19162,G59961,G15219);
  nand GNAME19163(G19163,G59953,G15220);
  nand GNAME19164(G19164,G59945,G15221);
  nand GNAME19165(G19165,G59937,G15223);
  nand GNAME19166(G19166,G59929,G15224);
  nand GNAME19167(G19167,G59921,G15225);
  nand GNAME19168(G19168,G59913,G15226);
  nand GNAME19169(G19169,G59905,G15228);
  nand GNAME19170(G19170,G59897,G15229);
  nand GNAME19171(G19171,G59889,G15230);
  nand GNAME19172(G19172,G59881,G15231);
  nand GNAME19173(G19173,G60001,G15232);
  nand GNAME19174(G19174,G15703,G15704,G15705,G15706);
  nand GNAME19175(G19175,G59993,G15187);
  nand GNAME19176(G19176,G59985,G15190);
  nand GNAME19177(G19177,G59977,G15191);
  nand GNAME19178(G19178,G59969,G15193);
  nand GNAME19179(G19179,G59961,G15195);
  nand GNAME19180(G19180,G59953,G15196);
  nand GNAME19181(G19181,G59945,G15197);
  nand GNAME19182(G19182,G59937,G15199);
  nand GNAME19183(G19183,G59929,G15200);
  nand GNAME19184(G19184,G59921,G15202);
  nand GNAME19185(G19185,G59913,G15203);
  nand GNAME19186(G19186,G59905,G15204);
  nand GNAME19187(G19187,G59897,G15205);
  nand GNAME19188(G19188,G59889,G15206);
  nand GNAME19189(G19189,G59881,G15207);
  nand GNAME19190(G19190,G60001,G15208);
  nand GNAME19191(G19191,G15699,G15700,G15701,G15702);
  nand GNAME19192(G19192,G59993,G17265);
  nand GNAME19193(G19193,G59985,G17326);
  nand GNAME19194(G19194,G59977,G17387);
  nand GNAME19195(G19195,G59969,G17448);
  nand GNAME19196(G19196,G59961,G17509);
  nand GNAME19197(G19197,G59953,G17570);
  nand GNAME19198(G19198,G59945,G17631);
  nand GNAME19199(G19199,G59937,G17692);
  nand GNAME19200(G19200,G59929,G17753);
  nand GNAME19201(G19201,G59921,G17814);
  nand GNAME19202(G19202,G59913,G17875);
  nand GNAME19203(G19203,G59905,G17936);
  nand GNAME19204(G19204,G59897,G17997);
  nand GNAME19205(G19205,G59889,G18058);
  nand GNAME19206(G19206,G59881,G18119);
  nand GNAME19207(G19207,G60001,G17183);
  nand GNAME19208(G19208,G15695,G15696,G15697,G15698);
  or GNAME19209(G19209,G15880,G19979);
  nand GNAME19210(G19210,G15181,G23423);
  nand GNAME19211(G19211,G19208,G15234);
  nand GNAME19212(G19212,G19191,G14821);
  nand GNAME19213(G19213,G19174,G15233);
  nand GNAME19214(G19214,G59994,G15211);
  nand GNAME19215(G19215,G59986,G15213);
  nand GNAME19216(G19216,G59978,G15215);
  nand GNAME19217(G19217,G59970,G15218);
  nand GNAME19218(G19218,G59962,G15219);
  nand GNAME19219(G19219,G59954,G15220);
  nand GNAME19220(G19220,G59946,G15221);
  nand GNAME19221(G19221,G59938,G15223);
  nand GNAME19222(G19222,G59930,G15224);
  nand GNAME19223(G19223,G59922,G15225);
  nand GNAME19224(G19224,G59914,G15226);
  nand GNAME19225(G19225,G59906,G15228);
  nand GNAME19226(G19226,G59898,G15229);
  nand GNAME19227(G19227,G59890,G15230);
  nand GNAME19228(G19228,G59882,G15231);
  nand GNAME19229(G19229,G60002,G15232);
  nand GNAME19230(G19230,G15715,G15716,G15717,G15718);
  nand GNAME19231(G19231,G59994,G15187);
  nand GNAME19232(G19232,G59986,G15190);
  nand GNAME19233(G19233,G59978,G15191);
  nand GNAME19234(G19234,G59970,G15193);
  nand GNAME19235(G19235,G59962,G15195);
  nand GNAME19236(G19236,G59954,G15196);
  nand GNAME19237(G19237,G59946,G15197);
  nand GNAME19238(G19238,G59938,G15199);
  nand GNAME19239(G19239,G59930,G15200);
  nand GNAME19240(G19240,G59922,G15202);
  nand GNAME19241(G19241,G59914,G15203);
  nand GNAME19242(G19242,G59906,G15204);
  nand GNAME19243(G19243,G59898,G15205);
  nand GNAME19244(G19244,G59890,G15206);
  nand GNAME19245(G19245,G59882,G15207);
  nand GNAME19246(G19246,G60002,G15208);
  nand GNAME19247(G19247,G15711,G15712,G15713,G15714);
  nand GNAME19248(G19248,G59994,G17265);
  nand GNAME19249(G19249,G59986,G17326);
  nand GNAME19250(G19250,G59978,G17387);
  nand GNAME19251(G19251,G59970,G17448);
  nand GNAME19252(G19252,G59962,G17509);
  nand GNAME19253(G19253,G59954,G17570);
  nand GNAME19254(G19254,G59946,G17631);
  nand GNAME19255(G19255,G59938,G17692);
  nand GNAME19256(G19256,G59930,G17753);
  nand GNAME19257(G19257,G59922,G17814);
  nand GNAME19258(G19258,G59914,G17875);
  nand GNAME19259(G19259,G59906,G17936);
  nand GNAME19260(G19260,G59898,G17997);
  nand GNAME19261(G19261,G59890,G18058);
  nand GNAME19262(G19262,G59882,G18119);
  nand GNAME19263(G19263,G60002,G17183);
  nand GNAME19264(G19264,G15707,G15708,G15709,G15710);
  nand GNAME19265(G19265,G15181,G23421);
  nand GNAME19266(G19266,G19264,G15234);
  nand GNAME19267(G19267,G19247,G14821);
  nand GNAME19268(G19268,G19230,G15233);
  nand GNAME19269(G19269,G14778,G60007);
  nand GNAME19270(G19270,G60003,G15232);
  nand GNAME19271(G19271,G59995,G15211);
  nand GNAME19272(G19272,G59987,G15213);
  nand GNAME19273(G19273,G59979,G15215);
  nand GNAME19274(G19274,G59971,G15218);
  nand GNAME19275(G19275,G59963,G15219);
  nand GNAME19276(G19276,G59955,G15220);
  nand GNAME19277(G19277,G59947,G15221);
  nand GNAME19278(G19278,G59939,G15223);
  nand GNAME19279(G19279,G59931,G15224);
  nand GNAME19280(G19280,G59923,G15225);
  nand GNAME19281(G19281,G59915,G15226);
  nand GNAME19282(G19282,G59907,G15228);
  nand GNAME19283(G19283,G59899,G15229);
  nand GNAME19284(G19284,G59891,G15230);
  nand GNAME19285(G19285,G59883,G15231);
  nand GNAME19286(G19286,G15727,G15728,G15729,G15730);
  nand GNAME19287(G19287,G60003,G15208);
  nand GNAME19288(G19288,G59995,G15187);
  nand GNAME19289(G19289,G59987,G15190);
  nand GNAME19290(G19290,G59979,G15191);
  nand GNAME19291(G19291,G59971,G15193);
  nand GNAME19292(G19292,G59963,G15195);
  nand GNAME19293(G19293,G59955,G15196);
  nand GNAME19294(G19294,G59947,G15197);
  nand GNAME19295(G19295,G59939,G15199);
  nand GNAME19296(G19296,G59931,G15200);
  nand GNAME19297(G19297,G59923,G15202);
  nand GNAME19298(G19298,G59915,G15203);
  nand GNAME19299(G19299,G59907,G15204);
  nand GNAME19300(G19300,G59899,G15205);
  nand GNAME19301(G19301,G59891,G15206);
  nand GNAME19302(G19302,G59883,G15207);
  nand GNAME19303(G19303,G15723,G15724,G15725,G15726);
  nand GNAME19304(G19304,G60003,G17183);
  nand GNAME19305(G19305,G59995,G17265);
  nand GNAME19306(G19306,G59987,G17326);
  nand GNAME19307(G19307,G59979,G17387);
  nand GNAME19308(G19308,G59971,G17448);
  nand GNAME19309(G19309,G59963,G17509);
  nand GNAME19310(G19310,G59955,G17570);
  nand GNAME19311(G19311,G59947,G17631);
  nand GNAME19312(G19312,G59939,G17692);
  nand GNAME19313(G19313,G59931,G17753);
  nand GNAME19314(G19314,G59923,G17814);
  nand GNAME19315(G19315,G59915,G17875);
  nand GNAME19316(G19316,G59907,G17936);
  nand GNAME19317(G19317,G59899,G17997);
  nand GNAME19318(G19318,G59891,G18058);
  nand GNAME19319(G19319,G59883,G18119);
  nand GNAME19320(G19320,G15719,G15720,G15721,G15722);
  nand GNAME19321(G19321,G15181,G23422);
  nand GNAME19322(G19322,G19320,G15234);
  nand GNAME19323(G19323,G19303,G14821);
  nand GNAME19324(G19324,G19286,G15233);
  nand GNAME19325(G19325,G14778,G60008);
  nand GNAME19326(G19326,G60004,G15232);
  nand GNAME19327(G19327,G59996,G15211);
  nand GNAME19328(G19328,G59988,G15213);
  nand GNAME19329(G19329,G59980,G15215);
  nand GNAME19330(G19330,G59972,G15218);
  nand GNAME19331(G19331,G59964,G15219);
  nand GNAME19332(G19332,G59956,G15220);
  nand GNAME19333(G19333,G59948,G15221);
  nand GNAME19334(G19334,G59940,G15223);
  nand GNAME19335(G19335,G59932,G15224);
  nand GNAME19336(G19336,G59924,G15225);
  nand GNAME19337(G19337,G59916,G15226);
  nand GNAME19338(G19338,G59908,G15228);
  nand GNAME19339(G19339,G59900,G15229);
  nand GNAME19340(G19340,G59892,G15230);
  nand GNAME19341(G19341,G59884,G15231);
  nand GNAME19342(G19342,G15740,G15741,G15742,G15743);
  nand GNAME19343(G19343,G60004,G15208);
  nand GNAME19344(G19344,G59996,G15187);
  nand GNAME19345(G19345,G59988,G15190);
  nand GNAME19346(G19346,G59980,G15191);
  nand GNAME19347(G19347,G59972,G15193);
  nand GNAME19348(G19348,G59964,G15195);
  nand GNAME19349(G19349,G59956,G15196);
  nand GNAME19350(G19350,G59948,G15197);
  nand GNAME19351(G19351,G59940,G15199);
  nand GNAME19352(G19352,G59932,G15200);
  nand GNAME19353(G19353,G59924,G15202);
  nand GNAME19354(G19354,G59916,G15203);
  nand GNAME19355(G19355,G59908,G15204);
  nand GNAME19356(G19356,G59900,G15205);
  nand GNAME19357(G19357,G59892,G15206);
  nand GNAME19358(G19358,G59884,G15207);
  nand GNAME19359(G19359,G15736,G15737,G15738,G15739);
  nand GNAME19360(G19360,G60004,G17183);
  nand GNAME19361(G19361,G59996,G17265);
  nand GNAME19362(G19362,G59988,G17326);
  nand GNAME19363(G19363,G59980,G17387);
  nand GNAME19364(G19364,G59972,G17448);
  nand GNAME19365(G19365,G59964,G17509);
  nand GNAME19366(G19366,G59956,G17570);
  nand GNAME19367(G19367,G59948,G17631);
  nand GNAME19368(G19368,G59940,G17692);
  nand GNAME19369(G19369,G59932,G17753);
  nand GNAME19370(G19370,G59924,G17814);
  nand GNAME19371(G19371,G59916,G17875);
  nand GNAME19372(G19372,G59908,G17936);
  nand GNAME19373(G19373,G59900,G17997);
  nand GNAME19374(G19374,G59892,G18058);
  nand GNAME19375(G19375,G59884,G18119);
  nand GNAME19376(G19376,G15732,G15733,G15734,G15735);
  nand GNAME19377(G19377,G15181,G23417);
  nand GNAME19378(G19378,G19376,G15234);
  nand GNAME19379(G19379,G19359,G14821);
  nand GNAME19380(G19380,G19342,G15233);
  nand GNAME19381(G19381,G14778,G60009);
  nand GNAME19382(G19382,G60005,G15232);
  nand GNAME19383(G19383,G59997,G15211);
  nand GNAME19384(G19384,G59989,G15213);
  nand GNAME19385(G19385,G59981,G15215);
  nand GNAME19386(G19386,G59973,G15218);
  nand GNAME19387(G19387,G59965,G15219);
  nand GNAME19388(G19388,G59957,G15220);
  nand GNAME19389(G19389,G59949,G15221);
  nand GNAME19390(G19390,G59941,G15223);
  nand GNAME19391(G19391,G59933,G15224);
  nand GNAME19392(G19392,G59925,G15225);
  nand GNAME19393(G19393,G59917,G15226);
  nand GNAME19394(G19394,G59909,G15228);
  nand GNAME19395(G19395,G59901,G15229);
  nand GNAME19396(G19396,G59893,G15230);
  nand GNAME19397(G19397,G59885,G15231);
  nand GNAME19398(G19398,G15753,G15754,G15755,G15756);
  nand GNAME19399(G19399,G60005,G15208);
  nand GNAME19400(G19400,G59997,G15187);
  nand GNAME19401(G19401,G59989,G15190);
  nand GNAME19402(G19402,G59981,G15191);
  nand GNAME19403(G19403,G59973,G15193);
  nand GNAME19404(G19404,G59965,G15195);
  nand GNAME19405(G19405,G59957,G15196);
  nand GNAME19406(G19406,G59949,G15197);
  nand GNAME19407(G19407,G59941,G15199);
  nand GNAME19408(G19408,G59933,G15200);
  nand GNAME19409(G19409,G59925,G15202);
  nand GNAME19410(G19410,G59917,G15203);
  nand GNAME19411(G19411,G59909,G15204);
  nand GNAME19412(G19412,G59901,G15205);
  nand GNAME19413(G19413,G59893,G15206);
  nand GNAME19414(G19414,G59885,G15207);
  nand GNAME19415(G19415,G15749,G15750,G15751,G15752);
  nand GNAME19416(G19416,G60005,G17183);
  nand GNAME19417(G19417,G59997,G17265);
  nand GNAME19418(G19418,G59989,G17326);
  nand GNAME19419(G19419,G59981,G17387);
  nand GNAME19420(G19420,G59973,G17448);
  nand GNAME19421(G19421,G59965,G17509);
  nand GNAME19422(G19422,G59957,G17570);
  nand GNAME19423(G19423,G59949,G17631);
  nand GNAME19424(G19424,G59941,G17692);
  nand GNAME19425(G19425,G59933,G17753);
  nand GNAME19426(G19426,G59925,G17814);
  nand GNAME19427(G19427,G59917,G17875);
  nand GNAME19428(G19428,G59909,G17936);
  nand GNAME19429(G19429,G59901,G17997);
  nand GNAME19430(G19430,G59893,G18058);
  nand GNAME19431(G19431,G59885,G18119);
  nand GNAME19432(G19432,G15745,G15746,G15747,G15748);
  nand GNAME19433(G19433,G15181,G23420);
  nand GNAME19434(G19434,G19432,G15234);
  nand GNAME19435(G19435,G19415,G14821);
  nand GNAME19436(G19436,G19398,G15233);
  nand GNAME19437(G19437,G14778,G60010);
  nand GNAME19438(G19438,G14795,G15234,G59877,G14779,G15897);
  nand GNAME19439(G19439,G60003,G14853);
  or GNAME19440(G19440,G14784,G15914,G14747);
  nand GNAME19441(G19441,G14781,G59877,G14795,G19984);
  nand GNAME19442(G19442,G60004,G14853);
  nand GNAME19443(G19443,G14778,G15829);
  nand GNAME19444(G19444,G14788,G14884);
  nand GNAME19445(G19445,G15759,G19829,G19964,G14889,G15237);
  nand GNAME19446(G19446,G19445,G59877);
  nand GNAME19447(G19447,G60005,G14853);
  nand GNAME19448(G19448,G14849,G14857);
  nand GNAME19449(G19449,G15846,G14850);
  nand GNAME19450(G19450,G14777,G15948);
  nand GNAME19451(G19451,G19450,G19448,G19449);
  nand GNAME19452(G19452,G14743,G14789);
  nand GNAME19453(G19453,G14740,G14779);
  nand GNAME19454(G19454,G19453,G15780);
  nand GNAME19455(G19455,G19454,G14884);
  nand GNAME19456(G19456,G19452,G14824);
  nand GNAME19457(G19457,G14850,G14891);
  nand GNAME19458(G19458,G14789,G19451);
  nand GNAME19459(G19459,G14818,G14821);
  nand GNAME19460(G19460,G15760,G14892,G19458,G19459);
  nand GNAME19461(G19461,G19460,G59877);
  or GNAME19462(G19462,G14896,G14784);
  nand GNAME19463(G19463,G15804,G19438,G19462,G15238);
  nand GNAME19464(G19464,G15793,G15776);
  nand GNAME19465(G19465,G19464,G23199);
  nand GNAME19466(G19466,G19463,G60025);
  nand GNAME19467(G19467,G15777,G60057);
  nand GNAME19468(G19468,G14785,G60216);
  nand GNAME19469(G19469,G19464,G23156);
  nand GNAME19470(G19470,G19463,G60024);
  nand GNAME19471(G19471,G15777,G60056);
  nand GNAME19472(G19472,G14785,G60215);
  nand GNAME19473(G19473,G19464,G23157);
  nand GNAME19474(G19474,G19463,G60023);
  nand GNAME19475(G19475,G15777,G60055);
  nand GNAME19476(G19476,G14785,G60214);
  nand GNAME19477(G19477,G19464,G23123);
  nand GNAME19478(G19478,G19463,G60022);
  nand GNAME19479(G19479,G15777,G60054);
  nand GNAME19480(G19480,G14785,G60213);
  nand GNAME19481(G19481,G19464,G23158);
  nand GNAME19482(G19482,G19463,G60021);
  nand GNAME19483(G19483,G15777,G60053);
  nand GNAME19484(G19484,G14785,G60212);
  nand GNAME19485(G19485,G59877,G14868);
  nand GNAME19486(G19486,G19485,G14860);
  nand GNAME19487(G19487,G19486,G60006);
  nand GNAME19488(G19488,G19464,G23159);
  nand GNAME19489(G19489,G19463,G60020);
  nand GNAME19490(G19490,G15777,G60052);
  nand GNAME19491(G19491,G14785,G60211);
  nand GNAME19492(G19492,G19463,G60047);
  nand GNAME19493(G19493,G15777,G60079);
  nand GNAME19494(G19494,G14830,G23190);
  nand GNAME19495(G19495,G14785,G60238);
  nand GNAME19496(G19496,G19464,G23122);
  nand GNAME19497(G19497,G19463,G60046);
  nand GNAME19498(G19498,G15777,G60078);
  nand GNAME19499(G19499,G14785,G60237);
  nand GNAME19500(G19500,G18576,G14861);
  nand GNAME19501(G19501,G16827,G16828);
  nand GNAME19502(G19502,G19501,G59877);
  nand GNAME19503(G19503,G15180,G15235);
  or GNAME19504(G19504,G14899,G14784);
  nand GNAME19505(G19505,G19504,G15239,G19503,G15794,G16317);
  nand GNAME19506(G19506,G19505,G60007);
  nand GNAME19507(G19507,G19464,G23160);
  nand GNAME19508(G19508,G19463,G60019);
  nand GNAME19509(G19509,G15777,G60051);
  nand GNAME19510(G19510,G14785,G60210);
  nand GNAME19511(G19511,G19464,G23176);
  nand GNAME19512(G19512,G19463,G60045);
  nand GNAME19513(G19513,G15777,G60077);
  nand GNAME19514(G19514,G14785,G60236);
  nand GNAME19515(G19515,G18593,G14861);
  nand GNAME19516(G19516,G19464,G23177);
  nand GNAME19517(G19517,G19463,G60044);
  nand GNAME19518(G19518,G15777,G60076);
  nand GNAME19519(G19519,G14785,G60235);
  nand GNAME19520(G19520,G18610,G14861);
  nand GNAME19521(G19521,G19464,G23178);
  nand GNAME19522(G19522,G19463,G60043);
  nand GNAME19523(G19523,G15777,G60075);
  nand GNAME19524(G19524,G14785,G60234);
  nand GNAME19525(G19525,G18627,G14861);
  nand GNAME19526(G19526,G19464,G23179);
  nand GNAME19527(G19527,G19463,G60042);
  nand GNAME19528(G19528,G15777,G60074);
  nand GNAME19529(G19529,G14785,G60233);
  nand GNAME19530(G19530,G18644,G14861);
  nand GNAME19531(G19531,G19464,G23180);
  nand GNAME19532(G19532,G19463,G60041);
  nand GNAME19533(G19533,G15777,G60073);
  nand GNAME19534(G19534,G14785,G60232);
  nand GNAME19535(G19535,G18661,G14861);
  nand GNAME19536(G19536,G19464,G23181);
  nand GNAME19537(G19537,G19463,G60040);
  nand GNAME19538(G19538,G15777,G60072);
  nand GNAME19539(G19539,G14785,G60231);
  nand GNAME19540(G19540,G18678,G14861);
  nand GNAME19541(G19541,G19464,G23182);
  nand GNAME19542(G19542,G19463,G60039);
  nand GNAME19543(G19543,G15777,G60071);
  nand GNAME19544(G19544,G14785,G60230);
  nand GNAME19545(G19545,G18695,G14861);
  nand GNAME19546(G19546,G19464,G23183);
  nand GNAME19547(G19547,G19463,G60038);
  nand GNAME19548(G19548,G15777,G60070);
  nand GNAME19549(G19549,G14785,G60229);
  nand GNAME19550(G19550,G19464,G23184);
  nand GNAME19551(G19551,G19463,G60037);
  nand GNAME19552(G19552,G15777,G60069);
  nand GNAME19553(G19553,G14785,G60228);
  nand GNAME19554(G19554,G19464,G23185);
  nand GNAME19555(G19555,G19463,G60036);
  nand GNAME19556(G19556,G15777,G60068);
  nand GNAME19557(G19557,G14785,G60227);
  nand GNAME19558(G19558,G19505,G60008);
  nand GNAME19559(G19559,G19464,G23121);
  nand GNAME19560(G19560,G19463,G60018);
  nand GNAME19561(G19561,G15777,G60050);
  nand GNAME19562(G19562,G14785,G60209);
  nand GNAME19563(G19563,G19464,G23186);
  nand GNAME19564(G19564,G19463,G60035);
  nand GNAME19565(G19565,G15777,G60067);
  nand GNAME19566(G19566,G14785,G60226);
  nand GNAME19567(G19567,G19464,G23187);
  nand GNAME19568(G19568,G19463,G60034);
  nand GNAME19569(G19569,G15777,G60066);
  nand GNAME19570(G19570,G14785,G60225);
  nand GNAME19571(G19571,G19464,G23188);
  nand GNAME19572(G19572,G19463,G60033);
  nand GNAME19573(G19573,G15777,G60065);
  nand GNAME19574(G19574,G14785,G60224);
  nand GNAME19575(G19575,G19464,G23216);
  nand GNAME19576(G19576,G19463,G60032);
  nand GNAME19577(G19577,G15777,G60064);
  nand GNAME19578(G19578,G14785,G60223);
  nand GNAME19579(G19579,G19464,G23219);
  nand GNAME19580(G19580,G19463,G60031);
  nand GNAME19581(G19581,G15777,G60063);
  nand GNAME19582(G19582,G14785,G60222);
  nand GNAME19583(G19583,G19464,G23191);
  nand GNAME19584(G19584,G19463,G60030);
  nand GNAME19585(G19585,G15777,G60062);
  nand GNAME19586(G19586,G14785,G60221);
  nand GNAME19587(G19587,G19464,G23223);
  nand GNAME19588(G19588,G19463,G60029);
  nand GNAME19589(G19589,G15777,G60061);
  nand GNAME19590(G19590,G14785,G60220);
  nand GNAME19591(G19591,G19464,G23226);
  nand GNAME19592(G19592,G19463,G60028);
  nand GNAME19593(G19593,G15777,G60060);
  nand GNAME19594(G19594,G14785,G60219);
  nand GNAME19595(G19595,G19464,G23192);
  nand GNAME19596(G19596,G19463,G60027);
  nand GNAME19597(G19597,G15777,G60059);
  nand GNAME19598(G19598,G14785,G60218);
  nand GNAME19599(G19599,G19464,G23120);
  nand GNAME19600(G19600,G19463,G60026);
  nand GNAME19601(G19601,G15777,G60058);
  nand GNAME19602(G19602,G14785,G60217);
  nand GNAME19603(G19603,G19505,G60009);
  nand GNAME19604(G19604,G19464,G23213);
  nand GNAME19605(G19605,G19463,G60017);
  nand GNAME19606(G19606,G15777,G60049);
  nand GNAME19607(G19607,G14785,G60208);
  nand GNAME19608(G19608,G19505,G60010);
  nand GNAME19609(G19609,G19464,G23189);
  nand GNAME19610(G19610,G19463,G60016);
  nand GNAME19611(G19611,G15777,G60048);
  nand GNAME19612(G19612,G14785,G60207);
  nand GNAME19613(G19613,G14780,G19967,G19968);
  or GNAME19614(G19614,G15948,G14820);
  nand GNAME19615(G19615,G15880,G14788);
  nand GNAME19616(G19616,G15761,G15237,G19969,G19970);
  nand GNAME19617(G19617,G19616,G59877);
  nand GNAME19618(G19618,G14798,G15235);
  nand GNAME19619(G19619,G59877,G14893);
  nand GNAME19620(G19620,G15806,G19618,G19619,G15239);
  nand GNAME19621(G19621,G16218,G15950);
  nand GNAME19622(G19622,G19621,G60184);
  nand GNAME19623(G19623,G19620,G60025);
  nand GNAME19624(G19624,G60152,G15241);
  nand GNAME19625(G19625,G14830,G60057);
  nand GNAME19626(G19626,G14853,G13988);
  nand GNAME19627(G19627,G19621,G60183);
  nand GNAME19628(G19628,G19620,G60024);
  nand GNAME19629(G19629,G60151,G15241);
  nand GNAME19630(G19630,G14830,G60056);
  nand GNAME19631(G19631,G14853,G8114);
  nand GNAME19632(G19632,G19621,G60182);
  nand GNAME19633(G19633,G19620,G60023);
  nand GNAME19634(G19634,G60150,G15241);
  nand GNAME19635(G19635,G14830,G60055);
  nand GNAME19636(G19636,G14853,G8113);
  nand GNAME19637(G19637,G19621,G60181);
  nand GNAME19638(G19638,G19620,G60022);
  nand GNAME19639(G19639,G60149,G15241);
  nand GNAME19640(G19640,G14830,G60054);
  nand GNAME19641(G19641,G14853,G8112);
  nand GNAME19642(G19642,G19621,G60180);
  nand GNAME19643(G19643,G19620,G60021);
  nand GNAME19644(G19644,G60148,G15241);
  nand GNAME19645(G19645,G14830,G60053);
  nand GNAME19646(G19646,G14853,G8111);
  nand GNAME19647(G19647,G19621,G60179);
  nand GNAME19648(G19648,G19620,G60020);
  nand GNAME19649(G19649,G60147,G15241);
  nand GNAME19650(G19650,G14830,G60052);
  nand GNAME19651(G19651,G14853,G8110);
  nand GNAME19652(G19652,G19621,G60206);
  nand GNAME19653(G19653,G19620,G60047);
  nand GNAME19654(G19654,G60174,G15241);
  nand GNAME19655(G19655,G14830,G60079);
  nand GNAME19656(G19656,G19621,G60205);
  nand GNAME19657(G19657,G19620,G60046);
  nand GNAME19658(G19658,G60173,G15241);
  nand GNAME19659(G19659,G14830,G60078);
  nand GNAME19660(G19660,G14853,G8107);
  nand GNAME19661(G19661,G23088,G15235);
  nand GNAME19662(G19662,G15238,G15988,G19661);
  nand GNAME19663(G19663,G19662,G60007);
  nand GNAME19664(G19664,G19621,G60178);
  nand GNAME19665(G19665,G19620,G60019);
  nand GNAME19666(G19666,G60146,G15241);
  nand GNAME19667(G19667,G14830,G60051);
  nand GNAME19668(G19668,G14853,G8109);
  nand GNAME19669(G19669,G14810,G19876);
  nand GNAME19670(G19670,G14938,G14937);
  nand GNAME19671(G19671,G14799,G60012);
  nand GNAME19672(G19672,G19621,G60204);
  nand GNAME19673(G19673,G19620,G60045);
  nand GNAME19674(G19674,G60172,G15241);
  nand GNAME19675(G19675,G14830,G60077);
  nand GNAME19676(G19676,G14853,G14029);
  nand GNAME19677(G19677,G19621,G60203);
  nand GNAME19678(G19678,G19620,G60044);
  nand GNAME19679(G19679,G60171,G15241);
  nand GNAME19680(G19680,G14830,G60076);
  nand GNAME19681(G19681,G14853,G14030);
  nand GNAME19682(G19682,G19621,G60202);
  nand GNAME19683(G19683,G19620,G60043);
  nand GNAME19684(G19684,G60170,G15241);
  nand GNAME19685(G19685,G14830,G60075);
  nand GNAME19686(G19686,G14853,G8105);
  nand GNAME19687(G19687,G19621,G60201);
  nand GNAME19688(G19688,G19620,G60042);
  nand GNAME19689(G19689,G60169,G15241);
  nand GNAME19690(G19690,G14830,G60074);
  nand GNAME19691(G19691,G14853,G14031);
  nand GNAME19692(G19692,G19621,G60200);
  nand GNAME19693(G19693,G19620,G60041);
  nand GNAME19694(G19694,G60168,G15241);
  nand GNAME19695(G19695,G14830,G60073);
  nand GNAME19696(G19696,G14853,G14032);
  nand GNAME19697(G19697,G19621,G60199);
  nand GNAME19698(G19698,G19620,G60040);
  nand GNAME19699(G19699,G60167,G15241);
  nand GNAME19700(G19700,G14830,G60072);
  nand GNAME19701(G19701,G14853,G8081);
  nand GNAME19702(G19702,G19621,G60198);
  nand GNAME19703(G19703,G19620,G60039);
  nand GNAME19704(G19704,G60166,G15241);
  nand GNAME19705(G19705,G14830,G60071);
  nand GNAME19706(G19706,G14853,G8080);
  nand GNAME19707(G19707,G19621,G60197);
  nand GNAME19708(G19708,G19620,G60038);
  nand GNAME19709(G19709,G60165,G15241);
  nand GNAME19710(G19710,G14830,G60070);
  nand GNAME19711(G19711,G14853,G8079);
  nand GNAME19712(G19712,G19621,G60196);
  nand GNAME19713(G19713,G19620,G60037);
  nand GNAME19714(G19714,G60164,G15241);
  nand GNAME19715(G19715,G14830,G60069);
  nand GNAME19716(G19716,G14853,G8078);
  nand GNAME19717(G19717,G19621,G60195);
  nand GNAME19718(G19718,G19620,G60036);
  nand GNAME19719(G19719,G60163,G15241);
  nand GNAME19720(G19720,G14830,G60068);
  nand GNAME19721(G19721,G14853,G8077);
  nand GNAME19722(G19722,G19662,G60008);
  nand GNAME19723(G19723,G19621,G60177);
  nand GNAME19724(G19724,G19620,G60018);
  nand GNAME19725(G19725,G60145,G15241);
  nand GNAME19726(G19726,G14830,G60050);
  nand GNAME19727(G19727,G14853,G8106);
  nand GNAME19728(G19728,G19889,G14937);
  nand GNAME19729(G19729,G14810,G17063);
  nand GNAME19730(G19730,G14799,G60013);
  nand GNAME19731(G19731,G19621,G60194);
  nand GNAME19732(G19732,G19620,G60035);
  nand GNAME19733(G19733,G60162,G15241);
  nand GNAME19734(G19734,G14830,G60067);
  nand GNAME19735(G19735,G14853,G8075);
  nand GNAME19736(G19736,G19621,G60193);
  nand GNAME19737(G19737,G19620,G60034);
  nand GNAME19738(G19738,G60161,G15241);
  nand GNAME19739(G19739,G14830,G60066);
  nand GNAME19740(G19740,G14853,G8074);
  nand GNAME19741(G19741,G19621,G60192);
  nand GNAME19742(G19742,G19620,G60033);
  nand GNAME19743(G19743,G60160,G15241);
  nand GNAME19744(G19744,G14830,G60065);
  nand GNAME19745(G19745,G14853,G8073);
  nand GNAME19746(G19746,G19621,G60191);
  nand GNAME19747(G19747,G19620,G60032);
  nand GNAME19748(G19748,G60159,G15241);
  nand GNAME19749(G19749,G14830,G60064);
  nand GNAME19750(G19750,G14853,G8103);
  nand GNAME19751(G19751,G19621,G60190);
  nand GNAME19752(G19752,G19620,G60031);
  nand GNAME19753(G19753,G60158,G15241);
  nand GNAME19754(G19754,G14830,G60063);
  nand GNAME19755(G19755,G14853,G8102);
  nand GNAME19756(G19756,G19621,G60189);
  nand GNAME19757(G19757,G19620,G60030);
  nand GNAME19758(G19758,G60157,G15241);
  nand GNAME19759(G19759,G14830,G60062);
  nand GNAME19760(G19760,G14853,G8101);
  nand GNAME19761(G19761,G19621,G60188);
  nand GNAME19762(G19762,G19620,G60029);
  nand GNAME19763(G19763,G60156,G15241);
  nand GNAME19764(G19764,G14830,G60061);
  nand GNAME19765(G19765,G14853,G8100);
  nand GNAME19766(G19766,G19621,G60187);
  nand GNAME19767(G19767,G19620,G60028);
  nand GNAME19768(G19768,G60155,G15241);
  nand GNAME19769(G19769,G14830,G60060);
  nand GNAME19770(G19770,G14853,G8099);
  nand GNAME19771(G19771,G19621,G60186);
  nand GNAME19772(G19772,G19620,G60027);
  nand GNAME19773(G19773,G60154,G15241);
  nand GNAME19774(G19774,G14830,G60059);
  nand GNAME19775(G19775,G14853,G8098);
  nand GNAME19776(G19776,G19621,G60185);
  nand GNAME19777(G19777,G19620,G60026);
  nand GNAME19778(G19778,G60153,G15241);
  nand GNAME19779(G19779,G14830,G60058);
  nand GNAME19780(G19780,G14853,G8097);
  nand GNAME19781(G19781,G19662,G60009);
  nand GNAME19782(G19782,G19621,G60176);
  nand GNAME19783(G19783,G19620,G60017);
  nand GNAME19784(G19784,G60144,G15241);
  nand GNAME19785(G19785,G14830,G60049);
  nand GNAME19786(G19786,G14853,G8104);
  nand GNAME19787(G19787,G15247,G14810);
  nand GNAME19788(G19788,G19883,G14937);
  nand GNAME19789(G19789,G14799,G60014);
  nand GNAME19790(G19790,G19662,G60010);
  nand GNAME19791(G19791,G19621,G60175);
  nand GNAME19792(G19792,G19620,G60016);
  nand GNAME19793(G19793,G60143,G15241);
  nand GNAME19794(G19794,G14830,G60048);
  nand GNAME19795(G19795,G14853,G8096);
  nand GNAME19796(G19796,G17093,G14937);
  nand GNAME19797(G19797,G14810,G17041);
  nand GNAME19798(G19798,G14799,G60015);
  not GNAME19799(G19799,G15242);
  or GNAME19800(G19800,G14831,G19979);
  nand GNAME19801(G19801,G19208,G19799);
  nand GNAME19802(G19802,G19264,G19799);
  nand GNAME19803(G19803,G60007,G59874);
  nand GNAME19804(G19804,G14777,G15914);
  nand GNAME19805(G19805,G19804,G15787);
  nand GNAME19806(G19806,G19805,G15105);
  nand GNAME19807(G19807,G19320,G19799);
  nand GNAME19808(G19808,G60008,G59874);
  nand GNAME19809(G19809,G14777,G19971,G19972);
  nand GNAME19810(G19810,G19376,G19799);
  nand GNAME19811(G19811,G19432,G19799);
  nand GNAME19812(G19812,G15787,G15243);
  nand GNAME19813(G19813,G23784,G15244);
  nand GNAME19814(G19814,G59876,G14112);
  nand GNAME19815(G19815,G15244,G23798);
  nand GNAME19816(G19816,G59876,G14034);
  nand GNAME19817(G19817,G15244,G23799);
  nand GNAME19818(G19818,G59876,G14033);
  nand GNAME19819(G19819,G15244,G23800);
  nand GNAME19820(G19820,G59876,G14036);
  nand GNAME19821(G19821,G15244,G23797);
  nand GNAME19822(G19822,G59876,G14035);
  nand GNAME19823(G19823,G15244,G23785);
  nand GNAME19824(G19824,G14779,G15243);
  nand GNAME19825(G19825,G14831,G19824);
  nand GNAME19826(G19826,G59840,G18206,G18207);
  nand GNAME19827(G19827,G60247,G15107,G59841);
  nand GNAME19828(G19828,G59840,G1589,G18211);
  nand GNAME19829(G19829,G14779,G15180);
  nand GNAME19830(G19830,G19978,G60253);
  nand GNAME19831(G19831,G15766,G15955);
  nand GNAME19832(G19832,G60252,G19978);
  nand GNAME19833(G19833,G15766,G15956);
  nand GNAME19834(G19834,G15781,G60249);
  nand GNAME19835(G19835,G14808,G60253);
  or GNAME19836(G19836,G60250,G15781);
  nand GNAME19837(G19837,G15781,G60248);
  nand GNAME19838(G19838,G60247,G15767);
  or GNAME19839(G19839,G15767,G15984);
  nand GNAME19840(G19840,G14804,G35);
  nand GNAME19841(G19841,G15958,G60246);
  nand GNAME19842(G19842,G14778,G15846);
  nand GNAME19843(G19843,G14793,G15880);
  not GNAME19844(G19844,G15246);
  nand GNAME19845(G19845,G15781,G60243);
  or GNAME19846(G19846,G60252,G15781);
  nand GNAME19847(G19847,G19982,G60242);
  nand GNAME19848(G19848,G14826,G60207);
  nand GNAME19849(G19849,G14777,G14780,G14779);
  nand GNAME19850(G19850,G15829,G14780,G14743);
  nand GNAME19851(G19851,G14780,G14891);
  nand GNAME19852(G19852,G16838,G15897);
  nand GNAME19853(G19853,G14789,G16830,G15948);
  nand GNAME19854(G19854,G14742,G15863);
  nand GNAME19855(G19855,G14811,G14810);
  nand GNAME19856(G19856,G59876,G14748,G14784);
  nand GNAME19857(G19857,G14914,G59877,G23088);
  nand GNAME19858(G19858,G60015,G17037);
  nand GNAME19859(G19859,G14835,G60016);
  nand GNAME19860(G19860,G15279,G60016);
  nand GNAME19861(G19861,G19859,G19860);
  or GNAME19862(G19862,G60015,G59875);
  nand GNAME19863(G19863,G14810,G60015);
  or GNAME19864(G19864,G15279,G60017);
  or GNAME19865(G19865,G14835,G2084);
  nand GNAME19866(G19866,G14917,G15798);
  nand GNAME19867(G19867,G14916,G17048);
  nand GNAME19868(G19868,G17052,G15396);
  or GNAME19869(G19869,G17052,G15396);
  not GNAME19870(G19870,G15247);
  or GNAME19871(G19871,G14920,G14919);
  nand GNAME19872(G19872,G14919,G14920);
  not GNAME19873(G19873,G15248);
  or GNAME19874(G19874,G15770,G15769);
  nand GNAME19875(G19875,G15769,G15770);
  not GNAME19876(G19876,G15249);
  or GNAME19877(G19877,G14749,G15771);
  nand GNAME19878(G19878,G15771,G17113);
  or GNAME19879(G19879,G17091,G15772);
  nand GNAME19880(G19880,G15772,G17091);
  nand GNAME19881(G19881,G17116,G15397);
  or GNAME19882(G19882,G17116,G15397);
  not GNAME19883(G19883,G15250);
  or GNAME19884(G19884,G14753,G15771);
  nand GNAME19885(G19885,G15771,G17131);
  nand GNAME19886(G19886,G17157,G17160);
  nand GNAME19887(G19887,G14933,G19886);
  nand GNAME19888(G19888,G17135,G17157,G17160);
  not GNAME19889(G19889,G15261);
  nand GNAME19890(G19890,G14789,G60008);
  nand GNAME19891(G19891,G14758,G15863);
  not GNAME19892(G19892,G15252);
  nand GNAME19893(G19893,G17141,G60008);
  nand GNAME19894(G19894,G14758,G15773);
  not GNAME19895(G19895,G15251);
  or GNAME19896(G19896,G14758,G15771);
  nand GNAME19897(G19897,G15771,G17152);
  or GNAME19898(G19898,G14765,G15774);
  nand GNAME19899(G19899,G15774,G17167);
  or GNAME19900(G19900,G14765,G15771);
  nand GNAME19901(G19901,G15771,G17179);
  nand GNAME19902(G19902,G15771,G14859,G14787,G23503);
  or GNAME19903(G19903,G19979,G15771);
  nand GNAME19904(G19904,G18184,G59877);
  nand GNAME19905(G19905,G14784,G18185);
  or GNAME19906(G19906,G14784,G15104);
  nand GNAME19907(G19907,G15104,G18191);
  nand GNAME19908(G19908,G15958,G59843);
  nand GNAME19909(G19909,G14804,G18201);
  nand GNAME19910(G19910,G14804,G15768,G18200);
  nand GNAME19911(G19911,G15958,G59842);
  nand GNAME19912(G19912,G14801,G18204);
  nand GNAME19913(G19913,G59840,G18202,G59841);
  or GNAME19914(G19914,G14803,G14745,G59840,G60247);
  nand GNAME19915(G19915,G14803,G15106,G59839);
  nand GNAME19916(G19916,G15781,G59808);
  nand GNAME19917(G19917,G14808,G60242);
  nand GNAME19918(G19918,G15781,G59807);
  nand GNAME19919(G19919,G14808,G60241);
  nand GNAME19920(G19920,G15781,G59806);
  nand GNAME19921(G19921,G14808,G60240);
  nand GNAME19922(G19922,G15781,G59805);
  nand GNAME19923(G19923,G14808,G60239);
  nand GNAME19924(G19924,G14758,G60009);
  nand GNAME19925(G19925,G14753,G60008);
  not GNAME19926(G19926,G15253);
  nand GNAME19927(G19927,G14753,G60007);
  nand GNAME19928(G19928,G60009,G14759);
  or GNAME19929(G19929,G60244,G14758);
  nand GNAME19930(G19930,G60244,G19861,G17063);
  or GNAME19931(G19931,G60244,G14753);
  nand GNAME19932(G19932,G60244,G19861,G15247);
  or GNAME19933(G19933,G60244,G14749);
  nand GNAME19934(G19934,G17109,G60244);
  nand GNAME19935(G19935,G15775,G23503,G14859);
  or GNAME19936(G19936,G19979,G15775);
  or GNAME19937(G19937,G14765,G15775);
  nand GNAME19938(G19938,G15775,G17176);
  or GNAME19939(G19939,G14758,G15775);
  nand GNAME19940(G19940,G15775,G17148);
  or GNAME19941(G19941,G14753,G15775);
  nand GNAME19942(G19942,G15775,G17127);
  or GNAME19943(G19943,G14749,G15775);
  nand GNAME19944(G19944,G15775,G17108);
  nand GNAME19945(G19945,G14811,G60206);
  nand GNAME19946(G19946,G59876,G60047);
  nand GNAME19947(G19947,G15863,G60046);
  nand GNAME19948(G19948,G14789,G18712);
  nand GNAME19949(G19949,G15863,G60045);
  nand GNAME19950(G19950,G14789,G18729);
  nand GNAME19951(G19951,G15863,G60044);
  nand GNAME19952(G19952,G14789,G18746);
  nand GNAME19953(G19953,G15863,G60043);
  nand GNAME19954(G19954,G14789,G18763);
  nand GNAME19955(G19955,G15863,G60042);
  nand GNAME19956(G19956,G14789,G18780);
  nand GNAME19957(G19957,G15863,G60041);
  nand GNAME19958(G19958,G14789,G18797);
  nand GNAME19959(G19959,G15863,G60040);
  nand GNAME19960(G19960,G14789,G18814);
  nand GNAME19961(G19961,G15863,G60039);
  nand GNAME19962(G19962,G14789,G18831);
  nand GNAME19963(G19963,G15948,G15914);
  nand GNAME19964(G19964,G14743,G14857);
  nand GNAME19965(G19965,G14789,G15948);
  nand GNAME19966(G19966,G14781,G15863);
  nand GNAME19967(G19967,G14779,G15829);
  nand GNAME19968(G19968,G14777,G14743);
  nand GNAME19969(G19969,G14793,G14884);
  nand GNAME19970(G19970,G15846,G15931);
  nand GNAME19971(G19971,G14779,G15846);
  nand GNAME19972(G19972,G14793,G15948);
  nand GNAME19973(G19973,G60009,G59874);
  nand GNAME19974(G19974,G14831,G19809);
  nand GNAME19975(G19975,G60010,G59874);
  nand GNAME19976(G19976,G14831,G19805);
  not GNAME19977(G19977,G14800);
  not GNAME19978(G19978,G15766);
  not GNAME19979(G19979,G60006);
  not GNAME19980(G19980,G14941);
  not GNAME19981(G19981,G14905);
  not GNAME19982(G19982,G14826);
  not GNAME19983(G19983,G14791);
  not GNAME19984(G19984,G15182);
  nand GNAME19985(G19985,G19986,G23484);
  nand GNAME19986(G19986,G20058,G20059);
  or GNAME19987(G19987,G20061,G20060);
  nand GNAME19988(G19988,G19989,G23424);
  nand GNAME19989(G19989,G20060,G20061);
  nand GNAME19990(G19990,G23461,G14128);
  nand GNAME19991(G19991,G19992,G20062);
  or GNAME19992(G19992,G23461,G14128);
  nand GNAME19993(G19993,G23481,G14122);
  not GNAME19994(G19994,G20037);
  not GNAME19995(G19995,G20003);
  and GNAME19996(G19996,G14042,G14041);
  and GNAME19997(G19997,G14046,G14045);
  and GNAME19998(G19998,G14050,G14049);
  and GNAME19999(G19999,G14054,G14053);
  and GNAME20000(G20000,G14058,G14057);
  not GNAME20001(G20001,G23425);
  and GNAME20002(G20002,G14062,G14061);
  nor GNAME20003(G20003,G14040,G20031);
  and GNAME20004(G20004,G20049,G23541);
  and GNAME20005(G20005,G20045,G23529);
  and GNAME20006(G20006,G20041,G23520);
  and GNAME20007(G20007,G23479,G19994);
  nand GNAME20008(G20008,G20033,G23475);
  and GNAME20009(G20009,G14044,G14043);
  and GNAME20010(G20010,G14048,G14047);
  and GNAME20011(G20011,G14052,G14051);
  and GNAME20012(G20012,G14056,G14055);
  and GNAME20013(G20013,G14060,G14059);
  and GNAME20014(G20014,G14096,G14095);
  nand GNAME20015(G20015,G14064,G14063);
  nand GNAME20016(G20016,G14066,G14065);
  nand GNAME20017(G20017,G14068,G14067);
  nand GNAME20018(G20018,G14070,G14069);
  nand GNAME20019(G20019,G14072,G14071);
  nand GNAME20020(G20020,G14074,G14073);
  nand GNAME20021(G20021,G14076,G14075);
  nand GNAME20022(G20022,G14078,G14077);
  nand GNAME20023(G20023,G14080,G14079);
  nand GNAME20024(G20024,G14082,G14081);
  nand GNAME20025(G20025,G14084,G14083);
  nand GNAME20026(G20026,G14086,G14085);
  nand GNAME20027(G20027,G14088,G14087);
  nand GNAME20028(G20028,G14090,G14089);
  nand GNAME20029(G20029,G14092,G14091);
  nand GNAME20030(G20030,G14094,G14093);
  and GNAME20031(G20031,G14100,G20051);
  not GNAME20032(G20032,G23475);
  and GNAME20033(G20033,G20035,G23476);
  not GNAME20034(G20034,G23476);
  and GNAME20035(G20035,G23477,G14037);
  nand GNAME20036(G20036,G19994,G23478,G23479);
  nand GNAME20037(G20037,G23520,G20041,G23517);
  not GNAME20038(G20038,G23478);
  not GNAME20039(G20039,G23520);
  not GNAME20040(G20040,G23517);
  and GNAME20041(G20041,G23523,G14038);
  nand GNAME20042(G20042,G23529,G20045,G23526);
  not GNAME20043(G20043,G23529);
  not GNAME20044(G20044,G23526);
  and GNAME20045(G20045,G23535,G14039);
  nand GNAME20046(G20046,G23541,G20049,G23538);
  not GNAME20047(G20047,G23541);
  not GNAME20048(G20048,G23538);
  nor GNAME20049(G20049,G20003,G20050);
  not GNAME20050(G20050,G23480);
  and GNAME20051(G20051,G14102,G14101);
  and GNAME20052(G20052,G14106,G14105);
  not GNAME20053(G20053,G14123);
  not GNAME20054(G20054,G14124);
  and GNAME20055(G20055,G14109,G14108);
  not GNAME20056(G20056,G14125);
  and GNAME20057(G20057,G19985,G14111);
  not GNAME20058(G20058,G14126);
  and GNAME20059(G20059,G19988,G19987);
  not GNAME20060(G20060,G14127);
  and GNAME20061(G20061,G19991,G19990);
  and GNAME20062(G20062,G14129,G23496);
  not GNAME20063(G20063,G14128);
  not GNAME20064(G20064,G23496);
  and GNAME20065(G20065,G14098,G14097);
  not GNAME20066(G20066,G23896);
  not GNAME20067(G20067,G23988);
  not GNAME20068(G20068,G23980);
  nand GNAME20069(G20069,G23842,G24082);
  nand GNAME20070(G20070,G23960,G15181);
  nand GNAME20071(G20071,G20073,G20072);
  nand GNAME20072(G20072,G23842,G14264);
  nand GNAME20073(G20073,G23855,G15181);
  or GNAME20074(G20074,G23856,G23922);
  nand GNAME20075(G20075,G23856,G23922);
  nand GNAME20076(G20076,G23842,G14263);
  nand GNAME20077(G20077,G23857,G15181);
  or GNAME20078(G20078,G24006,G23921);
  nand GNAME20079(G20079,G24006,G23921);
  nand GNAME20080(G20080,G23842,G14262);
  nand GNAME20081(G20081,G20082,G59243);
  not GNAME20082(G20082,G59244);
  not GNAME20083(G20083,G59360);
  nand GNAME20084(G20084,G20085,G59692);
  not GNAME20085(G20085,G59693);
  and GNAME20086(G20086,G20095,G59809);
  or GNAME20087(G20087,G59816,G59831,G59819,G59821);
  nor GNAME20088(G20088,G59814,G59828,G59829,G59813,G20087);
  or GNAME20089(G20089,G59830,G59820,G59827,G59837);
  nor GNAME20090(G20090,G59838,G59822,G59815,G20089);
  or GNAME20091(G20091,G59832,G59810,G59834,G59824);
  nor GNAME20092(G20092,G59817,G59812,G59826,G20091);
  or GNAME20093(G20093,G59811,G59835,G59823,G59825);
  nor GNAME20094(G20094,G59818,G59836,G59833,G20093);
  nand GNAME20095(G20095,G20088,G20090,G20092,G20094);
  and GNAME20096(G20096,G20105,G59360);
  or GNAME20097(G20097,G59367,G59382,G59370,G59372);
  nor GNAME20098(G20098,G59365,G59379,G59380,G59364,G20097);
  or GNAME20099(G20099,G59381,G59371,G59378,G59388);
  nor GNAME20100(G20100,G59389,G59373,G59366,G20099);
  or GNAME20101(G20101,G59383,G59361,G59385,G59375);
  nor GNAME20102(G20102,G59368,G59363,G59377,G20101);
  or GNAME20103(G20103,G59362,G59386,G59374,G59376);
  nor GNAME20104(G20104,G59369,G59387,G59384,G20103);
  nand GNAME20105(G20105,G20098,G20100,G20102,G20104);
  nand GNAME20106(G20106,G20107,G60141);
  not GNAME20107(G20107,G60142);
  nand GNAME20108(G20108,G20135,G20138,G20139);
  not GNAME20109(G20109,G2138);
  not GNAME20110(G20110,G2142);
  not GNAME20111(G20111,G2149);
  not GNAME20112(G20112,G2140);
  not GNAME20113(G20113,G2147);
  not GNAME20114(G20114,G2137);
  not GNAME20115(G20115,G2143);
  nand GNAME20116(G20116,G20117,G20134);
  or GNAME20117(G20117,G2145,G20109);
  or GNAME20118(G20118,G2150,G20110);
  nand GNAME20119(G20119,G2151,G20115,G20118);
  or GNAME20120(G20120,G2141,G20111);
  nand GNAME20121(G20121,G20110,G2150);
  nand GNAME20122(G20122,G20121,G20119,G20120);
  or GNAME20123(G20123,G2148,G20112);
  nand GNAME20124(G20124,G20111,G2141);
  nand GNAME20125(G20125,G20124,G20122,G20123);
  or GNAME20126(G20126,G2139,G20113);
  nand GNAME20127(G20127,G20112,G2148);
  nand GNAME20128(G20128,G20127,G20125,G20126);
  or GNAME20129(G20129,G2146,G20109);
  nand GNAME20130(G20130,G20113,G2139);
  nand GNAME20131(G20131,G20130,G20128,G20129);
  or GNAME20132(G20132,G2146,G2145);
  nand GNAME20133(G20133,G20109,G20132);
  nand GNAME20134(G20134,G20133,G20131);
  nand GNAME20135(G20135,G20116,G20136,G20137);
  nand GNAME20136(G20136,G20114,G2144);
  or GNAME20137(G20137,G2144,G20114);
  nand GNAME20138(G20138,G20114,G2144,G2136);
  or GNAME20139(G20139,G20114,G2144,G2136);
  and GNAME20140(G20140,G20305,G20306);
  and GNAME20141(G20141,G20264,G20302);
  and GNAME20142(G20142,G20254,G20300);
  and GNAME20143(G20143,G20266,G20273);
  not GNAME20144(G20144,G2791);
  not GNAME20145(G20145,G2192);
  not GNAME20146(G20146,G2193);
  nor GNAME20147(G20147,G20263,G20175);
  nor GNAME20148(G20148,G20174,G20264);
  nor GNAME20149(G20149,G20173,G20249);
  nor GNAME20150(G20150,G20265,G20171,G20172);
  nor GNAME20151(G20151,G20170,G20266);
  not GNAME20152(G20152,G2191);
  not GNAME20153(G20153,G2190);
  not GNAME20154(G20154,G2189);
  not GNAME20155(G20155,G2188);
  not GNAME20156(G20156,G2187);
  not GNAME20157(G20157,G2186);
  not GNAME20158(G20158,G2185);
  not GNAME20159(G20159,G2184);
  nor GNAME20160(G20160,G20235,G20195);
  nor GNAME20161(G20161,G20422,G20193,G20194);
  nor GNAME20162(G20162,G20192,G20250);
  nor GNAME20163(G20163,G20297,G20190,G20191);
  nor GNAME20164(G20164,G20189,G20251);
  nor GNAME20165(G20165,G20298,G20187,G20188);
  nor GNAME20166(G20166,G20186,G20252);
  nor GNAME20167(G20167,G20299,G20184,G20185);
  or GNAME20168(G20168,G20253,G20182,G20183);
  and GNAME20169(G20169,G20284,G20256);
  and GNAME20170(G20170,G20312,G20313);
  and GNAME20171(G20171,G20326,G20327);
  and GNAME20172(G20172,G20328,G20329);
  and GNAME20173(G20173,G20314,G20315);
  and GNAME20174(G20174,G20316,G20317);
  and GNAME20175(G20175,G20324,G20325);
  nand GNAME20176(G20176,G20336,G20337);
  nand GNAME20177(G20177,G20338,G20339);
  nand GNAME20178(G20178,G20340,G20341);
  nand GNAME20179(G20179,G20342,G20343);
  nand GNAME20180(G20180,G20344,G20345);
  and GNAME20181(G20181,G20349,G20350);
  and GNAME20182(G20182,G20387,G20388);
  and GNAME20183(G20183,G20389,G20390);
  and GNAME20184(G20184,G20383,G20384);
  and GNAME20185(G20185,G20385,G20386);
  and GNAME20186(G20186,G20351,G20352);
  and GNAME20187(G20187,G20379,G20380);
  and GNAME20188(G20188,G20381,G20382);
  and GNAME20189(G20189,G20353,G20354);
  and GNAME20190(G20190,G20375,G20376);
  and GNAME20191(G20191,G20377,G20378);
  and GNAME20192(G20192,G20355,G20356);
  and GNAME20193(G20193,G20371,G20372);
  and GNAME20194(G20194,G20373,G20374);
  and GNAME20195(G20195,G20369,G20370);
  nand GNAME20196(G20196,G20393,G20394);
  nand GNAME20197(G20197,G20395,G20396);
  nand GNAME20198(G20198,G20397,G20398);
  nand GNAME20199(G20199,G20399,G20400);
  nand GNAME20200(G20200,G20401,G20402);
  nand GNAME20201(G20201,G20403,G20404);
  nand GNAME20202(G20202,G20405,G20406);
  nand GNAME20203(G20203,G20407,G20408);
  nand GNAME20204(G20204,G20409,G20410);
  nand GNAME20205(G20205,G20411,G20412);
  nand GNAME20206(G20206,G20415,G20416);
  nand GNAME20207(G20207,G20417,G20418);
  nand GNAME20208(G20208,G20419,G20420);
  nand GNAME20209(G20209,G20433,G20434);
  nand GNAME20210(G20210,G20391,G20392);
  nand GNAME20211(G20211,G20425,G20426);
  nand GNAME20212(G20212,G20431,G20432);
  not GNAME20213(G20213,G2175);
  not GNAME20214(G20214,G2182);
  not GNAME20215(G20215,G2183);
  not GNAME20216(G20216,G2174);
  nand GNAME20217(G20217,G20269,G20267);
  and GNAME20218(G20218,G20271,G20270);
  and GNAME20219(G20219,G20334,G20335);
  nand GNAME20220(G20220,G20268,G20267);
  not GNAME20221(G20221,G2152);
  not GNAME20222(G20222,G2172);
  not GNAME20223(G20223,G2171);
  not GNAME20224(G20224,G2170);
  not GNAME20225(G20225,G2168);
  nor GNAME20226(G20226,G20181,G20168);
  nor GNAME20227(G20227,G20183,G20253);
  nor GNAME20228(G20228,G20184,G20299);
  nor GNAME20229(G20229,G20187,G20298);
  nor GNAME20230(G20230,G20190,G20297);
  nand GNAME20231(G20231,G20261,G20259);
  and GNAME20232(G20232,G20262,G20258);
  and GNAME20233(G20233,G20413,G20414);
  nor GNAME20234(G20234,G20193,G20422);
  and GNAME20235(G20235,G20296,G20274);
  and GNAME20236(G20236,G20421,G20422);
  nand GNAME20237(G20237,G20294,G20257);
  and GNAME20238(G20238,G20295,G20274);
  and GNAME20239(G20239,G20423,G20424);
  and GNAME20240(G20240,G20292,G20278);
  nand GNAME20241(G20241,G20290,G20279);
  and GNAME20242(G20242,G20291,G20278);
  and GNAME20243(G20243,G20427,G20428);
  nand GNAME20244(G20244,G20288,G20280);
  and GNAME20245(G20245,G20289,G20279);
  and GNAME20246(G20246,G20429,G20430);
  nor GNAME20247(G20247,G20435,G20169);
  and GNAME20248(G20248,G20260,G20259);
  not GNAME20249(G20249,G20148);
  not GNAME20250(G20250,G20161);
  not GNAME20251(G20251,G20163);
  not GNAME20252(G20252,G20165);
  not GNAME20253(G20253,G20167);
  not GNAME20254(G20254,G20226);
  nand GNAME20255(G20255,G20276,G20158,G20275);
  nand GNAME20256(G20256,G20283,G20154,G20282);
  nand GNAME20257(G20257,G20277,G2185);
  nand GNAME20258(G20258,G20320,G2192);
  nand GNAME20259(G20259,G20323,G2193);
  nand GNAME20260(G20260,G20146,G20321,G20322);
  nand GNAME20261(G20261,G20260,G2791);
  nand GNAME20262(G20262,G20145,G20318,G20319);
  and GNAME20263(G20263,G20258,G20301);
  not GNAME20264(G20264,G20147);
  not GNAME20265(G20265,G20149);
  not GNAME20266(G20266,G20150);
  nand GNAME20267(G20267,G20330,G2191);
  nand GNAME20268(G20268,G20152,G20310,G20311);
  nand GNAME20269(G20269,G20268,G20151);
  nand GNAME20270(G20270,G20333,G2190);
  nand GNAME20271(G20271,G20153,G20331,G20332);
  or GNAME20272(G20272,G20171,G20265);
  nand GNAME20273(G20273,G20272,G20172);
  nand GNAME20274(G20274,G20368,G2184);
  or GNAME20275(G20275,G2169,G20144);
  nand GNAME20276(G20276,G20144,G2169);
  nand GNAME20277(G20277,G20276,G20275);
  nand GNAME20278(G20278,G20365,G2186);
  nand GNAME20279(G20279,G20362,G2187);
  nand GNAME20280(G20280,G20359,G2188);
  nand GNAME20281(G20281,G20155,G20357,G20358);
  or GNAME20282(G20282,G2173,G20144);
  nand GNAME20283(G20283,G20144,G2173);
  nand GNAME20284(G20284,G20270,G20304);
  nand GNAME20285(G20285,G20282,G20283);
  nand GNAME20286(G20286,G20285,G2189);
  not GNAME20287(G20287,G20247);
  nand GNAME20288(G20288,G20281,G20287);
  nand GNAME20289(G20289,G20156,G20360,G20361);
  nand GNAME20290(G20290,G20244,G20289);
  nand GNAME20291(G20291,G20157,G20363,G20364);
  nand GNAME20292(G20292,G20241,G20291);
  not GNAME20293(G20293,G20240);
  nand GNAME20294(G20294,G20255,G20293);
  nand GNAME20295(G20295,G20159,G20366,G20367);
  nand GNAME20296(G20296,G20237,G20295);
  not GNAME20297(G20297,G20162);
  not GNAME20298(G20298,G20164);
  not GNAME20299(G20299,G20166);
  nand GNAME20300(G20300,G20168,G20181);
  nand GNAME20301(G20301,G20231,G20262);
  nand GNAME20302(G20302,G20175,G20258,G20301);
  nand GNAME20303(G20303,G20256,G20286);
  nand GNAME20304(G20304,G20217,G20271);
  nand GNAME20305(G20305,G20304,G20270,G20303);
  nand GNAME20306(G20306,G20286,G20169);
  not GNAME20307(G20307,G20248);
  nand GNAME20308(G20308,G20255,G20257);
  nand GNAME20309(G20309,G20280,G20281);
  or GNAME20310(G20310,G2175,G20144);
  or GNAME20311(G20311,G2791,G20213);
  or GNAME20312(G20312,G2176,G20144);
  nand GNAME20313(G20313,G20144,G2176);
  or GNAME20314(G20314,G2179,G20144);
  nand GNAME20315(G20315,G20144,G2179);
  or GNAME20316(G20316,G2180,G20144);
  nand GNAME20317(G20317,G20144,G2180);
  or GNAME20318(G20318,G2182,G20144);
  or GNAME20319(G20319,G2791,G20214);
  nand GNAME20320(G20320,G20318,G20319);
  or GNAME20321(G20321,G2183,G20144);
  or GNAME20322(G20322,G2791,G20215);
  nand GNAME20323(G20323,G20321,G20322);
  or GNAME20324(G20324,G2181,G20144);
  nand GNAME20325(G20325,G20144,G2181);
  or GNAME20326(G20326,G2178,G20144);
  nand GNAME20327(G20327,G20144,G2178);
  or GNAME20328(G20328,G2177,G20144);
  nand GNAME20329(G20329,G20144,G2177);
  nand GNAME20330(G20330,G20310,G20311);
  or GNAME20331(G20331,G2174,G20144);
  or GNAME20332(G20332,G2791,G20216);
  nand GNAME20333(G20333,G20331,G20332);
  or GNAME20334(G20334,G20218,G20217);
  nand GNAME20335(G20335,G20217,G20218);
  nand GNAME20336(G20336,G20220,G20151);
  or GNAME20337(G20337,G20151,G20220);
  nand GNAME20338(G20338,G20150,G20170);
  or GNAME20339(G20339,G20150,G20170);
  nand GNAME20340(G20340,G20149,G20171);
  or GNAME20341(G20341,G20149,G20171);
  nand GNAME20342(G20342,G20148,G20173);
  or GNAME20343(G20343,G20148,G20173);
  nand GNAME20344(G20344,G20147,G20174);
  or GNAME20345(G20345,G20147,G20174);
  or GNAME20346(G20346,G2152,G20144);
  or GNAME20347(G20347,G2791,G20221);
  nand GNAME20348(G20348,G20346,G20347);
  or GNAME20349(G20349,G2153,G20144);
  nand GNAME20350(G20350,G20144,G2153);
  or GNAME20351(G20351,G2158,G20144);
  nand GNAME20352(G20352,G20144,G2158);
  or GNAME20353(G20353,G2161,G20144);
  nand GNAME20354(G20354,G20144,G2161);
  or GNAME20355(G20355,G2164,G20144);
  nand GNAME20356(G20356,G20144,G2164);
  or GNAME20357(G20357,G2172,G20144);
  or GNAME20358(G20358,G2791,G20222);
  nand GNAME20359(G20359,G20357,G20358);
  or GNAME20360(G20360,G2171,G20144);
  or GNAME20361(G20361,G2791,G20223);
  nand GNAME20362(G20362,G20360,G20361);
  or GNAME20363(G20363,G2170,G20144);
  or GNAME20364(G20364,G2791,G20224);
  nand GNAME20365(G20365,G20363,G20364);
  or GNAME20366(G20366,G2168,G20144);
  or GNAME20367(G20367,G2791,G20225);
  nand GNAME20368(G20368,G20366,G20367);
  or GNAME20369(G20369,G2167,G20144);
  nand GNAME20370(G20370,G20144,G2167);
  or GNAME20371(G20371,G2166,G20144);
  nand GNAME20372(G20372,G20144,G2166);
  or GNAME20373(G20373,G2165,G20144);
  nand GNAME20374(G20374,G20144,G2165);
  or GNAME20375(G20375,G2163,G20144);
  nand GNAME20376(G20376,G20144,G2163);
  or GNAME20377(G20377,G2162,G20144);
  nand GNAME20378(G20378,G20144,G2162);
  or GNAME20379(G20379,G2160,G20144);
  nand GNAME20380(G20380,G20144,G2160);
  or GNAME20381(G20381,G2159,G20144);
  nand GNAME20382(G20382,G20144,G2159);
  or GNAME20383(G20383,G2157,G20144);
  nand GNAME20384(G20384,G20144,G2157);
  or GNAME20385(G20385,G2156,G20144);
  nand GNAME20386(G20386,G20144,G2156);
  or GNAME20387(G20387,G2154,G20144);
  nand GNAME20388(G20388,G20144,G2154);
  or GNAME20389(G20389,G2155,G20144);
  nand GNAME20390(G20390,G20144,G2155);
  nand GNAME20391(G20391,G20254,G20348);
  nand GNAME20392(G20392,G20226,G20346,G20347);
  nand GNAME20393(G20393,G20182,G20227);
  or GNAME20394(G20394,G20227,G20182);
  nand GNAME20395(G20395,G20167,G20183);
  or GNAME20396(G20396,G20167,G20183);
  nand GNAME20397(G20397,G20185,G20228);
  or GNAME20398(G20398,G20228,G20185);
  nand GNAME20399(G20399,G20166,G20184);
  or GNAME20400(G20400,G20166,G20184);
  nand GNAME20401(G20401,G20165,G20186);
  or GNAME20402(G20402,G20165,G20186);
  nand GNAME20403(G20403,G20188,G20229);
  or GNAME20404(G20404,G20229,G20188);
  nand GNAME20405(G20405,G20164,G20187);
  or GNAME20406(G20406,G20164,G20187);
  nand GNAME20407(G20407,G20163,G20189);
  or GNAME20408(G20408,G20163,G20189);
  nand GNAME20409(G20409,G20191,G20230);
  or GNAME20410(G20410,G20230,G20191);
  nand GNAME20411(G20411,G20162,G20190);
  or GNAME20412(G20412,G20162,G20190);
  or GNAME20413(G20413,G20232,G20231);
  nand GNAME20414(G20414,G20231,G20232);
  nand GNAME20415(G20415,G20161,G20192);
  or GNAME20416(G20416,G20161,G20192);
  nand GNAME20417(G20417,G20194,G20234);
  or GNAME20418(G20418,G20234,G20194);
  nand GNAME20419(G20419,G20160,G20193);
  or GNAME20420(G20420,G20160,G20193);
  nand GNAME20421(G20421,G20195,G20235);
  or GNAME20422(G20422,G20235,G20195);
  or GNAME20423(G20423,G20238,G20237);
  nand GNAME20424(G20424,G20237,G20238);
  nand GNAME20425(G20425,G20293,G20308);
  nand GNAME20426(G20426,G20240,G20255,G20257);
  or GNAME20427(G20427,G20242,G20241);
  nand GNAME20428(G20428,G20241,G20242);
  or GNAME20429(G20429,G20245,G20244);
  nand GNAME20430(G20430,G20244,G20245);
  nand GNAME20431(G20431,G20287,G20309);
  nand GNAME20432(G20432,G20247,G20280,G20281);
  or GNAME20433(G20433,G20248,G20144);
  or GNAME20434(G20434,G2791,G20307);
  not GNAME20435(G20435,G20286);
  not GNAME20436(G20436,G2121);
  not GNAME20437(G20437,G2126);
  not GNAME20438(G20438,G2120);
  not GNAME20439(G20439,G2122);
  not GNAME20440(G20440,G2127);
  not GNAME20441(G20441,G2124);
  not GNAME20442(G20442,G2125);
  not GNAME20443(G20443,G2123);
  and GNAME20444(G20444,G20611,G20635);
  and GNAME20445(G20445,G20565,G20633);
  and GNAME20446(G20446,G20630,G20631);
  and GNAME20447(G20447,G20566,G20627);
  and GNAME20448(G20448,G20600,G20601);
  not GNAME20449(G20449,G2836);
  not GNAME20450(G20450,G2235);
  not GNAME20451(G20451,G2236);
  not GNAME20452(G20452,G2239);
  not GNAME20453(G20453,G2240);
  not GNAME20454(G20454,G2241);
  not GNAME20455(G20455,G2238);
  not GNAME20456(G20456,G2237);
  not GNAME20457(G20457,G2234);
  nor GNAME20458(G20458,G20515,G20480);
  and GNAME20459(G20459,G20593,G20567);
  nor GNAME20460(G20460,G20664,G20479,G20493);
  nor GNAME20461(G20461,G20492,G20611);
  nor GNAME20462(G20462,G20491,G20564);
  nor GNAME20463(G20463,G20569,G20489,G20490);
  nor GNAME20464(G20464,G20488,G20565);
  not GNAME20465(G20465,G2233);
  not GNAME20466(G20466,G2232);
  not GNAME20467(G20467,G2231);
  not GNAME20468(G20468,G2230);
  not GNAME20469(G20469,G2229);
  not GNAME20470(G20470,G2228);
  not GNAME20471(G20471,G2227);
  not GNAME20472(G20472,G2226);
  nor GNAME20473(G20473,G20536,G20494);
  nor GNAME20474(G20474,G20739,G20486,G20487);
  and GNAME20475(G20475,G20770,G20474);
  nor GNAME20476(G20476,G20484,G20771);
  nand GNAME20477(G20477,G20772,G20476);
  and GNAME20478(G20478,G20585,G20568);
  and GNAME20479(G20479,G20659,G20660);
  and GNAME20480(G20480,G20657,G20658);
  nand GNAME20481(G20481,G20661,G20662);
  and GNAME20482(G20482,G20676,G20677);
  and GNAME20483(G20483,G20678,G20679);
  and GNAME20484(G20484,G20680,G20681);
  and GNAME20485(G20485,G20682,G20683);
  and GNAME20486(G20486,G20722,G20723);
  and GNAME20487(G20487,G20724,G20725);
  and GNAME20488(G20488,G20686,G20687);
  and GNAME20489(G20489,G20694,G20695);
  and GNAME20490(G20490,G20696,G20697);
  and GNAME20491(G20491,G20688,G20689);
  and GNAME20492(G20492,G20690,G20691);
  and GNAME20493(G20493,G20692,G20693);
  and GNAME20494(G20494,G20720,G20721);
  nand GNAME20495(G20495,G20728,G20729);
  nand GNAME20496(G20496,G20730,G20731);
  nand GNAME20497(G20497,G20732,G20733);
  nand GNAME20498(G20498,G20734,G20735);
  nand GNAME20499(G20499,G20736,G20737);
  nand GNAME20500(G20500,G20756,G20757);
  nand GNAME20501(G20501,G20758,G20759);
  nand GNAME20502(G20502,G20760,G20761);
  nand GNAME20503(G20503,G20762,G20763);
  nand GNAME20504(G20504,G20764,G20765);
  nand GNAME20505(G20505,G20766,G20767);
  nand GNAME20506(G20506,G20665,G20666);
  nand GNAME20507(G20507,G20671,G20672);
  nand GNAME20508(G20508,G20726,G20727);
  not GNAME20509(G20509,G2218);
  not GNAME20510(G20510,G2220);
  not GNAME20511(G20511,G2222);
  not GNAME20512(G20512,G2224);
  not GNAME20513(G20513,G2225);
  not GNAME20514(G20514,G2221);
  and GNAME20515(G20515,G20597,G20570);
  and GNAME20516(G20516,G20663,G20664);
  nor GNAME20517(G20517,G20769,G20459);
  nand GNAME20518(G20518,G20591,G20575);
  and GNAME20519(G20519,G20592,G20572);
  and GNAME20520(G20520,G20667,G20668);
  nand GNAME20521(G20521,G20589,G20576);
  and GNAME20522(G20522,G20590,G20575);
  and GNAME20523(G20523,G20669,G20670);
  nor GNAME20524(G20524,G20768,G20478);
  not GNAME20525(G20525,G2194);
  not GNAME20526(G20526,G2209);
  not GNAME20527(G20527,G2208);
  not GNAME20528(G20528,G2207);
  not GNAME20529(G20529,G2206);
  not GNAME20530(G20530,G2205);
  not GNAME20531(G20531,G2204);
  not GNAME20532(G20532,G2203);
  not GNAME20533(G20533,G2202);
  nor GNAME20534(G20534,G20482,G20477);
  nor GNAME20535(G20535,G20487,G20739);
  and GNAME20536(G20536,G20626,G20602);
  and GNAME20537(G20537,G20738,G20739);
  nand GNAME20538(G20538,G20624,G20603);
  and GNAME20539(G20539,G20625,G20602);
  and GNAME20540(G20540,G20740,G20741);
  nand GNAME20541(G20541,G20622,G20604);
  and GNAME20542(G20542,G20623,G20603);
  and GNAME20543(G20543,G20742,G20743);
  nand GNAME20544(G20544,G20620,G20605);
  and GNAME20545(G20545,G20621,G20604);
  and GNAME20546(G20546,G20744,G20745);
  nand GNAME20547(G20547,G20618,G20606);
  and GNAME20548(G20548,G20619,G20605);
  and GNAME20549(G20549,G20746,G20747);
  nand GNAME20550(G20550,G20583,G20581);
  and GNAME20551(G20551,G20584,G20578);
  and GNAME20552(G20552,G20748,G20749);
  nand GNAME20553(G20553,G20616,G20607);
  and GNAME20554(G20554,G20617,G20606);
  and GNAME20555(G20555,G20750,G20751);
  nand GNAME20556(G20556,G20614,G20608);
  and GNAME20557(G20557,G20615,G20607);
  and GNAME20558(G20558,G20752,G20753);
  nand GNAME20559(G20559,G20612,G20609);
  and GNAME20560(G20560,G20613,G20608);
  and GNAME20561(G20561,G20754,G20755);
  nand GNAME20562(G20562,G20610,G20609);
  and GNAME20563(G20563,G20582,G20581);
  not GNAME20564(G20564,G20461);
  not GNAME20565(G20565,G20463);
  not GNAME20566(G20566,G20534);
  nand GNAME20567(G20567,G20574,G20450,G20573);
  nand GNAME20568(G20568,G20580,G20452,G20579);
  not GNAME20569(G20569,G20462);
  nand GNAME20570(G20570,G20656,G2234);
  nand GNAME20571(G20571,G20457,G20639,G20640);
  nand GNAME20572(G20572,G20643,G2236);
  or GNAME20573(G20573,G2219,G20449);
  nand GNAME20574(G20574,G20449,G2219);
  nand GNAME20575(G20575,G20655,G2237);
  nand GNAME20576(G20576,G20652,G2238);
  nand GNAME20577(G20577,G20455,G20644,G20645);
  nand GNAME20578(G20578,G20648,G2240);
  or GNAME20579(G20579,G2223,G20449);
  nand GNAME20580(G20580,G20449,G2223);
  nand GNAME20581(G20581,G20651,G2241);
  nand GNAME20582(G20582,G20454,G20649,G20650);
  nand GNAME20583(G20583,G20582,G2836);
  nand GNAME20584(G20584,G20453,G20646,G20647);
  nand GNAME20585(G20585,G20578,G20628);
  nand GNAME20586(G20586,G20579,G20580);
  nand GNAME20587(G20587,G20586,G2239);
  not GNAME20588(G20588,G20524);
  nand GNAME20589(G20589,G20577,G20588);
  nand GNAME20590(G20590,G20456,G20653,G20654);
  nand GNAME20591(G20591,G20521,G20590);
  nand GNAME20592(G20592,G20451,G20641,G20642);
  nand GNAME20593(G20593,G20572,G20598);
  nand GNAME20594(G20594,G20573,G20574);
  nand GNAME20595(G20595,G20594,G2235);
  not GNAME20596(G20596,G20517);
  nand GNAME20597(G20597,G20571,G20596);
  nand GNAME20598(G20598,G20518,G20592);
  nand GNAME20599(G20599,G20567,G20595);
  nand GNAME20600(G20600,G20599,G20572,G20598);
  nand GNAME20601(G20601,G20595,G20459);
  nand GNAME20602(G20602,G20719,G2226);
  nand GNAME20603(G20603,G20716,G2227);
  nand GNAME20604(G20604,G20713,G2228);
  nand GNAME20605(G20605,G20710,G2229);
  nand GNAME20606(G20606,G20707,G2230);
  nand GNAME20607(G20607,G20704,G2231);
  nand GNAME20608(G20608,G20701,G2232);
  nand GNAME20609(G20609,G20698,G2233);
  nand GNAME20610(G20610,G20465,G20684,G20685);
  not GNAME20611(G20611,G20460);
  nand GNAME20612(G20612,G20610,G20464);
  nand GNAME20613(G20613,G20466,G20699,G20700);
  nand GNAME20614(G20614,G20559,G20613);
  nand GNAME20615(G20615,G20467,G20702,G20703);
  nand GNAME20616(G20616,G20556,G20615);
  nand GNAME20617(G20617,G20468,G20705,G20706);
  nand GNAME20618(G20618,G20553,G20617);
  nand GNAME20619(G20619,G20469,G20708,G20709);
  nand GNAME20620(G20620,G20547,G20619);
  nand GNAME20621(G20621,G20470,G20711,G20712);
  nand GNAME20622(G20622,G20544,G20621);
  nand GNAME20623(G20623,G20471,G20714,G20715);
  nand GNAME20624(G20624,G20541,G20623);
  nand GNAME20625(G20625,G20472,G20717,G20718);
  nand GNAME20626(G20626,G20538,G20625);
  nand GNAME20627(G20627,G20477,G20482);
  nand GNAME20628(G20628,G20550,G20584);
  nand GNAME20629(G20629,G20568,G20587);
  nand GNAME20630(G20630,G20629,G20578,G20628);
  nand GNAME20631(G20631,G20587,G20478);
  or GNAME20632(G20632,G20489,G20569);
  nand GNAME20633(G20633,G20632,G20490);
  or GNAME20634(G20634,G20479,G20664);
  nand GNAME20635(G20635,G20634,G20493);
  not GNAME20636(G20636,G20563);
  nand GNAME20637(G20637,G20570,G20571);
  nand GNAME20638(G20638,G20576,G20577);
  or GNAME20639(G20639,G2218,G20449);
  or GNAME20640(G20640,G2836,G20509);
  or GNAME20641(G20641,G2220,G20449);
  or GNAME20642(G20642,G2836,G20510);
  nand GNAME20643(G20643,G20641,G20642);
  or GNAME20644(G20644,G2222,G20449);
  or GNAME20645(G20645,G2836,G20511);
  or GNAME20646(G20646,G2224,G20449);
  or GNAME20647(G20647,G2836,G20512);
  nand GNAME20648(G20648,G20646,G20647);
  or GNAME20649(G20649,G2225,G20449);
  or GNAME20650(G20650,G2836,G20513);
  nand GNAME20651(G20651,G20649,G20650);
  nand GNAME20652(G20652,G20644,G20645);
  or GNAME20653(G20653,G2221,G20449);
  or GNAME20654(G20654,G2836,G20514);
  nand GNAME20655(G20655,G20653,G20654);
  nand GNAME20656(G20656,G20639,G20640);
  or GNAME20657(G20657,G2217,G20449);
  nand GNAME20658(G20658,G20449,G2217);
  or GNAME20659(G20659,G2216,G20449);
  nand GNAME20660(G20660,G20449,G2216);
  nand GNAME20661(G20661,G20458,G20479);
  or GNAME20662(G20662,G20458,G20479);
  nand GNAME20663(G20663,G20480,G20515);
  or GNAME20664(G20664,G20515,G20480);
  nand GNAME20665(G20665,G20596,G20637);
  nand GNAME20666(G20666,G20517,G20570,G20571);
  or GNAME20667(G20667,G20519,G20518);
  nand GNAME20668(G20668,G20518,G20519);
  or GNAME20669(G20669,G20522,G20521);
  nand GNAME20670(G20670,G20521,G20522);
  nand GNAME20671(G20671,G20588,G20638);
  nand GNAME20672(G20672,G20524,G20576,G20577);
  or GNAME20673(G20673,G2194,G20449);
  or GNAME20674(G20674,G2836,G20525);
  nand GNAME20675(G20675,G20673,G20674);
  or GNAME20676(G20676,G2195,G20449);
  nand GNAME20677(G20677,G20449,G2195);
  or GNAME20678(G20678,G2196,G20449);
  nand GNAME20679(G20679,G20449,G2196);
  or GNAME20680(G20680,G2197,G20449);
  nand GNAME20681(G20681,G20449,G2197);
  or GNAME20682(G20682,G2198,G20449);
  nand GNAME20683(G20683,G20449,G2198);
  or GNAME20684(G20684,G2209,G20449);
  or GNAME20685(G20685,G2836,G20526);
  or GNAME20686(G20686,G2210,G20449);
  nand GNAME20687(G20687,G20449,G2210);
  or GNAME20688(G20688,G2213,G20449);
  nand GNAME20689(G20689,G20449,G2213);
  or GNAME20690(G20690,G2214,G20449);
  nand GNAME20691(G20691,G20449,G2214);
  or GNAME20692(G20692,G2215,G20449);
  nand GNAME20693(G20693,G20449,G2215);
  or GNAME20694(G20694,G2212,G20449);
  nand GNAME20695(G20695,G20449,G2212);
  or GNAME20696(G20696,G2211,G20449);
  nand GNAME20697(G20697,G20449,G2211);
  nand GNAME20698(G20698,G20684,G20685);
  or GNAME20699(G20699,G2208,G20449);
  or GNAME20700(G20700,G2836,G20527);
  nand GNAME20701(G20701,G20699,G20700);
  or GNAME20702(G20702,G2207,G20449);
  or GNAME20703(G20703,G2836,G20528);
  nand GNAME20704(G20704,G20702,G20703);
  or GNAME20705(G20705,G2206,G20449);
  or GNAME20706(G20706,G2836,G20529);
  nand GNAME20707(G20707,G20705,G20706);
  or GNAME20708(G20708,G2205,G20449);
  or GNAME20709(G20709,G2836,G20530);
  nand GNAME20710(G20710,G20708,G20709);
  or GNAME20711(G20711,G2204,G20449);
  or GNAME20712(G20712,G2836,G20531);
  nand GNAME20713(G20713,G20711,G20712);
  or GNAME20714(G20714,G2203,G20449);
  or GNAME20715(G20715,G2836,G20532);
  nand GNAME20716(G20716,G20714,G20715);
  or GNAME20717(G20717,G2202,G20449);
  or GNAME20718(G20718,G2836,G20533);
  nand GNAME20719(G20719,G20717,G20718);
  or GNAME20720(G20720,G2201,G20449);
  nand GNAME20721(G20721,G20449,G2201);
  or GNAME20722(G20722,G2199,G20449);
  nand GNAME20723(G20723,G20449,G2199);
  or GNAME20724(G20724,G2200,G20449);
  nand GNAME20725(G20725,G20449,G2200);
  nand GNAME20726(G20726,G20566,G20675);
  nand GNAME20727(G20727,G20534,G20673,G20674);
  nand GNAME20728(G20728,G20476,G20483);
  or GNAME20729(G20729,G20476,G20483);
  nand GNAME20730(G20730,G20475,G20484);
  or GNAME20731(G20731,G20475,G20484);
  nand GNAME20732(G20732,G20474,G20485);
  or GNAME20733(G20733,G20474,G20485);
  nand GNAME20734(G20734,G20486,G20535);
  or GNAME20735(G20735,G20535,G20486);
  nand GNAME20736(G20736,G20473,G20487);
  or GNAME20737(G20737,G20473,G20487);
  nand GNAME20738(G20738,G20494,G20536);
  or GNAME20739(G20739,G20536,G20494);
  or GNAME20740(G20740,G20539,G20538);
  nand GNAME20741(G20741,G20538,G20539);
  or GNAME20742(G20742,G20542,G20541);
  nand GNAME20743(G20743,G20541,G20542);
  or GNAME20744(G20744,G20545,G20544);
  nand GNAME20745(G20745,G20544,G20545);
  or GNAME20746(G20746,G20548,G20547);
  nand GNAME20747(G20747,G20547,G20548);
  or GNAME20748(G20748,G20551,G20550);
  nand GNAME20749(G20749,G20550,G20551);
  or GNAME20750(G20750,G20554,G20553);
  nand GNAME20751(G20751,G20553,G20554);
  or GNAME20752(G20752,G20557,G20556);
  nand GNAME20753(G20753,G20556,G20557);
  or GNAME20754(G20754,G20560,G20559);
  nand GNAME20755(G20755,G20559,G20560);
  nand GNAME20756(G20756,G20562,G20464);
  or GNAME20757(G20757,G20464,G20562);
  nand GNAME20758(G20758,G20463,G20488);
  or GNAME20759(G20759,G20463,G20488);
  nand GNAME20760(G20760,G20462,G20489);
  or GNAME20761(G20761,G20462,G20489);
  nand GNAME20762(G20762,G20461,G20491);
  or GNAME20763(G20763,G20461,G20491);
  nand GNAME20764(G20764,G20460,G20492);
  or GNAME20765(G20765,G20460,G20492);
  or GNAME20766(G20766,G20563,G20449);
  or GNAME20767(G20767,G2836,G20636);
  not GNAME20768(G20768,G20587);
  not GNAME20769(G20769,G20595);
  not GNAME20770(G20770,G20485);
  not GNAME20771(G20771,G20475);
  not GNAME20772(G20772,G20483);
  nor GNAME20773(G20773,G20776,G20804);
  and GNAME20774(G20774,G20783,G20781,G20782);
  and GNAME20775(G20775,G20778,G20820);
  nor GNAME20776(G20776,G20775,G20774,G20819,G20818);
  not GNAME20777(G20777,G20817);
  not GNAME20778(G20778,G3852);
  not GNAME20779(G20779,G20805);
  or GNAME20780(G20780,G3784,G20777);
  nand GNAME20781(G20781,G3785,G20779,G20780);
  or GNAME20782(G20782,G20820,G20778);
  nand GNAME20783(G20783,G20777,G3784);
  or GNAME20784(G20784,G3280,G20785);
  nor GNAME20785(G20785,G21596,G21597);
  and GNAME20786(G20786,G20802,G20803);
  not GNAME20787(G20787,G3283);
  not GNAME20788(G20788,G59115);
  not GNAME20789(G20789,G3281);
  not GNAME20790(G20790,G3280);
  not GNAME20791(G20791,G3284);
  or GNAME20792(G20792,G59116,G20787);
  nand GNAME20793(G20793,G59117,G20791,G20792);
  or GNAME20794(G20794,G3282,G20788);
  nand GNAME20795(G20795,G20787,G59116);
  nand GNAME20796(G20796,G20795,G20793,G20794);
  or GNAME20797(G20797,G59114,G20789);
  nand GNAME20798(G20798,G20788,G3282);
  nand GNAME20799(G20799,G20798,G20796,G20797);
  nand GNAME20800(G20800,G20790,G59113);
  nand GNAME20801(G20801,G20789,G59114);
  nand GNAME20802(G20802,G20801,G20799,G20800);
  or GNAME20803(G20803,G59113,G20790);
  nand GNAME20804(G20804,G20836,G20837);
  nand GNAME20805(G20805,G20838,G20824);
  not GNAME20806(G20806,G59112);
  not GNAME20807(G20807,G59111);
  not GNAME20808(G20808,G59116);
  and GNAME20809(G20809,G20825,G20855);
  not GNAME20810(G20810,G59110);
  not GNAME20811(G20811,G59115);
  and GNAME20812(G20812,G20828,G20829);
  not GNAME20813(G20813,G59109);
  not GNAME20814(G20814,G59114);
  and GNAME20815(G20815,G20832,G20833);
  not GNAME20816(G20816,G59108);
  nand GNAME20817(G20817,G20856,G20857);
  nand GNAME20818(G20818,G20842,G20843);
  nand GNAME20819(G20819,G20847,G20848);
  nand GNAME20820(G20820,G20852,G20853);
  and GNAME20821(G20821,G20854,G20855);
  not GNAME20822(G20822,G59113);
  nor GNAME20823(G20823,G59117,G20806);
  not GNAME20824(G20824,G20823);
  nand GNAME20825(G20825,G20824,G20854);
  not GNAME20826(G20826,G20809);
  or GNAME20827(G20827,G20826,G20810);
  nand GNAME20828(G20828,G20827,G59115);
  or GNAME20829(G20829,G59110,G20809);
  not GNAME20830(G20830,G20812);
  or GNAME20831(G20831,G20830,G20813);
  nand GNAME20832(G20832,G20831,G59114);
  or GNAME20833(G20833,G59109,G20812);
  not GNAME20834(G20834,G20815);
  or GNAME20835(G20835,G20815,G59108);
  nand GNAME20836(G20836,G20822,G20835);
  or GNAME20837(G20837,G20834,G20816);
  nand GNAME20838(G20838,G20806,G59117);
  or GNAME20839(G20839,G59108,G20822);
  or GNAME20840(G20840,G59113,G20816);
  nand GNAME20841(G20841,G20839,G20840);
  nand GNAME20842(G20842,G20834,G20841);
  nand GNAME20843(G20843,G20815,G20839,G20840);
  or GNAME20844(G20844,G59109,G20814);
  or GNAME20845(G20845,G59114,G20813);
  nand GNAME20846(G20846,G20844,G20845);
  nand GNAME20847(G20847,G20830,G20846);
  nand GNAME20848(G20848,G20812,G20844,G20845);
  or GNAME20849(G20849,G59110,G20811);
  or GNAME20850(G20850,G59115,G20810);
  nand GNAME20851(G20851,G20849,G20850);
  nand GNAME20852(G20852,G20826,G20851);
  nand GNAME20853(G20853,G20809,G20849,G20850);
  or GNAME20854(G20854,G59116,G20807);
  or GNAME20855(G20855,G59111,G20808);
  nand GNAME20856(G20856,G20821,G20823);
  or GNAME20857(G20857,G20823,G20821);
  and GNAME20858(G20858,G21100,G21101);
  and GNAME20859(G20859,G21095,G21096);
  and GNAME20860(G20860,G21089,G21090);
  and GNAME20861(G20861,G21016,G21017);
  not GNAME20862(G20862,G3187);
  not GNAME20863(G20863,G2275);
  not GNAME20864(G20864,G2276);
  not GNAME20865(G20865,G2279);
  not GNAME20866(G20866,G2280);
  not GNAME20867(G20867,G2281);
  not GNAME20868(G20868,G2278);
  not GNAME20869(G20869,G2277);
  not GNAME20870(G20870,G2274);
  and GNAME20871(G20871,G21010,G20983);
  not GNAME20872(G20872,G2273);
  and GNAME20873(G20873,G21006,G20981);
  or GNAME20874(G20874,G21018,G20949);
  not GNAME20875(G20875,G2270);
  and GNAME20876(G20876,G21021,G21022);
  not GNAME20877(G20877,G2269);
  not GNAME20878(G20878,G2268);
  nand GNAME20879(G20879,G21024,G21025);
  nand GNAME20880(G20880,G21028,G21029);
  not GNAME20881(G20881,G2267);
  and GNAME20882(G20882,G21032,G21033);
  not GNAME20883(G20883,G2266);
  and GNAME20884(G20884,G21035,G21036);
  not GNAME20885(G20885,G2265);
  and GNAME20886(G20886,G21038,G21039);
  not GNAME20887(G20887,G2264);
  and GNAME20888(G20888,G21041,G21042);
  not GNAME20889(G20889,G2263);
  and GNAME20890(G20890,G21044,G21045);
  not GNAME20891(G20891,G2262);
  and GNAME20892(G20892,G21047,G21048);
  not GNAME20893(G20893,G2261);
  and GNAME20894(G20894,G21050,G21051);
  not GNAME20895(G20895,G2260);
  and GNAME20896(G20896,G21053,G21054);
  not GNAME20897(G20897,G2259);
  and GNAME20898(G20898,G21056,G21057);
  not GNAME20899(G20899,G2258);
  and GNAME20900(G20900,G21059,G21060);
  not GNAME20901(G20901,G2257);
  and GNAME20902(G20902,G21062,G21063);
  not GNAME20903(G20903,G2256);
  and GNAME20904(G20904,G21065,G21066);
  not GNAME20905(G20905,G2255);
  and GNAME20906(G20906,G21068,G21069);
  not GNAME20907(G20907,G2254);
  and GNAME20908(G20908,G21071,G21072);
  not GNAME20909(G20909,G2253);
  not GNAME20910(G20910,G2252);
  nand GNAME20911(G20911,G21074,G21075);
  nand GNAME20912(G20912,G21078,G21079);
  not GNAME20913(G20913,G2251);
  not GNAME20914(G20914,G2250);
  and GNAME20915(G20915,G20998,G20982);
  nand GNAME20916(G20916,G3187,G2271);
  nand GNAME20917(G20917,G21092,G21093);
  nand GNAME20918(G20918,G21225,G21226);
  nand GNAME20919(G20919,G21132,G21133);
  nand GNAME20920(G20920,G21138,G21139);
  nand GNAME20921(G20921,G21140,G21141);
  nand GNAME20922(G20922,G21145,G21146);
  nand GNAME20923(G20923,G21212,G21213);
  and GNAME20924(G20924,G21124,G21125);
  and GNAME20925(G20925,G21128,G21129);
  and GNAME20926(G20926,G21147,G21148);
  and GNAME20927(G20927,G21151,G21152);
  and GNAME20928(G20928,G21155,G21156);
  and GNAME20929(G20929,G21159,G21160);
  and GNAME20930(G20930,G21163,G21164);
  and GNAME20931(G20931,G21167,G21168);
  and GNAME20932(G20932,G21171,G21172);
  and GNAME20933(G20933,G21175,G21176);
  and GNAME20934(G20934,G21179,G21180);
  and GNAME20935(G20935,G21183,G21184);
  and GNAME20936(G20936,G21189,G21190);
  and GNAME20937(G20937,G21193,G21194);
  and GNAME20938(G20938,G21197,G21198);
  and GNAME20939(G20939,G21201,G21202);
  and GNAME20940(G20940,G21205,G21206);
  and GNAME20941(G20941,G21214,G21215);
  and GNAME20942(G20942,G21218,G21219);
  not GNAME20943(G20943,G2242);
  not GNAME20944(G20944,G2244);
  not GNAME20945(G20945,G2246);
  not GNAME20946(G20946,G2248);
  not GNAME20947(G20947,G2249);
  not GNAME20948(G20948,G2245);
  and GNAME20949(G20949,G21012,G21013);
  and GNAME20950(G20950,G21126,G21127);
  and GNAME20951(G20951,G21130,G21131);
  or GNAME20952(G20952,G21008,G20873);
  nand GNAME20953(G20953,G21004,G20988);
  and GNAME20954(G20954,G21005,G20985);
  and GNAME20955(G20955,G21134,G21135);
  nand GNAME20956(G20956,G21002,G20989);
  and GNAME20957(G20957,G21003,G20988);
  and GNAME20958(G20958,G21136,G21137);
  or GNAME20959(G20959,G21000,G20915);
  and GNAME20960(G20960,G21149,G21150);
  and GNAME20961(G20961,G21153,G21154);
  and GNAME20962(G20962,G21157,G21158);
  and GNAME20963(G20963,G21161,G21162);
  and GNAME20964(G20964,G21165,G21166);
  and GNAME20965(G20965,G21169,G21170);
  and GNAME20966(G20966,G21173,G21174);
  and GNAME20967(G20967,G21177,G21178);
  and GNAME20968(G20968,G21181,G21182);
  and GNAME20969(G20969,G21185,G21186);
  nand GNAME20970(G20970,G20996,G20994);
  and GNAME20971(G20971,G20997,G20991);
  and GNAME20972(G20972,G21187,G21188);
  and GNAME20973(G20973,G21191,G21192);
  and GNAME20974(G20974,G21195,G21196);
  and GNAME20975(G20975,G21199,G21200);
  and GNAME20976(G20976,G21203,G21204);
  and GNAME20977(G20977,G21207,G21208);
  and GNAME20978(G20978,G21216,G21217);
  and GNAME20979(G20979,G21220,G21221);
  nand GNAME20980(G20980,G20995,G20994);
  nand GNAME20981(G20981,G20987,G20863,G20986);
  nand GNAME20982(G20982,G20993,G20865,G20992);
  nand GNAME20983(G20983,G21123,G2274);
  nand GNAME20984(G20984,G20870,G21106,G21107);
  nand GNAME20985(G20985,G21110,G2276);
  or GNAME20986(G20986,G2243,G20862);
  nand GNAME20987(G20987,G20862,G2243);
  nand GNAME20988(G20988,G21122,G2277);
  nand GNAME20989(G20989,G21119,G2278);
  nand GNAME20990(G20990,G20868,G21111,G21112);
  nand GNAME20991(G20991,G21115,G2280);
  or GNAME20992(G20992,G2247,G20862);
  nand GNAME20993(G20993,G20862,G2247);
  nand GNAME20994(G20994,G21118,G2281);
  nand GNAME20995(G20995,G20867,G21116,G21117);
  nand GNAME20996(G20996,G20995,G3187);
  nand GNAME20997(G20997,G20866,G21113,G21114);
  nand GNAME20998(G20998,G20991,G21087);
  nand GNAME20999(G20999,G20992,G20993);
  and GNAME21000(G21000,G20999,G2279);
  not GNAME21001(G21001,G20959);
  nand GNAME21002(G21002,G20990,G20959);
  nand GNAME21003(G21003,G20869,G21120,G21121);
  nand GNAME21004(G21004,G20956,G21003);
  nand GNAME21005(G21005,G20864,G21108,G21109);
  nand GNAME21006(G21006,G20985,G21014);
  nand GNAME21007(G21007,G20986,G20987);
  and GNAME21008(G21008,G21007,G2275);
  not GNAME21009(G21009,G20952);
  nand GNAME21010(G21010,G20984,G20952);
  nand GNAME21011(G21011,G20872,G20871);
  nand GNAME21012(G21012,G21011,G3187);
  or GNAME21013(G21013,G20871,G20872);
  nand GNAME21014(G21014,G20953,G21005);
  nand GNAME21015(G21015,G20981,G21228);
  nand GNAME21016(G21016,G21015,G20985,G21014);
  nand GNAME21017(G21017,G21228,G20873);
  nor GNAME21018(G21018,G2272,G3187);
  not GNAME21019(G21019,G20874);
  or GNAME21020(G21020,G2272,G2270,G21019,G21229);
  nand GNAME21021(G21021,G2270,G21019,G2271);
  nand GNAME21022(G21022,G21020,G3187);
  nand GNAME21023(G21023,G20877,G20876);
  nand GNAME21024(G21024,G21023,G3187);
  or GNAME21025(G21025,G20876,G20877);
  not GNAME21026(G21026,G20879);
  nand GNAME21027(G21027,G20879,G2268);
  nand GNAME21028(G21028,G20862,G21027);
  nand GNAME21029(G21029,G20878,G21026);
  not GNAME21030(G21030,G20880);
  nand GNAME21031(G21031,G20880,G20881);
  nand GNAME21032(G21032,G21031,G3187);
  nand GNAME21033(G21033,G21030,G2267);
  nand GNAME21034(G21034,G20883,G20882);
  nand GNAME21035(G21035,G21034,G3187);
  or GNAME21036(G21036,G20882,G20883);
  nand GNAME21037(G21037,G20885,G20884);
  nand GNAME21038(G21038,G21037,G3187);
  or GNAME21039(G21039,G20884,G20885);
  nand GNAME21040(G21040,G20887,G20886);
  nand GNAME21041(G21041,G21040,G3187);
  or GNAME21042(G21042,G20886,G20887);
  nand GNAME21043(G21043,G20889,G20888);
  nand GNAME21044(G21044,G21043,G3187);
  or GNAME21045(G21045,G20888,G20889);
  nand GNAME21046(G21046,G20891,G20890);
  nand GNAME21047(G21047,G21046,G3187);
  or GNAME21048(G21048,G20890,G20891);
  nand GNAME21049(G21049,G20893,G20892);
  nand GNAME21050(G21050,G21049,G3187);
  or GNAME21051(G21051,G20892,G20893);
  nand GNAME21052(G21052,G20895,G20894);
  nand GNAME21053(G21053,G21052,G3187);
  or GNAME21054(G21054,G20894,G20895);
  nand GNAME21055(G21055,G20897,G20896);
  nand GNAME21056(G21056,G21055,G3187);
  or GNAME21057(G21057,G20896,G20897);
  nand GNAME21058(G21058,G20899,G20898);
  nand GNAME21059(G21059,G21058,G3187);
  or GNAME21060(G21060,G20898,G20899);
  nand GNAME21061(G21061,G20901,G20900);
  nand GNAME21062(G21062,G21061,G3187);
  or GNAME21063(G21063,G20900,G20901);
  nand GNAME21064(G21064,G20903,G20902);
  nand GNAME21065(G21065,G21064,G3187);
  or GNAME21066(G21066,G20902,G20903);
  nand GNAME21067(G21067,G20905,G20904);
  nand GNAME21068(G21068,G21067,G3187);
  or GNAME21069(G21069,G20904,G20905);
  nand GNAME21070(G21070,G20907,G20906);
  nand GNAME21071(G21071,G21070,G3187);
  or GNAME21072(G21072,G20906,G20907);
  nand GNAME21073(G21073,G20909,G20908);
  nand GNAME21074(G21074,G21073,G3187);
  or GNAME21075(G21075,G20908,G20909);
  not GNAME21076(G21076,G20911);
  nand GNAME21077(G21077,G20911,G2252);
  nand GNAME21078(G21078,G20862,G21077);
  nand GNAME21079(G21079,G20910,G21076);
  not GNAME21080(G21080,G20912);
  nand GNAME21081(G21081,G21080,G2251);
  nand GNAME21082(G21082,G20862,G21081);
  nand GNAME21083(G21083,G20913,G20912);
  nand GNAME21084(G21084,G2250,G21082,G21083);
  nand GNAME21085(G21085,G21083,G3187);
  nand GNAME21086(G21086,G21081,G20914,G21085);
  nand GNAME21087(G21087,G20970,G20997);
  nand GNAME21088(G21088,G20982,G21227);
  nand GNAME21089(G21089,G21088,G20991,G21087);
  nand GNAME21090(G21090,G21227,G20915);
  nand GNAME21091(G21091,G21019,G2271);
  nand GNAME21092(G21092,G20862,G21091);
  or GNAME21093(G21093,G2272,G21019);
  nand GNAME21094(G21094,G20916,G20917);
  nand GNAME21095(G21095,G21094,G21224);
  nand GNAME21096(G21096,G21222,G21223,G20916,G20917);
  or GNAME21097(G21097,G2272,G20916);
  nand GNAME21098(G21098,G21097,G3187);
  nand GNAME21099(G21099,G20916,G2271);
  nand GNAME21100(G21100,G21099,G20874,G21098);
  or GNAME21101(G21101,G21229,G20917);
  not GNAME21102(G21102,G20980);
  nand GNAME21103(G21103,G20983,G20984);
  nand GNAME21104(G21104,G20989,G20990);
  nand GNAME21105(G21105,G21084,G21086);
  nand GNAME21106(G21106,G20943,G3187);
  nand GNAME21107(G21107,G20862,G2242);
  nand GNAME21108(G21108,G20944,G3187);
  nand GNAME21109(G21109,G20862,G2244);
  nand GNAME21110(G21110,G21108,G21109);
  nand GNAME21111(G21111,G20945,G3187);
  nand GNAME21112(G21112,G20862,G2246);
  nand GNAME21113(G21113,G20946,G3187);
  nand GNAME21114(G21114,G20862,G2248);
  nand GNAME21115(G21115,G21113,G21114);
  nand GNAME21116(G21116,G20947,G3187);
  nand GNAME21117(G21117,G20862,G2249);
  nand GNAME21118(G21118,G21116,G21117);
  nand GNAME21119(G21119,G21111,G21112);
  nand GNAME21120(G21120,G20948,G3187);
  nand GNAME21121(G21121,G20862,G2245);
  nand GNAME21122(G21122,G21120,G21121);
  nand GNAME21123(G21123,G21106,G21107);
  or GNAME21124(G21124,G2272,G20862);
  nand GNAME21125(G21125,G20862,G2272);
  nand GNAME21126(G21126,G20924,G20949);
  or GNAME21127(G21127,G20949,G20924);
  nand GNAME21128(G21128,G20872,G3187);
  nand GNAME21129(G21129,G20862,G2273);
  nand GNAME21130(G21130,G20871,G20925);
  or GNAME21131(G21131,G20871,G20925);
  nand GNAME21132(G21132,G20952,G21103);
  nand GNAME21133(G21133,G21009,G20983,G20984);
  or GNAME21134(G21134,G20954,G20953);
  nand GNAME21135(G21135,G20953,G20954);
  or GNAME21136(G21136,G20957,G20956);
  nand GNAME21137(G21137,G20956,G20957);
  nand GNAME21138(G21138,G20959,G21104);
  nand GNAME21139(G21139,G21001,G20989,G20990);
  nand GNAME21140(G21140,G21105,G3187);
  nand GNAME21141(G21141,G20862,G21084,G21086);
  nand GNAME21142(G21142,G20913,G3187);
  nand GNAME21143(G21143,G20862,G2251);
  nand GNAME21144(G21144,G21142,G21143);
  nand GNAME21145(G21145,G20912,G21144);
  nand GNAME21146(G21146,G21080,G21142,G21143);
  nand GNAME21147(G21147,G20910,G3187);
  nand GNAME21148(G21148,G20862,G2252);
  nand GNAME21149(G21149,G21076,G20926);
  or GNAME21150(G21150,G21076,G20926);
  nand GNAME21151(G21151,G20909,G3187);
  nand GNAME21152(G21152,G20862,G2253);
  nand GNAME21153(G21153,G20908,G20927);
  or GNAME21154(G21154,G20908,G20927);
  nand GNAME21155(G21155,G20907,G3187);
  nand GNAME21156(G21156,G20862,G2254);
  nand GNAME21157(G21157,G20906,G20928);
  or GNAME21158(G21158,G20906,G20928);
  nand GNAME21159(G21159,G20905,G3187);
  nand GNAME21160(G21160,G20862,G2255);
  nand GNAME21161(G21161,G20904,G20929);
  or GNAME21162(G21162,G20904,G20929);
  nand GNAME21163(G21163,G20903,G3187);
  nand GNAME21164(G21164,G20862,G2256);
  nand GNAME21165(G21165,G20902,G20930);
  or GNAME21166(G21166,G20902,G20930);
  nand GNAME21167(G21167,G20901,G3187);
  nand GNAME21168(G21168,G20862,G2257);
  nand GNAME21169(G21169,G20900,G20931);
  or GNAME21170(G21170,G20900,G20931);
  nand GNAME21171(G21171,G20899,G3187);
  nand GNAME21172(G21172,G20862,G2258);
  nand GNAME21173(G21173,G20898,G20932);
  or GNAME21174(G21174,G20898,G20932);
  nand GNAME21175(G21175,G20897,G3187);
  nand GNAME21176(G21176,G20862,G2259);
  nand GNAME21177(G21177,G20896,G20933);
  or GNAME21178(G21178,G20896,G20933);
  nand GNAME21179(G21179,G20895,G3187);
  nand GNAME21180(G21180,G20862,G2260);
  nand GNAME21181(G21181,G20894,G20934);
  or GNAME21182(G21182,G20894,G20934);
  nand GNAME21183(G21183,G20893,G3187);
  nand GNAME21184(G21184,G20862,G2261);
  nand GNAME21185(G21185,G20892,G20935);
  or GNAME21186(G21186,G20892,G20935);
  or GNAME21187(G21187,G20971,G20970);
  nand GNAME21188(G21188,G20970,G20971);
  nand GNAME21189(G21189,G20891,G3187);
  nand GNAME21190(G21190,G20862,G2262);
  nand GNAME21191(G21191,G20890,G20936);
  or GNAME21192(G21192,G20890,G20936);
  nand GNAME21193(G21193,G20889,G3187);
  nand GNAME21194(G21194,G20862,G2263);
  nand GNAME21195(G21195,G20888,G20937);
  or GNAME21196(G21196,G20888,G20937);
  nand GNAME21197(G21197,G20887,G3187);
  nand GNAME21198(G21198,G20862,G2264);
  nand GNAME21199(G21199,G20886,G20938);
  or GNAME21200(G21200,G20886,G20938);
  nand GNAME21201(G21201,G20885,G3187);
  nand GNAME21202(G21202,G20862,G2265);
  nand GNAME21203(G21203,G20884,G20939);
  or GNAME21204(G21204,G20884,G20939);
  nand GNAME21205(G21205,G20883,G3187);
  nand GNAME21206(G21206,G20862,G2266);
  nand GNAME21207(G21207,G20882,G20940);
  or GNAME21208(G21208,G20882,G20940);
  nand GNAME21209(G21209,G20881,G3187);
  nand GNAME21210(G21210,G20862,G2267);
  nand GNAME21211(G21211,G21209,G21210);
  nand GNAME21212(G21212,G20880,G21211);
  nand GNAME21213(G21213,G21030,G21209,G21210);
  nand GNAME21214(G21214,G20878,G3187);
  nand GNAME21215(G21215,G20862,G2268);
  nand GNAME21216(G21216,G21026,G20941);
  or GNAME21217(G21217,G21026,G20941);
  nand GNAME21218(G21218,G20877,G3187);
  nand GNAME21219(G21219,G20862,G2269);
  nand GNAME21220(G21220,G20876,G20942);
  or GNAME21221(G21221,G20876,G20942);
  nand GNAME21222(G21222,G20875,G3187);
  nand GNAME21223(G21223,G20862,G2270);
  nand GNAME21224(G21224,G21222,G21223);
  nand GNAME21225(G21225,G20980,G3187);
  nand GNAME21226(G21226,G20862,G21102);
  not GNAME21227(G21227,G21000);
  not GNAME21228(G21228,G21008);
  not GNAME21229(G21229,G20916);
  and GNAME21230(G21230,G21324,G21325);
  not GNAME21231(G21231,G20516);
  not GNAME21232(G21232,G2134);
  and GNAME21233(G21233,G2135,G20516);
  and GNAME21234(G21234,G21304,G21305);
  not GNAME21235(G21235,G2133);
  and GNAME21236(G21236,G21307,G21308);
  not GNAME21237(G21237,G2132);
  and GNAME21238(G21238,G21310,G21311);
  not GNAME21239(G21239,G2131);
  and GNAME21240(G21240,G21313,G21314);
  not GNAME21241(G21241,G2130);
  not GNAME21242(G21242,G2129);
  and GNAME21243(G21243,G21316,G21317);
  and GNAME21244(G21244,G21320,G21321);
  not GNAME21245(G21245,G20500);
  nor GNAME21246(G21246,G21292,G21245);
  not GNAME21247(G21247,G20558);
  not GNAME21248(G21248,G20561);
  nand GNAME21249(G21249,G20561,G21246,G20558);
  and GNAME21250(G21250,G20555,G21383);
  not GNAME21251(G21251,G20546);
  not GNAME21252(G21252,G20549);
  nand GNAME21253(G21253,G20549,G21250,G20546);
  and GNAME21254(G21254,G20543,G21384);
  not GNAME21255(G21255,G20537);
  not GNAME21256(G21256,G20540);
  not GNAME21257(G21257,G20498);
  nand GNAME21258(G21258,G20540,G21254,G20537);
  nand GNAME21259(G21259,G21301,G20498,G20499);
  and GNAME21260(G21260,G20497,G21385);
  not GNAME21261(G21261,G20496);
  and GNAME21262(G21262,G21260,G20496);
  not GNAME21263(G21263,G20495);
  and GNAME21264(G21264,G21322,G21244);
  nand GNAME21265(G21265,G21328,G21329);
  nand GNAME21266(G21266,G21330,G21331);
  nand GNAME21267(G21267,G21332,G21333);
  nand GNAME21268(G21268,G21334,G21335);
  nand GNAME21269(G21269,G21336,G21337);
  nand GNAME21270(G21270,G21338,G21339);
  nand GNAME21271(G21271,G21340,G21341);
  nand GNAME21272(G21272,G21342,G21343);
  nand GNAME21273(G21273,G21344,G21345);
  nand GNAME21274(G21274,G21346,G21347);
  nand GNAME21275(G21275,G21348,G21349);
  nand GNAME21276(G21276,G21350,G21351);
  nand GNAME21277(G21277,G21352,G21353);
  nand GNAME21278(G21278,G21354,G21355);
  nand GNAME21279(G21279,G21356,G21357);
  nand GNAME21280(G21280,G21358,G21359);
  and GNAME21281(G21281,G21326,G21327);
  and GNAME21282(G21282,G21362,G21363);
  and GNAME21283(G21283,G21366,G21367);
  and GNAME21284(G21284,G21370,G21371);
  and GNAME21285(G21285,G21374,G21375);
  and GNAME21286(G21286,G21378,G21379);
  nand GNAME21287(G21287,G21262,G20495);
  and GNAME21288(G21288,G20499,G21301);
  and GNAME21289(G21289,G21254,G20540);
  and GNAME21290(G21290,G21250,G20549);
  and GNAME21291(G21291,G21246,G20561);
  nor GNAME21292(G21292,G21382,G21264);
  and GNAME21293(G21293,G21360,G21361);
  not GNAME21294(G21294,G20445);
  and GNAME21295(G21295,G21364,G21365);
  and GNAME21296(G21296,G21368,G21369);
  and GNAME21297(G21297,G21372,G21373);
  and GNAME21298(G21298,G21376,G21377);
  and GNAME21299(G21299,G21380,G21381);
  not GNAME21300(G21300,G21292);
  not GNAME21301(G21301,G21258);
  nand GNAME21302(G21302,G20501,G2128);
  or GNAME21303(G21303,G20481,G2134);
  nand GNAME21304(G21304,G21303,G21233);
  nand GNAME21305(G21305,G20481,G2134);
  nand GNAME21306(G21306,G21235,G21234);
  nand GNAME21307(G21307,G21306,G20444);
  or GNAME21308(G21308,G21234,G21235);
  nand GNAME21309(G21309,G21237,G21236);
  nand GNAME21310(G21310,G21309,G20504);
  or GNAME21311(G21311,G21236,G21237);
  nand GNAME21312(G21312,G21239,G21238);
  nand GNAME21313(G21313,G21312,G20503);
  or GNAME21314(G21314,G21238,G21239);
  nand GNAME21315(G21315,G21241,G21240);
  nand GNAME21316(G21316,G21315,G20502);
  or GNAME21317(G21317,G21240,G21241);
  not GNAME21318(G21318,G21243);
  or GNAME21319(G21319,G21243,G21242);
  nand GNAME21320(G21320,G21294,G21319);
  or GNAME21321(G21321,G2129,G21318);
  or GNAME21322(G21322,G2128,G20501);
  and GNAME21323(G21323,G21302,G21322);
  or GNAME21324(G21324,G21323,G21244);
  nand GNAME21325(G21325,G21302,G21264);
  nand GNAME21326(G21326,G21232,G20481);
  or GNAME21327(G21327,G20481,G21232);
  nand GNAME21328(G21328,G21233,G21281);
  or GNAME21329(G21329,G21233,G21281);
  or GNAME21330(G21330,G2135,G21231);
  nand GNAME21331(G21331,G21231,G2135);
  nand GNAME21332(G21332,G21287,G20447);
  or GNAME21333(G21333,G20447,G21287);
  or GNAME21334(G21334,G21262,G21263);
  nand GNAME21335(G21335,G21263,G21262);
  or GNAME21336(G21336,G21260,G21261);
  nand GNAME21337(G21337,G21261,G21260);
  or GNAME21338(G21338,G20497,G21259);
  nand GNAME21339(G21339,G21259,G20497);
  or GNAME21340(G21340,G21288,G21257);
  nand GNAME21341(G21341,G21257,G21288);
  or GNAME21342(G21342,G20499,G21258);
  nand GNAME21343(G21343,G21258,G20499);
  or GNAME21344(G21344,G21289,G21255);
  nand GNAME21345(G21345,G21255,G21289);
  or GNAME21346(G21346,G21254,G21256);
  nand GNAME21347(G21347,G21256,G21254);
  or GNAME21348(G21348,G20543,G21253);
  nand GNAME21349(G21349,G21253,G20543);
  or GNAME21350(G21350,G21290,G21251);
  nand GNAME21351(G21351,G21251,G21290);
  or GNAME21352(G21352,G21250,G21252);
  nand GNAME21353(G21353,G21252,G21250);
  or GNAME21354(G21354,G20555,G21249);
  nand GNAME21355(G21355,G21249,G20555);
  or GNAME21356(G21356,G21291,G21247);
  nand GNAME21357(G21357,G21247,G21291);
  or GNAME21358(G21358,G21246,G21248);
  nand GNAME21359(G21359,G21248,G21246);
  or GNAME21360(G21360,G21292,G21245);
  or GNAME21361(G21361,G20500,G21300);
  or GNAME21362(G21362,G2129,G21294);
  or GNAME21363(G21363,G20445,G21242);
  nand GNAME21364(G21364,G21243,G21282);
  or GNAME21365(G21365,G21243,G21282);
  nand GNAME21366(G21366,G21241,G20502);
  or GNAME21367(G21367,G20502,G21241);
  nand GNAME21368(G21368,G21240,G21283);
  or GNAME21369(G21369,G21240,G21283);
  nand GNAME21370(G21370,G21239,G20503);
  or GNAME21371(G21371,G20503,G21239);
  nand GNAME21372(G21372,G21238,G21284);
  or GNAME21373(G21373,G21238,G21284);
  nand GNAME21374(G21374,G21237,G20504);
  or GNAME21375(G21375,G20504,G21237);
  nand GNAME21376(G21376,G21236,G21285);
  or GNAME21377(G21377,G21236,G21285);
  nand GNAME21378(G21378,G21235,G20444);
  or GNAME21379(G21379,G20444,G21235);
  nand GNAME21380(G21380,G21234,G21286);
  or GNAME21381(G21381,G21234,G21286);
  not GNAME21382(G21382,G21302);
  not GNAME21383(G21383,G21249);
  not GNAME21384(G21384,G21253);
  not GNAME21385(G21385,G21259);
  not GNAME21386(G21386,G3278);
  not GNAME21387(G21387,G3279);
  not GNAME21388(G21388,G2119);
  not GNAME21389(G21389,G3277);
  nor GNAME21390(G21390,G21430,G21516);
  and GNAME21391(G21391,G21483,G21514);
  nor GNAME21392(G21392,G21432,G21513);
  and GNAME21393(G21393,G21591,G21511);
  nand GNAME21394(G21394,G21484,G3869);
  not GNAME21395(G21395,G2304);
  not GNAME21396(G21396,G2305);
  not GNAME21397(G21397,G2302);
  and GNAME21398(G21398,G21485,G2302);
  not GNAME21399(G21399,G2301);
  not GNAME21400(G21400,G2300);
  and GNAME21401(G21401,G2300,G21398,G2301);
  and GNAME21402(G21402,G2299,G21401);
  not GNAME21403(G21403,G2297);
  not GNAME21404(G21404,G2298);
  and GNAME21405(G21405,G2298,G21402,G2297);
  not GNAME21406(G21406,G2296);
  nand GNAME21407(G21407,G21405,G2296);
  not GNAME21408(G21408,G2295);
  not GNAME21409(G21409,G2294);
  and GNAME21410(G21410,G2294,G21486,G2295);
  not GNAME21411(G21411,G2292);
  and GNAME21412(G21412,G2292,G2293,G21410);
  not GNAME21413(G21413,G2290);
  and GNAME21414(G21414,G2290,G2291,G21412);
  not GNAME21415(G21415,G2289);
  and GNAME21416(G21416,G21488,G21489);
  not GNAME21417(G21417,G2312);
  and GNAME21418(G21418,G21491,G21492);
  not GNAME21419(G21419,G2311);
  and GNAME21420(G21420,G21494,G21495);
  not GNAME21421(G21421,G2310);
  and GNAME21422(G21422,G21497,G21498);
  not GNAME21423(G21423,G2309);
  and GNAME21424(G21424,G21500,G21501);
  not GNAME21425(G21425,G2308);
  and GNAME21426(G21426,G21503,G21504);
  not GNAME21427(G21427,G2307);
  and GNAME21428(G21428,G21506,G21507);
  not GNAME21429(G21429,G2306);
  and GNAME21430(G21430,G3291,G21467,G3292);
  and GNAME21431(G21431,G3290,G21430);
  and GNAME21432(G21432,G21431,G3289,G3288);
  and GNAME21433(G21433,G3287,G21432);
  nand GNAME21434(G21434,G21518,G21519);
  nand GNAME21435(G21435,G21520,G21521);
  nand GNAME21436(G21436,G21522,G21523);
  nand GNAME21437(G21437,G21524,G21525);
  nand GNAME21438(G21438,G21526,G21527);
  nand GNAME21439(G21439,G21528,G21529);
  nand GNAME21440(G21440,G21530,G21531);
  nand GNAME21441(G21441,G21532,G21533);
  nand GNAME21442(G21442,G21534,G21535);
  nand GNAME21443(G21443,G21536,G21537);
  nand GNAME21444(G21444,G21538,G21539);
  nand GNAME21445(G21445,G21558,G21559);
  nand GNAME21446(G21446,G21574,G21575);
  nand GNAME21447(G21447,G21576,G21577);
  nand GNAME21448(G21448,G21578,G21579);
  nand GNAME21449(G21449,G21580,G21581);
  nand GNAME21450(G21450,G21582,G21583);
  nand GNAME21451(G21451,G21584,G21585);
  nand GNAME21452(G21452,G21586,G21587);
  nand GNAME21453(G21453,G21588,G21589);
  and GNAME21454(G21454,G21542,G21543);
  and GNAME21455(G21455,G21546,G21547);
  and GNAME21456(G21456,G21550,G21551);
  and GNAME21457(G21457,G21554,G21555);
  and GNAME21458(G21458,G21560,G21561);
  and GNAME21459(G21459,G21564,G21565);
  and GNAME21460(G21460,G21568,G21569);
  and GNAME21461(G21461,G21572,G21573);
  and GNAME21462(G21462,G21402,G2298);
  and GNAME21463(G21463,G21398,G2301);
  nand GNAME21464(G21464,G21433,G3286);
  not GNAME21465(G21465,G2303);
  nand GNAME21466(G21466,G21480,G3869);
  nand GNAME21467(G21467,G21509,G21510);
  and GNAME21468(G21468,G21540,G21541);
  and GNAME21469(G21469,G21544,G21545);
  and GNAME21470(G21470,G21548,G21549);
  and GNAME21471(G21471,G21552,G21553);
  and GNAME21472(G21472,G21556,G21557);
  and GNAME21473(G21473,G2305,G3869);
  and GNAME21474(G21474,G21562,G21563);
  and GNAME21475(G21475,G21566,G21567);
  and GNAME21476(G21476,G21570,G21571);
  and GNAME21477(G21477,G2291,G21412);
  and GNAME21478(G21478,G2293,G21410);
  and GNAME21479(G21479,G21486,G2295);
  nand GNAME21480(G21480,G2304,G2305);
  not GNAME21481(G21481,G21410);
  not GNAME21482(G21482,G21412);
  not GNAME21483(G21483,G21431);
  nand GNAME21484(G21484,G21465,G21480);
  not GNAME21485(G21485,G21394);
  not GNAME21486(G21486,G21407);
  or GNAME21487(G21487,G2289,G2313);
  nand GNAME21488(G21488,G21487,G21414);
  nand GNAME21489(G21489,G2313,G2289);
  nand GNAME21490(G21490,G21417,G21416);
  nand GNAME21491(G21491,G21490,G2288);
  or GNAME21492(G21492,G21416,G21417);
  nand GNAME21493(G21493,G21419,G21418);
  nand GNAME21494(G21494,G21493,G2287);
  or GNAME21495(G21495,G21418,G21419);
  nand GNAME21496(G21496,G21421,G21420);
  nand GNAME21497(G21497,G21496,G2286);
  or GNAME21498(G21498,G21420,G21421);
  nand GNAME21499(G21499,G21423,G21422);
  nand GNAME21500(G21500,G21499,G2285);
  or GNAME21501(G21501,G21422,G21423);
  nand GNAME21502(G21502,G21425,G21424);
  nand GNAME21503(G21503,G21502,G2284);
  or GNAME21504(G21504,G21424,G21425);
  nand GNAME21505(G21505,G21427,G21426);
  nand GNAME21506(G21506,G21505,G2283);
  or GNAME21507(G21507,G21426,G21427);
  nand GNAME21508(G21508,G21429,G21428);
  nand GNAME21509(G21509,G21508,G3293);
  or GNAME21510(G21510,G21428,G21429);
  or GNAME21511(G21511,G3287,G21432);
  and GNAME21512(G21512,G3289,G21431);
  nor GNAME21513(G21513,G21512,G3288);
  or GNAME21514(G21514,G3290,G21430);
  and GNAME21515(G21515,G21467,G3292);
  nor GNAME21516(G21516,G21515,G3291);
  not GNAME21517(G21517,G21466);
  nand GNAME21518(G21518,G21406,G21405);
  or GNAME21519(G21519,G21405,G21406);
  or GNAME21520(G21520,G21462,G21403);
  nand GNAME21521(G21521,G21403,G21462);
  or GNAME21522(G21522,G21402,G21404);
  nand GNAME21523(G21523,G21404,G21402);
  or GNAME21524(G21524,G2299,G21590);
  nand GNAME21525(G21525,G21590,G2299);
  or GNAME21526(G21526,G21463,G21400);
  nand GNAME21527(G21527,G21400,G21463);
  or GNAME21528(G21528,G21398,G21399);
  nand GNAME21529(G21529,G21399,G21398);
  nand GNAME21530(G21530,G21394,G2302);
  nand GNAME21531(G21531,G21397,G21485);
  nand GNAME21532(G21532,G21464,G2282);
  or GNAME21533(G21533,G2282,G21464);
  nand GNAME21534(G21534,G21591,G3286);
  or GNAME21535(G21535,G3286,G21591);
  nand GNAME21536(G21536,G21466,G2303);
  nand GNAME21537(G21537,G21465,G21517);
  or GNAME21538(G21538,G3289,G21483);
  nand GNAME21539(G21539,G21483,G3289);
  nand GNAME21540(G21540,G21467,G3292);
  or GNAME21541(G21541,G3292,G21467);
  nand GNAME21542(G21542,G21429,G3293);
  or GNAME21543(G21543,G3293,G21429);
  nand GNAME21544(G21544,G21428,G21454);
  or GNAME21545(G21545,G21428,G21454);
  nand GNAME21546(G21546,G21427,G2283);
  or GNAME21547(G21547,G2283,G21427);
  nand GNAME21548(G21548,G21426,G21455);
  or GNAME21549(G21549,G21426,G21455);
  nand GNAME21550(G21550,G21425,G2284);
  or GNAME21551(G21551,G2284,G21425);
  nand GNAME21552(G21552,G21424,G21456);
  or GNAME21553(G21553,G21424,G21456);
  nand GNAME21554(G21554,G21423,G2285);
  or GNAME21555(G21555,G2285,G21423);
  nand GNAME21556(G21556,G21422,G21457);
  or GNAME21557(G21557,G21422,G21457);
  or GNAME21558(G21558,G21473,G21395);
  nand GNAME21559(G21559,G21395,G21473);
  nand GNAME21560(G21560,G21421,G2286);
  or GNAME21561(G21561,G2286,G21421);
  nand GNAME21562(G21562,G21420,G21458);
  or GNAME21563(G21563,G21420,G21458);
  nand GNAME21564(G21564,G21419,G2287);
  or GNAME21565(G21565,G2287,G21419);
  nand GNAME21566(G21566,G21418,G21459);
  or GNAME21567(G21567,G21418,G21459);
  nand GNAME21568(G21568,G21417,G2288);
  or GNAME21569(G21569,G2288,G21417);
  nand GNAME21570(G21570,G21416,G21460);
  or GNAME21571(G21571,G21416,G21460);
  nand GNAME21572(G21572,G21415,G21414);
  or GNAME21573(G21573,G21414,G21415);
  nand GNAME21574(G21574,G2313,G21461);
  or GNAME21575(G21575,G2313,G21461);
  or GNAME21576(G21576,G21477,G21413);
  nand GNAME21577(G21577,G21413,G21477);
  or GNAME21578(G21578,G2291,G21482);
  nand GNAME21579(G21579,G21482,G2291);
  or GNAME21580(G21580,G21478,G21411);
  nand GNAME21581(G21581,G21411,G21478);
  or GNAME21582(G21582,G2293,G21481);
  nand GNAME21583(G21583,G21481,G2293);
  or GNAME21584(G21584,G21479,G21409);
  nand GNAME21585(G21585,G21409,G21479);
  nand GNAME21586(G21586,G21407,G2295);
  nand GNAME21587(G21587,G21408,G21486);
  or GNAME21588(G21588,G3869,G21396);
  nand GNAME21589(G21589,G21396,G3869);
  not GNAME21590(G21590,G21401);
  not GNAME21591(G21591,G21433);
  nand GNAME21592(G21592,G21594,G21595);
  not GNAME21593(G21593,G59118);
  nand GNAME21594(G21594,G21593,G59119);
  or GNAME21595(G21595,G59119,G21593);
  not GNAME21596(G21596,G3281);
  not GNAME21597(G21597,G3282);
  nand GNAME21598(G21598,G21625,G21628,G21629);
  not GNAME21599(G21599,G8135);
  not GNAME21600(G21600,G8139);
  not GNAME21601(G21601,G8146);
  not GNAME21602(G21602,G8137);
  not GNAME21603(G21603,G8144);
  not GNAME21604(G21604,G8134);
  not GNAME21605(G21605,G8140);
  nand GNAME21606(G21606,G21607,G21624);
  or GNAME21607(G21607,G8142,G21599);
  or GNAME21608(G21608,G8147,G21600);
  nand GNAME21609(G21609,G8148,G21605,G21608);
  or GNAME21610(G21610,G8138,G21601);
  nand GNAME21611(G21611,G21600,G8147);
  nand GNAME21612(G21612,G21611,G21609,G21610);
  or GNAME21613(G21613,G8145,G21602);
  nand GNAME21614(G21614,G21601,G8138);
  nand GNAME21615(G21615,G21614,G21612,G21613);
  or GNAME21616(G21616,G8136,G21603);
  nand GNAME21617(G21617,G21602,G8145);
  nand GNAME21618(G21618,G21617,G21615,G21616);
  or GNAME21619(G21619,G8143,G21599);
  nand GNAME21620(G21620,G21603,G8136);
  nand GNAME21621(G21621,G21620,G21618,G21619);
  or GNAME21622(G21622,G8143,G8142);
  nand GNAME21623(G21623,G21599,G21622);
  nand GNAME21624(G21624,G21623,G21621);
  nand GNAME21625(G21625,G21606,G21626,G21627);
  nand GNAME21626(G21626,G21604,G8141);
  or GNAME21627(G21627,G8141,G21604);
  nand GNAME21628(G21628,G21604,G8141,G8133);
  or GNAME21629(G21629,G21604,G8141,G8133);
  and GNAME21630(G21630,G21795,G21796);
  and GNAME21631(G21631,G21754,G21792);
  and GNAME21632(G21632,G21744,G21790);
  and GNAME21633(G21633,G21756,G21763);
  not GNAME21634(G21634,G8788);
  not GNAME21635(G21635,G8189);
  not GNAME21636(G21636,G8190);
  nor GNAME21637(G21637,G21753,G21665);
  nor GNAME21638(G21638,G21664,G21754);
  nor GNAME21639(G21639,G21663,G21739);
  nor GNAME21640(G21640,G21755,G21661,G21662);
  nor GNAME21641(G21641,G21660,G21756);
  not GNAME21642(G21642,G8188);
  not GNAME21643(G21643,G8187);
  not GNAME21644(G21644,G8186);
  not GNAME21645(G21645,G8185);
  not GNAME21646(G21646,G8184);
  not GNAME21647(G21647,G8183);
  not GNAME21648(G21648,G8182);
  not GNAME21649(G21649,G8181);
  nor GNAME21650(G21650,G21725,G21685);
  nor GNAME21651(G21651,G21912,G21683,G21684);
  nor GNAME21652(G21652,G21682,G21740);
  nor GNAME21653(G21653,G21787,G21680,G21681);
  nor GNAME21654(G21654,G21679,G21741);
  nor GNAME21655(G21655,G21788,G21677,G21678);
  nor GNAME21656(G21656,G21676,G21742);
  nor GNAME21657(G21657,G21789,G21674,G21675);
  or GNAME21658(G21658,G21743,G21672,G21673);
  and GNAME21659(G21659,G21774,G21746);
  and GNAME21660(G21660,G21802,G21803);
  and GNAME21661(G21661,G21816,G21817);
  and GNAME21662(G21662,G21818,G21819);
  and GNAME21663(G21663,G21804,G21805);
  and GNAME21664(G21664,G21806,G21807);
  and GNAME21665(G21665,G21814,G21815);
  nand GNAME21666(G21666,G21826,G21827);
  nand GNAME21667(G21667,G21828,G21829);
  nand GNAME21668(G21668,G21830,G21831);
  nand GNAME21669(G21669,G21832,G21833);
  nand GNAME21670(G21670,G21834,G21835);
  and GNAME21671(G21671,G21839,G21840);
  and GNAME21672(G21672,G21877,G21878);
  and GNAME21673(G21673,G21879,G21880);
  and GNAME21674(G21674,G21873,G21874);
  and GNAME21675(G21675,G21875,G21876);
  and GNAME21676(G21676,G21841,G21842);
  and GNAME21677(G21677,G21869,G21870);
  and GNAME21678(G21678,G21871,G21872);
  and GNAME21679(G21679,G21843,G21844);
  and GNAME21680(G21680,G21865,G21866);
  and GNAME21681(G21681,G21867,G21868);
  and GNAME21682(G21682,G21845,G21846);
  and GNAME21683(G21683,G21861,G21862);
  and GNAME21684(G21684,G21863,G21864);
  and GNAME21685(G21685,G21859,G21860);
  nand GNAME21686(G21686,G21883,G21884);
  nand GNAME21687(G21687,G21885,G21886);
  nand GNAME21688(G21688,G21887,G21888);
  nand GNAME21689(G21689,G21889,G21890);
  nand GNAME21690(G21690,G21891,G21892);
  nand GNAME21691(G21691,G21893,G21894);
  nand GNAME21692(G21692,G21895,G21896);
  nand GNAME21693(G21693,G21897,G21898);
  nand GNAME21694(G21694,G21899,G21900);
  nand GNAME21695(G21695,G21901,G21902);
  nand GNAME21696(G21696,G21905,G21906);
  nand GNAME21697(G21697,G21907,G21908);
  nand GNAME21698(G21698,G21909,G21910);
  nand GNAME21699(G21699,G21923,G21924);
  nand GNAME21700(G21700,G21881,G21882);
  nand GNAME21701(G21701,G21915,G21916);
  nand GNAME21702(G21702,G21921,G21922);
  not GNAME21703(G21703,G8172);
  not GNAME21704(G21704,G8179);
  not GNAME21705(G21705,G8180);
  not GNAME21706(G21706,G8171);
  nand GNAME21707(G21707,G21759,G21757);
  and GNAME21708(G21708,G21761,G21760);
  and GNAME21709(G21709,G21824,G21825);
  nand GNAME21710(G21710,G21758,G21757);
  not GNAME21711(G21711,G8149);
  not GNAME21712(G21712,G8169);
  not GNAME21713(G21713,G8168);
  not GNAME21714(G21714,G8167);
  not GNAME21715(G21715,G8165);
  nor GNAME21716(G21716,G21671,G21658);
  nor GNAME21717(G21717,G21673,G21743);
  nor GNAME21718(G21718,G21674,G21789);
  nor GNAME21719(G21719,G21677,G21788);
  nor GNAME21720(G21720,G21680,G21787);
  nand GNAME21721(G21721,G21751,G21749);
  and GNAME21722(G21722,G21752,G21748);
  and GNAME21723(G21723,G21903,G21904);
  nor GNAME21724(G21724,G21683,G21912);
  and GNAME21725(G21725,G21786,G21764);
  and GNAME21726(G21726,G21911,G21912);
  nand GNAME21727(G21727,G21784,G21747);
  and GNAME21728(G21728,G21785,G21764);
  and GNAME21729(G21729,G21913,G21914);
  and GNAME21730(G21730,G21782,G21768);
  nand GNAME21731(G21731,G21780,G21769);
  and GNAME21732(G21732,G21781,G21768);
  and GNAME21733(G21733,G21917,G21918);
  nand GNAME21734(G21734,G21778,G21770);
  and GNAME21735(G21735,G21779,G21769);
  and GNAME21736(G21736,G21919,G21920);
  nor GNAME21737(G21737,G21925,G21659);
  and GNAME21738(G21738,G21750,G21749);
  not GNAME21739(G21739,G21638);
  not GNAME21740(G21740,G21651);
  not GNAME21741(G21741,G21653);
  not GNAME21742(G21742,G21655);
  not GNAME21743(G21743,G21657);
  not GNAME21744(G21744,G21716);
  nand GNAME21745(G21745,G21766,G21648,G21765);
  nand GNAME21746(G21746,G21773,G21644,G21772);
  nand GNAME21747(G21747,G21767,G8182);
  nand GNAME21748(G21748,G21810,G8189);
  nand GNAME21749(G21749,G21813,G8190);
  nand GNAME21750(G21750,G21636,G21811,G21812);
  nand GNAME21751(G21751,G21750,G8788);
  nand GNAME21752(G21752,G21635,G21808,G21809);
  and GNAME21753(G21753,G21748,G21791);
  not GNAME21754(G21754,G21637);
  not GNAME21755(G21755,G21639);
  not GNAME21756(G21756,G21640);
  nand GNAME21757(G21757,G21820,G8188);
  nand GNAME21758(G21758,G21642,G21800,G21801);
  nand GNAME21759(G21759,G21758,G21641);
  nand GNAME21760(G21760,G21823,G8187);
  nand GNAME21761(G21761,G21643,G21821,G21822);
  or GNAME21762(G21762,G21661,G21755);
  nand GNAME21763(G21763,G21762,G21662);
  nand GNAME21764(G21764,G21858,G8181);
  or GNAME21765(G21765,G8166,G21634);
  nand GNAME21766(G21766,G21634,G8166);
  nand GNAME21767(G21767,G21766,G21765);
  nand GNAME21768(G21768,G21855,G8183);
  nand GNAME21769(G21769,G21852,G8184);
  nand GNAME21770(G21770,G21849,G8185);
  nand GNAME21771(G21771,G21645,G21847,G21848);
  or GNAME21772(G21772,G8170,G21634);
  nand GNAME21773(G21773,G21634,G8170);
  nand GNAME21774(G21774,G21760,G21794);
  nand GNAME21775(G21775,G21772,G21773);
  nand GNAME21776(G21776,G21775,G8186);
  not GNAME21777(G21777,G21737);
  nand GNAME21778(G21778,G21771,G21777);
  nand GNAME21779(G21779,G21646,G21850,G21851);
  nand GNAME21780(G21780,G21734,G21779);
  nand GNAME21781(G21781,G21647,G21853,G21854);
  nand GNAME21782(G21782,G21731,G21781);
  not GNAME21783(G21783,G21730);
  nand GNAME21784(G21784,G21745,G21783);
  nand GNAME21785(G21785,G21649,G21856,G21857);
  nand GNAME21786(G21786,G21727,G21785);
  not GNAME21787(G21787,G21652);
  not GNAME21788(G21788,G21654);
  not GNAME21789(G21789,G21656);
  nand GNAME21790(G21790,G21658,G21671);
  nand GNAME21791(G21791,G21721,G21752);
  nand GNAME21792(G21792,G21665,G21748,G21791);
  nand GNAME21793(G21793,G21746,G21776);
  nand GNAME21794(G21794,G21707,G21761);
  nand GNAME21795(G21795,G21794,G21760,G21793);
  nand GNAME21796(G21796,G21776,G21659);
  not GNAME21797(G21797,G21738);
  nand GNAME21798(G21798,G21745,G21747);
  nand GNAME21799(G21799,G21770,G21771);
  or GNAME21800(G21800,G8172,G21634);
  or GNAME21801(G21801,G8788,G21703);
  or GNAME21802(G21802,G8173,G21634);
  nand GNAME21803(G21803,G21634,G8173);
  or GNAME21804(G21804,G8176,G21634);
  nand GNAME21805(G21805,G21634,G8176);
  or GNAME21806(G21806,G8177,G21634);
  nand GNAME21807(G21807,G21634,G8177);
  or GNAME21808(G21808,G8179,G21634);
  or GNAME21809(G21809,G8788,G21704);
  nand GNAME21810(G21810,G21808,G21809);
  or GNAME21811(G21811,G8180,G21634);
  or GNAME21812(G21812,G8788,G21705);
  nand GNAME21813(G21813,G21811,G21812);
  or GNAME21814(G21814,G8178,G21634);
  nand GNAME21815(G21815,G21634,G8178);
  or GNAME21816(G21816,G8175,G21634);
  nand GNAME21817(G21817,G21634,G8175);
  or GNAME21818(G21818,G8174,G21634);
  nand GNAME21819(G21819,G21634,G8174);
  nand GNAME21820(G21820,G21800,G21801);
  or GNAME21821(G21821,G8171,G21634);
  or GNAME21822(G21822,G8788,G21706);
  nand GNAME21823(G21823,G21821,G21822);
  or GNAME21824(G21824,G21708,G21707);
  nand GNAME21825(G21825,G21707,G21708);
  nand GNAME21826(G21826,G21710,G21641);
  or GNAME21827(G21827,G21641,G21710);
  nand GNAME21828(G21828,G21640,G21660);
  or GNAME21829(G21829,G21640,G21660);
  nand GNAME21830(G21830,G21639,G21661);
  or GNAME21831(G21831,G21639,G21661);
  nand GNAME21832(G21832,G21638,G21663);
  or GNAME21833(G21833,G21638,G21663);
  nand GNAME21834(G21834,G21637,G21664);
  or GNAME21835(G21835,G21637,G21664);
  or GNAME21836(G21836,G8149,G21634);
  or GNAME21837(G21837,G8788,G21711);
  nand GNAME21838(G21838,G21836,G21837);
  or GNAME21839(G21839,G8150,G21634);
  nand GNAME21840(G21840,G21634,G8150);
  or GNAME21841(G21841,G8155,G21634);
  nand GNAME21842(G21842,G21634,G8155);
  or GNAME21843(G21843,G8158,G21634);
  nand GNAME21844(G21844,G21634,G8158);
  or GNAME21845(G21845,G8161,G21634);
  nand GNAME21846(G21846,G21634,G8161);
  or GNAME21847(G21847,G8169,G21634);
  or GNAME21848(G21848,G8788,G21712);
  nand GNAME21849(G21849,G21847,G21848);
  or GNAME21850(G21850,G8168,G21634);
  or GNAME21851(G21851,G8788,G21713);
  nand GNAME21852(G21852,G21850,G21851);
  or GNAME21853(G21853,G8167,G21634);
  or GNAME21854(G21854,G8788,G21714);
  nand GNAME21855(G21855,G21853,G21854);
  or GNAME21856(G21856,G8165,G21634);
  or GNAME21857(G21857,G8788,G21715);
  nand GNAME21858(G21858,G21856,G21857);
  or GNAME21859(G21859,G8164,G21634);
  nand GNAME21860(G21860,G21634,G8164);
  or GNAME21861(G21861,G8163,G21634);
  nand GNAME21862(G21862,G21634,G8163);
  or GNAME21863(G21863,G8162,G21634);
  nand GNAME21864(G21864,G21634,G8162);
  or GNAME21865(G21865,G8160,G21634);
  nand GNAME21866(G21866,G21634,G8160);
  or GNAME21867(G21867,G8159,G21634);
  nand GNAME21868(G21868,G21634,G8159);
  or GNAME21869(G21869,G8157,G21634);
  nand GNAME21870(G21870,G21634,G8157);
  or GNAME21871(G21871,G8156,G21634);
  nand GNAME21872(G21872,G21634,G8156);
  or GNAME21873(G21873,G8154,G21634);
  nand GNAME21874(G21874,G21634,G8154);
  or GNAME21875(G21875,G8153,G21634);
  nand GNAME21876(G21876,G21634,G8153);
  or GNAME21877(G21877,G8151,G21634);
  nand GNAME21878(G21878,G21634,G8151);
  or GNAME21879(G21879,G8152,G21634);
  nand GNAME21880(G21880,G21634,G8152);
  nand GNAME21881(G21881,G21744,G21838);
  nand GNAME21882(G21882,G21716,G21836,G21837);
  nand GNAME21883(G21883,G21672,G21717);
  or GNAME21884(G21884,G21717,G21672);
  nand GNAME21885(G21885,G21657,G21673);
  or GNAME21886(G21886,G21657,G21673);
  nand GNAME21887(G21887,G21675,G21718);
  or GNAME21888(G21888,G21718,G21675);
  nand GNAME21889(G21889,G21656,G21674);
  or GNAME21890(G21890,G21656,G21674);
  nand GNAME21891(G21891,G21655,G21676);
  or GNAME21892(G21892,G21655,G21676);
  nand GNAME21893(G21893,G21678,G21719);
  or GNAME21894(G21894,G21719,G21678);
  nand GNAME21895(G21895,G21654,G21677);
  or GNAME21896(G21896,G21654,G21677);
  nand GNAME21897(G21897,G21653,G21679);
  or GNAME21898(G21898,G21653,G21679);
  nand GNAME21899(G21899,G21681,G21720);
  or GNAME21900(G21900,G21720,G21681);
  nand GNAME21901(G21901,G21652,G21680);
  or GNAME21902(G21902,G21652,G21680);
  or GNAME21903(G21903,G21722,G21721);
  nand GNAME21904(G21904,G21721,G21722);
  nand GNAME21905(G21905,G21651,G21682);
  or GNAME21906(G21906,G21651,G21682);
  nand GNAME21907(G21907,G21684,G21724);
  or GNAME21908(G21908,G21724,G21684);
  nand GNAME21909(G21909,G21650,G21683);
  or GNAME21910(G21910,G21650,G21683);
  nand GNAME21911(G21911,G21685,G21725);
  or GNAME21912(G21912,G21725,G21685);
  or GNAME21913(G21913,G21728,G21727);
  nand GNAME21914(G21914,G21727,G21728);
  nand GNAME21915(G21915,G21783,G21798);
  nand GNAME21916(G21916,G21730,G21745,G21747);
  or GNAME21917(G21917,G21732,G21731);
  nand GNAME21918(G21918,G21731,G21732);
  or GNAME21919(G21919,G21735,G21734);
  nand GNAME21920(G21920,G21734,G21735);
  nand GNAME21921(G21921,G21777,G21799);
  nand GNAME21922(G21922,G21737,G21770,G21771);
  or GNAME21923(G21923,G21738,G21634);
  or GNAME21924(G21924,G8788,G21797);
  not GNAME21925(G21925,G21776);
  not GNAME21926(G21926,G8118);
  not GNAME21927(G21927,G8123);
  not GNAME21928(G21928,G8117);
  not GNAME21929(G21929,G8119);
  not GNAME21930(G21930,G8124);
  not GNAME21931(G21931,G8121);
  not GNAME21932(G21932,G8122);
  not GNAME21933(G21933,G8120);
  and GNAME21934(G21934,G22101,G22125);
  and GNAME21935(G21935,G22055,G22123);
  and GNAME21936(G21936,G22120,G22121);
  and GNAME21937(G21937,G22056,G22117);
  and GNAME21938(G21938,G22090,G22091);
  not GNAME21939(G21939,G8833);
  not GNAME21940(G21940,G8232);
  not GNAME21941(G21941,G8233);
  not GNAME21942(G21942,G8236);
  not GNAME21943(G21943,G8237);
  not GNAME21944(G21944,G8238);
  not GNAME21945(G21945,G8235);
  not GNAME21946(G21946,G8234);
  not GNAME21947(G21947,G8231);
  nor GNAME21948(G21948,G22005,G21970);
  and GNAME21949(G21949,G22083,G22057);
  nor GNAME21950(G21950,G22154,G21969,G21983);
  nor GNAME21951(G21951,G21982,G22101);
  nor GNAME21952(G21952,G21981,G22054);
  nor GNAME21953(G21953,G22059,G21979,G21980);
  nor GNAME21954(G21954,G21978,G22055);
  not GNAME21955(G21955,G8230);
  not GNAME21956(G21956,G8229);
  not GNAME21957(G21957,G8228);
  not GNAME21958(G21958,G8227);
  not GNAME21959(G21959,G8226);
  not GNAME21960(G21960,G8225);
  not GNAME21961(G21961,G8224);
  not GNAME21962(G21962,G8223);
  nor GNAME21963(G21963,G22026,G21984);
  nor GNAME21964(G21964,G22229,G21976,G21977);
  and GNAME21965(G21965,G22260,G21964);
  nor GNAME21966(G21966,G21974,G22261);
  nand GNAME21967(G21967,G22262,G21966);
  and GNAME21968(G21968,G22075,G22058);
  and GNAME21969(G21969,G22149,G22150);
  and GNAME21970(G21970,G22147,G22148);
  nand GNAME21971(G21971,G22151,G22152);
  and GNAME21972(G21972,G22166,G22167);
  and GNAME21973(G21973,G22168,G22169);
  and GNAME21974(G21974,G22170,G22171);
  and GNAME21975(G21975,G22172,G22173);
  and GNAME21976(G21976,G22212,G22213);
  and GNAME21977(G21977,G22214,G22215);
  and GNAME21978(G21978,G22176,G22177);
  and GNAME21979(G21979,G22184,G22185);
  and GNAME21980(G21980,G22186,G22187);
  and GNAME21981(G21981,G22178,G22179);
  and GNAME21982(G21982,G22180,G22181);
  and GNAME21983(G21983,G22182,G22183);
  and GNAME21984(G21984,G22210,G22211);
  nand GNAME21985(G21985,G22218,G22219);
  nand GNAME21986(G21986,G22220,G22221);
  nand GNAME21987(G21987,G22222,G22223);
  nand GNAME21988(G21988,G22224,G22225);
  nand GNAME21989(G21989,G22226,G22227);
  nand GNAME21990(G21990,G22246,G22247);
  nand GNAME21991(G21991,G22248,G22249);
  nand GNAME21992(G21992,G22250,G22251);
  nand GNAME21993(G21993,G22252,G22253);
  nand GNAME21994(G21994,G22254,G22255);
  nand GNAME21995(G21995,G22256,G22257);
  nand GNAME21996(G21996,G22155,G22156);
  nand GNAME21997(G21997,G22161,G22162);
  nand GNAME21998(G21998,G22216,G22217);
  not GNAME21999(G21999,G8215);
  not GNAME22000(G22000,G8217);
  not GNAME22001(G22001,G8219);
  not GNAME22002(G22002,G8221);
  not GNAME22003(G22003,G8222);
  not GNAME22004(G22004,G8218);
  and GNAME22005(G22005,G22087,G22060);
  and GNAME22006(G22006,G22153,G22154);
  nor GNAME22007(G22007,G22259,G21949);
  nand GNAME22008(G22008,G22081,G22065);
  and GNAME22009(G22009,G22082,G22062);
  and GNAME22010(G22010,G22157,G22158);
  nand GNAME22011(G22011,G22079,G22066);
  and GNAME22012(G22012,G22080,G22065);
  and GNAME22013(G22013,G22159,G22160);
  nor GNAME22014(G22014,G22258,G21968);
  not GNAME22015(G22015,G8191);
  not GNAME22016(G22016,G8206);
  not GNAME22017(G22017,G8205);
  not GNAME22018(G22018,G8204);
  not GNAME22019(G22019,G8203);
  not GNAME22020(G22020,G8202);
  not GNAME22021(G22021,G8201);
  not GNAME22022(G22022,G8200);
  not GNAME22023(G22023,G8199);
  nor GNAME22024(G22024,G21972,G21967);
  nor GNAME22025(G22025,G21977,G22229);
  and GNAME22026(G22026,G22116,G22092);
  and GNAME22027(G22027,G22228,G22229);
  nand GNAME22028(G22028,G22114,G22093);
  and GNAME22029(G22029,G22115,G22092);
  and GNAME22030(G22030,G22230,G22231);
  nand GNAME22031(G22031,G22112,G22094);
  and GNAME22032(G22032,G22113,G22093);
  and GNAME22033(G22033,G22232,G22233);
  nand GNAME22034(G22034,G22110,G22095);
  and GNAME22035(G22035,G22111,G22094);
  and GNAME22036(G22036,G22234,G22235);
  nand GNAME22037(G22037,G22108,G22096);
  and GNAME22038(G22038,G22109,G22095);
  and GNAME22039(G22039,G22236,G22237);
  nand GNAME22040(G22040,G22073,G22071);
  and GNAME22041(G22041,G22074,G22068);
  and GNAME22042(G22042,G22238,G22239);
  nand GNAME22043(G22043,G22106,G22097);
  and GNAME22044(G22044,G22107,G22096);
  and GNAME22045(G22045,G22240,G22241);
  nand GNAME22046(G22046,G22104,G22098);
  and GNAME22047(G22047,G22105,G22097);
  and GNAME22048(G22048,G22242,G22243);
  nand GNAME22049(G22049,G22102,G22099);
  and GNAME22050(G22050,G22103,G22098);
  and GNAME22051(G22051,G22244,G22245);
  nand GNAME22052(G22052,G22100,G22099);
  and GNAME22053(G22053,G22072,G22071);
  not GNAME22054(G22054,G21951);
  not GNAME22055(G22055,G21953);
  not GNAME22056(G22056,G22024);
  nand GNAME22057(G22057,G22064,G21940,G22063);
  nand GNAME22058(G22058,G22070,G21942,G22069);
  not GNAME22059(G22059,G21952);
  nand GNAME22060(G22060,G22146,G8231);
  nand GNAME22061(G22061,G21947,G22129,G22130);
  nand GNAME22062(G22062,G22133,G8233);
  or GNAME22063(G22063,G8216,G21939);
  nand GNAME22064(G22064,G21939,G8216);
  nand GNAME22065(G22065,G22145,G8234);
  nand GNAME22066(G22066,G22142,G8235);
  nand GNAME22067(G22067,G21945,G22134,G22135);
  nand GNAME22068(G22068,G22138,G8237);
  or GNAME22069(G22069,G8220,G21939);
  nand GNAME22070(G22070,G21939,G8220);
  nand GNAME22071(G22071,G22141,G8238);
  nand GNAME22072(G22072,G21944,G22139,G22140);
  nand GNAME22073(G22073,G22072,G8833);
  nand GNAME22074(G22074,G21943,G22136,G22137);
  nand GNAME22075(G22075,G22068,G22118);
  nand GNAME22076(G22076,G22069,G22070);
  nand GNAME22077(G22077,G22076,G8236);
  not GNAME22078(G22078,G22014);
  nand GNAME22079(G22079,G22067,G22078);
  nand GNAME22080(G22080,G21946,G22143,G22144);
  nand GNAME22081(G22081,G22011,G22080);
  nand GNAME22082(G22082,G21941,G22131,G22132);
  nand GNAME22083(G22083,G22062,G22088);
  nand GNAME22084(G22084,G22063,G22064);
  nand GNAME22085(G22085,G22084,G8232);
  not GNAME22086(G22086,G22007);
  nand GNAME22087(G22087,G22061,G22086);
  nand GNAME22088(G22088,G22008,G22082);
  nand GNAME22089(G22089,G22057,G22085);
  nand GNAME22090(G22090,G22089,G22062,G22088);
  nand GNAME22091(G22091,G22085,G21949);
  nand GNAME22092(G22092,G22209,G8223);
  nand GNAME22093(G22093,G22206,G8224);
  nand GNAME22094(G22094,G22203,G8225);
  nand GNAME22095(G22095,G22200,G8226);
  nand GNAME22096(G22096,G22197,G8227);
  nand GNAME22097(G22097,G22194,G8228);
  nand GNAME22098(G22098,G22191,G8229);
  nand GNAME22099(G22099,G22188,G8230);
  nand GNAME22100(G22100,G21955,G22174,G22175);
  not GNAME22101(G22101,G21950);
  nand GNAME22102(G22102,G22100,G21954);
  nand GNAME22103(G22103,G21956,G22189,G22190);
  nand GNAME22104(G22104,G22049,G22103);
  nand GNAME22105(G22105,G21957,G22192,G22193);
  nand GNAME22106(G22106,G22046,G22105);
  nand GNAME22107(G22107,G21958,G22195,G22196);
  nand GNAME22108(G22108,G22043,G22107);
  nand GNAME22109(G22109,G21959,G22198,G22199);
  nand GNAME22110(G22110,G22037,G22109);
  nand GNAME22111(G22111,G21960,G22201,G22202);
  nand GNAME22112(G22112,G22034,G22111);
  nand GNAME22113(G22113,G21961,G22204,G22205);
  nand GNAME22114(G22114,G22031,G22113);
  nand GNAME22115(G22115,G21962,G22207,G22208);
  nand GNAME22116(G22116,G22028,G22115);
  nand GNAME22117(G22117,G21967,G21972);
  nand GNAME22118(G22118,G22040,G22074);
  nand GNAME22119(G22119,G22058,G22077);
  nand GNAME22120(G22120,G22119,G22068,G22118);
  nand GNAME22121(G22121,G22077,G21968);
  or GNAME22122(G22122,G21979,G22059);
  nand GNAME22123(G22123,G22122,G21980);
  or GNAME22124(G22124,G21969,G22154);
  nand GNAME22125(G22125,G22124,G21983);
  not GNAME22126(G22126,G22053);
  nand GNAME22127(G22127,G22060,G22061);
  nand GNAME22128(G22128,G22066,G22067);
  or GNAME22129(G22129,G8215,G21939);
  or GNAME22130(G22130,G8833,G21999);
  or GNAME22131(G22131,G8217,G21939);
  or GNAME22132(G22132,G8833,G22000);
  nand GNAME22133(G22133,G22131,G22132);
  or GNAME22134(G22134,G8219,G21939);
  or GNAME22135(G22135,G8833,G22001);
  or GNAME22136(G22136,G8221,G21939);
  or GNAME22137(G22137,G8833,G22002);
  nand GNAME22138(G22138,G22136,G22137);
  or GNAME22139(G22139,G8222,G21939);
  or GNAME22140(G22140,G8833,G22003);
  nand GNAME22141(G22141,G22139,G22140);
  nand GNAME22142(G22142,G22134,G22135);
  or GNAME22143(G22143,G8218,G21939);
  or GNAME22144(G22144,G8833,G22004);
  nand GNAME22145(G22145,G22143,G22144);
  nand GNAME22146(G22146,G22129,G22130);
  or GNAME22147(G22147,G8214,G21939);
  nand GNAME22148(G22148,G21939,G8214);
  or GNAME22149(G22149,G8213,G21939);
  nand GNAME22150(G22150,G21939,G8213);
  nand GNAME22151(G22151,G21948,G21969);
  or GNAME22152(G22152,G21948,G21969);
  nand GNAME22153(G22153,G21970,G22005);
  or GNAME22154(G22154,G22005,G21970);
  nand GNAME22155(G22155,G22086,G22127);
  nand GNAME22156(G22156,G22007,G22060,G22061);
  or GNAME22157(G22157,G22009,G22008);
  nand GNAME22158(G22158,G22008,G22009);
  or GNAME22159(G22159,G22012,G22011);
  nand GNAME22160(G22160,G22011,G22012);
  nand GNAME22161(G22161,G22078,G22128);
  nand GNAME22162(G22162,G22014,G22066,G22067);
  or GNAME22163(G22163,G8191,G21939);
  or GNAME22164(G22164,G8833,G22015);
  nand GNAME22165(G22165,G22163,G22164);
  or GNAME22166(G22166,G8192,G21939);
  nand GNAME22167(G22167,G21939,G8192);
  or GNAME22168(G22168,G8193,G21939);
  nand GNAME22169(G22169,G21939,G8193);
  or GNAME22170(G22170,G8194,G21939);
  nand GNAME22171(G22171,G21939,G8194);
  or GNAME22172(G22172,G8195,G21939);
  nand GNAME22173(G22173,G21939,G8195);
  or GNAME22174(G22174,G8206,G21939);
  or GNAME22175(G22175,G8833,G22016);
  or GNAME22176(G22176,G8207,G21939);
  nand GNAME22177(G22177,G21939,G8207);
  or GNAME22178(G22178,G8210,G21939);
  nand GNAME22179(G22179,G21939,G8210);
  or GNAME22180(G22180,G8211,G21939);
  nand GNAME22181(G22181,G21939,G8211);
  or GNAME22182(G22182,G8212,G21939);
  nand GNAME22183(G22183,G21939,G8212);
  or GNAME22184(G22184,G8209,G21939);
  nand GNAME22185(G22185,G21939,G8209);
  or GNAME22186(G22186,G8208,G21939);
  nand GNAME22187(G22187,G21939,G8208);
  nand GNAME22188(G22188,G22174,G22175);
  or GNAME22189(G22189,G8205,G21939);
  or GNAME22190(G22190,G8833,G22017);
  nand GNAME22191(G22191,G22189,G22190);
  or GNAME22192(G22192,G8204,G21939);
  or GNAME22193(G22193,G8833,G22018);
  nand GNAME22194(G22194,G22192,G22193);
  or GNAME22195(G22195,G8203,G21939);
  or GNAME22196(G22196,G8833,G22019);
  nand GNAME22197(G22197,G22195,G22196);
  or GNAME22198(G22198,G8202,G21939);
  or GNAME22199(G22199,G8833,G22020);
  nand GNAME22200(G22200,G22198,G22199);
  or GNAME22201(G22201,G8201,G21939);
  or GNAME22202(G22202,G8833,G22021);
  nand GNAME22203(G22203,G22201,G22202);
  or GNAME22204(G22204,G8200,G21939);
  or GNAME22205(G22205,G8833,G22022);
  nand GNAME22206(G22206,G22204,G22205);
  or GNAME22207(G22207,G8199,G21939);
  or GNAME22208(G22208,G8833,G22023);
  nand GNAME22209(G22209,G22207,G22208);
  or GNAME22210(G22210,G8198,G21939);
  nand GNAME22211(G22211,G21939,G8198);
  or GNAME22212(G22212,G8196,G21939);
  nand GNAME22213(G22213,G21939,G8196);
  or GNAME22214(G22214,G8197,G21939);
  nand GNAME22215(G22215,G21939,G8197);
  nand GNAME22216(G22216,G22056,G22165);
  nand GNAME22217(G22217,G22024,G22163,G22164);
  nand GNAME22218(G22218,G21966,G21973);
  or GNAME22219(G22219,G21966,G21973);
  nand GNAME22220(G22220,G21965,G21974);
  or GNAME22221(G22221,G21965,G21974);
  nand GNAME22222(G22222,G21964,G21975);
  or GNAME22223(G22223,G21964,G21975);
  nand GNAME22224(G22224,G21976,G22025);
  or GNAME22225(G22225,G22025,G21976);
  nand GNAME22226(G22226,G21963,G21977);
  or GNAME22227(G22227,G21963,G21977);
  nand GNAME22228(G22228,G21984,G22026);
  or GNAME22229(G22229,G22026,G21984);
  or GNAME22230(G22230,G22029,G22028);
  nand GNAME22231(G22231,G22028,G22029);
  or GNAME22232(G22232,G22032,G22031);
  nand GNAME22233(G22233,G22031,G22032);
  or GNAME22234(G22234,G22035,G22034);
  nand GNAME22235(G22235,G22034,G22035);
  or GNAME22236(G22236,G22038,G22037);
  nand GNAME22237(G22237,G22037,G22038);
  or GNAME22238(G22238,G22041,G22040);
  nand GNAME22239(G22239,G22040,G22041);
  or GNAME22240(G22240,G22044,G22043);
  nand GNAME22241(G22241,G22043,G22044);
  or GNAME22242(G22242,G22047,G22046);
  nand GNAME22243(G22243,G22046,G22047);
  or GNAME22244(G22244,G22050,G22049);
  nand GNAME22245(G22245,G22049,G22050);
  nand GNAME22246(G22246,G22052,G21954);
  or GNAME22247(G22247,G21954,G22052);
  nand GNAME22248(G22248,G21953,G21978);
  or GNAME22249(G22249,G21953,G21978);
  nand GNAME22250(G22250,G21952,G21979);
  or GNAME22251(G22251,G21952,G21979);
  nand GNAME22252(G22252,G21951,G21981);
  or GNAME22253(G22253,G21951,G21981);
  nand GNAME22254(G22254,G21950,G21982);
  or GNAME22255(G22255,G21950,G21982);
  or GNAME22256(G22256,G22053,G21939);
  or GNAME22257(G22257,G8833,G22126);
  not GNAME22258(G22258,G22077);
  not GNAME22259(G22259,G22085);
  not GNAME22260(G22260,G21975);
  not GNAME22261(G22261,G21965);
  not GNAME22262(G22262,G21973);
  nor GNAME22263(G22263,G22266,G22294);
  and GNAME22264(G22264,G22273,G22271,G22272);
  and GNAME22265(G22265,G22268,G22310);
  nor GNAME22266(G22266,G22265,G22264,G22309,G22308);
  not GNAME22267(G22267,G22307);
  not GNAME22268(G22268,G9849);
  not GNAME22269(G22269,G22295);
  or GNAME22270(G22270,G9781,G22267);
  nand GNAME22271(G22271,G9782,G22269,G22270);
  or GNAME22272(G22272,G22310,G22268);
  nand GNAME22273(G22273,G22267,G9781);
  or GNAME22274(G22274,G9277,G22275);
  nor GNAME22275(G22275,G23086,G23087);
  and GNAME22276(G22276,G22292,G22293);
  not GNAME22277(G22277,G9280);
  not GNAME22278(G22278,G59564);
  not GNAME22279(G22279,G9278);
  not GNAME22280(G22280,G9277);
  not GNAME22281(G22281,G9281);
  or GNAME22282(G22282,G59565,G22277);
  nand GNAME22283(G22283,G59566,G22281,G22282);
  or GNAME22284(G22284,G9279,G22278);
  nand GNAME22285(G22285,G22277,G59565);
  nand GNAME22286(G22286,G22285,G22283,G22284);
  or GNAME22287(G22287,G59563,G22279);
  nand GNAME22288(G22288,G22278,G9279);
  nand GNAME22289(G22289,G22288,G22286,G22287);
  nand GNAME22290(G22290,G22280,G59562);
  nand GNAME22291(G22291,G22279,G59563);
  nand GNAME22292(G22292,G22291,G22289,G22290);
  or GNAME22293(G22293,G59562,G22280);
  nand GNAME22294(G22294,G22326,G22327);
  nand GNAME22295(G22295,G22328,G22314);
  not GNAME22296(G22296,G59561);
  not GNAME22297(G22297,G59560);
  not GNAME22298(G22298,G59565);
  and GNAME22299(G22299,G22315,G22345);
  not GNAME22300(G22300,G59559);
  not GNAME22301(G22301,G59564);
  and GNAME22302(G22302,G22318,G22319);
  not GNAME22303(G22303,G59558);
  not GNAME22304(G22304,G59563);
  and GNAME22305(G22305,G22322,G22323);
  not GNAME22306(G22306,G59557);
  nand GNAME22307(G22307,G22346,G22347);
  nand GNAME22308(G22308,G22332,G22333);
  nand GNAME22309(G22309,G22337,G22338);
  nand GNAME22310(G22310,G22342,G22343);
  and GNAME22311(G22311,G22344,G22345);
  not GNAME22312(G22312,G59562);
  nor GNAME22313(G22313,G59566,G22296);
  not GNAME22314(G22314,G22313);
  nand GNAME22315(G22315,G22314,G22344);
  not GNAME22316(G22316,G22299);
  or GNAME22317(G22317,G22316,G22300);
  nand GNAME22318(G22318,G22317,G59564);
  or GNAME22319(G22319,G59559,G22299);
  not GNAME22320(G22320,G22302);
  or GNAME22321(G22321,G22320,G22303);
  nand GNAME22322(G22322,G22321,G59563);
  or GNAME22323(G22323,G59558,G22302);
  not GNAME22324(G22324,G22305);
  or GNAME22325(G22325,G22305,G59557);
  nand GNAME22326(G22326,G22312,G22325);
  or GNAME22327(G22327,G22324,G22306);
  nand GNAME22328(G22328,G22296,G59566);
  or GNAME22329(G22329,G59557,G22312);
  or GNAME22330(G22330,G59562,G22306);
  nand GNAME22331(G22331,G22329,G22330);
  nand GNAME22332(G22332,G22324,G22331);
  nand GNAME22333(G22333,G22305,G22329,G22330);
  or GNAME22334(G22334,G59558,G22304);
  or GNAME22335(G22335,G59563,G22303);
  nand GNAME22336(G22336,G22334,G22335);
  nand GNAME22337(G22337,G22320,G22336);
  nand GNAME22338(G22338,G22302,G22334,G22335);
  or GNAME22339(G22339,G59559,G22301);
  or GNAME22340(G22340,G59564,G22300);
  nand GNAME22341(G22341,G22339,G22340);
  nand GNAME22342(G22342,G22316,G22341);
  nand GNAME22343(G22343,G22299,G22339,G22340);
  or GNAME22344(G22344,G59565,G22297);
  or GNAME22345(G22345,G59560,G22298);
  nand GNAME22346(G22346,G22311,G22313);
  or GNAME22347(G22347,G22313,G22311);
  and GNAME22348(G22348,G22590,G22591);
  and GNAME22349(G22349,G22585,G22586);
  and GNAME22350(G22350,G22579,G22580);
  and GNAME22351(G22351,G22506,G22507);
  not GNAME22352(G22352,G9184);
  not GNAME22353(G22353,G8272);
  not GNAME22354(G22354,G8273);
  not GNAME22355(G22355,G8276);
  not GNAME22356(G22356,G8277);
  not GNAME22357(G22357,G8278);
  not GNAME22358(G22358,G8275);
  not GNAME22359(G22359,G8274);
  not GNAME22360(G22360,G8271);
  and GNAME22361(G22361,G22500,G22473);
  not GNAME22362(G22362,G8270);
  and GNAME22363(G22363,G22496,G22471);
  or GNAME22364(G22364,G22508,G22439);
  not GNAME22365(G22365,G8267);
  and GNAME22366(G22366,G22511,G22512);
  not GNAME22367(G22367,G8266);
  not GNAME22368(G22368,G8265);
  nand GNAME22369(G22369,G22514,G22515);
  nand GNAME22370(G22370,G22518,G22519);
  not GNAME22371(G22371,G8264);
  and GNAME22372(G22372,G22522,G22523);
  not GNAME22373(G22373,G8263);
  and GNAME22374(G22374,G22525,G22526);
  not GNAME22375(G22375,G8262);
  and GNAME22376(G22376,G22528,G22529);
  not GNAME22377(G22377,G8261);
  and GNAME22378(G22378,G22531,G22532);
  not GNAME22379(G22379,G8260);
  and GNAME22380(G22380,G22534,G22535);
  not GNAME22381(G22381,G8259);
  and GNAME22382(G22382,G22537,G22538);
  not GNAME22383(G22383,G8258);
  and GNAME22384(G22384,G22540,G22541);
  not GNAME22385(G22385,G8257);
  and GNAME22386(G22386,G22543,G22544);
  not GNAME22387(G22387,G8256);
  and GNAME22388(G22388,G22546,G22547);
  not GNAME22389(G22389,G8255);
  and GNAME22390(G22390,G22549,G22550);
  not GNAME22391(G22391,G8254);
  and GNAME22392(G22392,G22552,G22553);
  not GNAME22393(G22393,G8253);
  and GNAME22394(G22394,G22555,G22556);
  not GNAME22395(G22395,G8252);
  and GNAME22396(G22396,G22558,G22559);
  not GNAME22397(G22397,G8251);
  and GNAME22398(G22398,G22561,G22562);
  not GNAME22399(G22399,G8250);
  not GNAME22400(G22400,G8249);
  nand GNAME22401(G22401,G22564,G22565);
  nand GNAME22402(G22402,G22568,G22569);
  not GNAME22403(G22403,G8248);
  not GNAME22404(G22404,G8247);
  and GNAME22405(G22405,G22488,G22472);
  nand GNAME22406(G22406,G9184,G8268);
  nand GNAME22407(G22407,G22582,G22583);
  nand GNAME22408(G22408,G22715,G22716);
  nand GNAME22409(G22409,G22622,G22623);
  nand GNAME22410(G22410,G22628,G22629);
  nand GNAME22411(G22411,G22630,G22631);
  nand GNAME22412(G22412,G22635,G22636);
  nand GNAME22413(G22413,G22702,G22703);
  and GNAME22414(G22414,G22614,G22615);
  and GNAME22415(G22415,G22618,G22619);
  and GNAME22416(G22416,G22637,G22638);
  and GNAME22417(G22417,G22641,G22642);
  and GNAME22418(G22418,G22645,G22646);
  and GNAME22419(G22419,G22649,G22650);
  and GNAME22420(G22420,G22653,G22654);
  and GNAME22421(G22421,G22657,G22658);
  and GNAME22422(G22422,G22661,G22662);
  and GNAME22423(G22423,G22665,G22666);
  and GNAME22424(G22424,G22669,G22670);
  and GNAME22425(G22425,G22673,G22674);
  and GNAME22426(G22426,G22679,G22680);
  and GNAME22427(G22427,G22683,G22684);
  and GNAME22428(G22428,G22687,G22688);
  and GNAME22429(G22429,G22691,G22692);
  and GNAME22430(G22430,G22695,G22696);
  and GNAME22431(G22431,G22704,G22705);
  and GNAME22432(G22432,G22708,G22709);
  not GNAME22433(G22433,G8239);
  not GNAME22434(G22434,G8241);
  not GNAME22435(G22435,G8243);
  not GNAME22436(G22436,G8245);
  not GNAME22437(G22437,G8246);
  not GNAME22438(G22438,G8242);
  and GNAME22439(G22439,G22502,G22503);
  and GNAME22440(G22440,G22616,G22617);
  and GNAME22441(G22441,G22620,G22621);
  or GNAME22442(G22442,G22498,G22363);
  nand GNAME22443(G22443,G22494,G22478);
  and GNAME22444(G22444,G22495,G22475);
  and GNAME22445(G22445,G22624,G22625);
  nand GNAME22446(G22446,G22492,G22479);
  and GNAME22447(G22447,G22493,G22478);
  and GNAME22448(G22448,G22626,G22627);
  or GNAME22449(G22449,G22490,G22405);
  and GNAME22450(G22450,G22639,G22640);
  and GNAME22451(G22451,G22643,G22644);
  and GNAME22452(G22452,G22647,G22648);
  and GNAME22453(G22453,G22651,G22652);
  and GNAME22454(G22454,G22655,G22656);
  and GNAME22455(G22455,G22659,G22660);
  and GNAME22456(G22456,G22663,G22664);
  and GNAME22457(G22457,G22667,G22668);
  and GNAME22458(G22458,G22671,G22672);
  and GNAME22459(G22459,G22675,G22676);
  nand GNAME22460(G22460,G22486,G22484);
  and GNAME22461(G22461,G22487,G22481);
  and GNAME22462(G22462,G22677,G22678);
  and GNAME22463(G22463,G22681,G22682);
  and GNAME22464(G22464,G22685,G22686);
  and GNAME22465(G22465,G22689,G22690);
  and GNAME22466(G22466,G22693,G22694);
  and GNAME22467(G22467,G22697,G22698);
  and GNAME22468(G22468,G22706,G22707);
  and GNAME22469(G22469,G22710,G22711);
  nand GNAME22470(G22470,G22485,G22484);
  nand GNAME22471(G22471,G22477,G22353,G22476);
  nand GNAME22472(G22472,G22483,G22355,G22482);
  nand GNAME22473(G22473,G22613,G8271);
  nand GNAME22474(G22474,G22360,G22596,G22597);
  nand GNAME22475(G22475,G22600,G8273);
  or GNAME22476(G22476,G8240,G22352);
  nand GNAME22477(G22477,G22352,G8240);
  nand GNAME22478(G22478,G22612,G8274);
  nand GNAME22479(G22479,G22609,G8275);
  nand GNAME22480(G22480,G22358,G22601,G22602);
  nand GNAME22481(G22481,G22605,G8277);
  or GNAME22482(G22482,G8244,G22352);
  nand GNAME22483(G22483,G22352,G8244);
  nand GNAME22484(G22484,G22608,G8278);
  nand GNAME22485(G22485,G22357,G22606,G22607);
  nand GNAME22486(G22486,G22485,G9184);
  nand GNAME22487(G22487,G22356,G22603,G22604);
  nand GNAME22488(G22488,G22481,G22577);
  nand GNAME22489(G22489,G22482,G22483);
  and GNAME22490(G22490,G22489,G8276);
  not GNAME22491(G22491,G22449);
  nand GNAME22492(G22492,G22480,G22449);
  nand GNAME22493(G22493,G22359,G22610,G22611);
  nand GNAME22494(G22494,G22446,G22493);
  nand GNAME22495(G22495,G22354,G22598,G22599);
  nand GNAME22496(G22496,G22475,G22504);
  nand GNAME22497(G22497,G22476,G22477);
  and GNAME22498(G22498,G22497,G8272);
  not GNAME22499(G22499,G22442);
  nand GNAME22500(G22500,G22474,G22442);
  nand GNAME22501(G22501,G22362,G22361);
  nand GNAME22502(G22502,G22501,G9184);
  or GNAME22503(G22503,G22361,G22362);
  nand GNAME22504(G22504,G22443,G22495);
  nand GNAME22505(G22505,G22471,G22718);
  nand GNAME22506(G22506,G22505,G22475,G22504);
  nand GNAME22507(G22507,G22718,G22363);
  nor GNAME22508(G22508,G8269,G9184);
  not GNAME22509(G22509,G22364);
  or GNAME22510(G22510,G8269,G8267,G22509,G22719);
  nand GNAME22511(G22511,G8267,G22509,G8268);
  nand GNAME22512(G22512,G22510,G9184);
  nand GNAME22513(G22513,G22367,G22366);
  nand GNAME22514(G22514,G22513,G9184);
  or GNAME22515(G22515,G22366,G22367);
  not GNAME22516(G22516,G22369);
  nand GNAME22517(G22517,G22369,G8265);
  nand GNAME22518(G22518,G22352,G22517);
  nand GNAME22519(G22519,G22368,G22516);
  not GNAME22520(G22520,G22370);
  nand GNAME22521(G22521,G22370,G22371);
  nand GNAME22522(G22522,G22521,G9184);
  nand GNAME22523(G22523,G22520,G8264);
  nand GNAME22524(G22524,G22373,G22372);
  nand GNAME22525(G22525,G22524,G9184);
  or GNAME22526(G22526,G22372,G22373);
  nand GNAME22527(G22527,G22375,G22374);
  nand GNAME22528(G22528,G22527,G9184);
  or GNAME22529(G22529,G22374,G22375);
  nand GNAME22530(G22530,G22377,G22376);
  nand GNAME22531(G22531,G22530,G9184);
  or GNAME22532(G22532,G22376,G22377);
  nand GNAME22533(G22533,G22379,G22378);
  nand GNAME22534(G22534,G22533,G9184);
  or GNAME22535(G22535,G22378,G22379);
  nand GNAME22536(G22536,G22381,G22380);
  nand GNAME22537(G22537,G22536,G9184);
  or GNAME22538(G22538,G22380,G22381);
  nand GNAME22539(G22539,G22383,G22382);
  nand GNAME22540(G22540,G22539,G9184);
  or GNAME22541(G22541,G22382,G22383);
  nand GNAME22542(G22542,G22385,G22384);
  nand GNAME22543(G22543,G22542,G9184);
  or GNAME22544(G22544,G22384,G22385);
  nand GNAME22545(G22545,G22387,G22386);
  nand GNAME22546(G22546,G22545,G9184);
  or GNAME22547(G22547,G22386,G22387);
  nand GNAME22548(G22548,G22389,G22388);
  nand GNAME22549(G22549,G22548,G9184);
  or GNAME22550(G22550,G22388,G22389);
  nand GNAME22551(G22551,G22391,G22390);
  nand GNAME22552(G22552,G22551,G9184);
  or GNAME22553(G22553,G22390,G22391);
  nand GNAME22554(G22554,G22393,G22392);
  nand GNAME22555(G22555,G22554,G9184);
  or GNAME22556(G22556,G22392,G22393);
  nand GNAME22557(G22557,G22395,G22394);
  nand GNAME22558(G22558,G22557,G9184);
  or GNAME22559(G22559,G22394,G22395);
  nand GNAME22560(G22560,G22397,G22396);
  nand GNAME22561(G22561,G22560,G9184);
  or GNAME22562(G22562,G22396,G22397);
  nand GNAME22563(G22563,G22399,G22398);
  nand GNAME22564(G22564,G22563,G9184);
  or GNAME22565(G22565,G22398,G22399);
  not GNAME22566(G22566,G22401);
  nand GNAME22567(G22567,G22401,G8249);
  nand GNAME22568(G22568,G22352,G22567);
  nand GNAME22569(G22569,G22400,G22566);
  not GNAME22570(G22570,G22402);
  nand GNAME22571(G22571,G22570,G8248);
  nand GNAME22572(G22572,G22352,G22571);
  nand GNAME22573(G22573,G22403,G22402);
  nand GNAME22574(G22574,G8247,G22572,G22573);
  nand GNAME22575(G22575,G22573,G9184);
  nand GNAME22576(G22576,G22571,G22404,G22575);
  nand GNAME22577(G22577,G22460,G22487);
  nand GNAME22578(G22578,G22472,G22717);
  nand GNAME22579(G22579,G22578,G22481,G22577);
  nand GNAME22580(G22580,G22717,G22405);
  nand GNAME22581(G22581,G22509,G8268);
  nand GNAME22582(G22582,G22352,G22581);
  or GNAME22583(G22583,G8269,G22509);
  nand GNAME22584(G22584,G22406,G22407);
  nand GNAME22585(G22585,G22584,G22714);
  nand GNAME22586(G22586,G22712,G22713,G22406,G22407);
  or GNAME22587(G22587,G8269,G22406);
  nand GNAME22588(G22588,G22587,G9184);
  nand GNAME22589(G22589,G22406,G8268);
  nand GNAME22590(G22590,G22589,G22364,G22588);
  or GNAME22591(G22591,G22719,G22407);
  not GNAME22592(G22592,G22470);
  nand GNAME22593(G22593,G22473,G22474);
  nand GNAME22594(G22594,G22479,G22480);
  nand GNAME22595(G22595,G22574,G22576);
  nand GNAME22596(G22596,G22433,G9184);
  nand GNAME22597(G22597,G22352,G8239);
  nand GNAME22598(G22598,G22434,G9184);
  nand GNAME22599(G22599,G22352,G8241);
  nand GNAME22600(G22600,G22598,G22599);
  nand GNAME22601(G22601,G22435,G9184);
  nand GNAME22602(G22602,G22352,G8243);
  nand GNAME22603(G22603,G22436,G9184);
  nand GNAME22604(G22604,G22352,G8245);
  nand GNAME22605(G22605,G22603,G22604);
  nand GNAME22606(G22606,G22437,G9184);
  nand GNAME22607(G22607,G22352,G8246);
  nand GNAME22608(G22608,G22606,G22607);
  nand GNAME22609(G22609,G22601,G22602);
  nand GNAME22610(G22610,G22438,G9184);
  nand GNAME22611(G22611,G22352,G8242);
  nand GNAME22612(G22612,G22610,G22611);
  nand GNAME22613(G22613,G22596,G22597);
  or GNAME22614(G22614,G8269,G22352);
  nand GNAME22615(G22615,G22352,G8269);
  nand GNAME22616(G22616,G22414,G22439);
  or GNAME22617(G22617,G22439,G22414);
  nand GNAME22618(G22618,G22362,G9184);
  nand GNAME22619(G22619,G22352,G8270);
  nand GNAME22620(G22620,G22361,G22415);
  or GNAME22621(G22621,G22361,G22415);
  nand GNAME22622(G22622,G22442,G22593);
  nand GNAME22623(G22623,G22499,G22473,G22474);
  or GNAME22624(G22624,G22444,G22443);
  nand GNAME22625(G22625,G22443,G22444);
  or GNAME22626(G22626,G22447,G22446);
  nand GNAME22627(G22627,G22446,G22447);
  nand GNAME22628(G22628,G22449,G22594);
  nand GNAME22629(G22629,G22491,G22479,G22480);
  nand GNAME22630(G22630,G22595,G9184);
  nand GNAME22631(G22631,G22352,G22574,G22576);
  nand GNAME22632(G22632,G22403,G9184);
  nand GNAME22633(G22633,G22352,G8248);
  nand GNAME22634(G22634,G22632,G22633);
  nand GNAME22635(G22635,G22402,G22634);
  nand GNAME22636(G22636,G22570,G22632,G22633);
  nand GNAME22637(G22637,G22400,G9184);
  nand GNAME22638(G22638,G22352,G8249);
  nand GNAME22639(G22639,G22566,G22416);
  or GNAME22640(G22640,G22566,G22416);
  nand GNAME22641(G22641,G22399,G9184);
  nand GNAME22642(G22642,G22352,G8250);
  nand GNAME22643(G22643,G22398,G22417);
  or GNAME22644(G22644,G22398,G22417);
  nand GNAME22645(G22645,G22397,G9184);
  nand GNAME22646(G22646,G22352,G8251);
  nand GNAME22647(G22647,G22396,G22418);
  or GNAME22648(G22648,G22396,G22418);
  nand GNAME22649(G22649,G22395,G9184);
  nand GNAME22650(G22650,G22352,G8252);
  nand GNAME22651(G22651,G22394,G22419);
  or GNAME22652(G22652,G22394,G22419);
  nand GNAME22653(G22653,G22393,G9184);
  nand GNAME22654(G22654,G22352,G8253);
  nand GNAME22655(G22655,G22392,G22420);
  or GNAME22656(G22656,G22392,G22420);
  nand GNAME22657(G22657,G22391,G9184);
  nand GNAME22658(G22658,G22352,G8254);
  nand GNAME22659(G22659,G22390,G22421);
  or GNAME22660(G22660,G22390,G22421);
  nand GNAME22661(G22661,G22389,G9184);
  nand GNAME22662(G22662,G22352,G8255);
  nand GNAME22663(G22663,G22388,G22422);
  or GNAME22664(G22664,G22388,G22422);
  nand GNAME22665(G22665,G22387,G9184);
  nand GNAME22666(G22666,G22352,G8256);
  nand GNAME22667(G22667,G22386,G22423);
  or GNAME22668(G22668,G22386,G22423);
  nand GNAME22669(G22669,G22385,G9184);
  nand GNAME22670(G22670,G22352,G8257);
  nand GNAME22671(G22671,G22384,G22424);
  or GNAME22672(G22672,G22384,G22424);
  nand GNAME22673(G22673,G22383,G9184);
  nand GNAME22674(G22674,G22352,G8258);
  nand GNAME22675(G22675,G22382,G22425);
  or GNAME22676(G22676,G22382,G22425);
  or GNAME22677(G22677,G22461,G22460);
  nand GNAME22678(G22678,G22460,G22461);
  nand GNAME22679(G22679,G22381,G9184);
  nand GNAME22680(G22680,G22352,G8259);
  nand GNAME22681(G22681,G22380,G22426);
  or GNAME22682(G22682,G22380,G22426);
  nand GNAME22683(G22683,G22379,G9184);
  nand GNAME22684(G22684,G22352,G8260);
  nand GNAME22685(G22685,G22378,G22427);
  or GNAME22686(G22686,G22378,G22427);
  nand GNAME22687(G22687,G22377,G9184);
  nand GNAME22688(G22688,G22352,G8261);
  nand GNAME22689(G22689,G22376,G22428);
  or GNAME22690(G22690,G22376,G22428);
  nand GNAME22691(G22691,G22375,G9184);
  nand GNAME22692(G22692,G22352,G8262);
  nand GNAME22693(G22693,G22374,G22429);
  or GNAME22694(G22694,G22374,G22429);
  nand GNAME22695(G22695,G22373,G9184);
  nand GNAME22696(G22696,G22352,G8263);
  nand GNAME22697(G22697,G22372,G22430);
  or GNAME22698(G22698,G22372,G22430);
  nand GNAME22699(G22699,G22371,G9184);
  nand GNAME22700(G22700,G22352,G8264);
  nand GNAME22701(G22701,G22699,G22700);
  nand GNAME22702(G22702,G22370,G22701);
  nand GNAME22703(G22703,G22520,G22699,G22700);
  nand GNAME22704(G22704,G22368,G9184);
  nand GNAME22705(G22705,G22352,G8265);
  nand GNAME22706(G22706,G22516,G22431);
  or GNAME22707(G22707,G22516,G22431);
  nand GNAME22708(G22708,G22367,G9184);
  nand GNAME22709(G22709,G22352,G8266);
  nand GNAME22710(G22710,G22366,G22432);
  or GNAME22711(G22711,G22366,G22432);
  nand GNAME22712(G22712,G22365,G9184);
  nand GNAME22713(G22713,G22352,G8267);
  nand GNAME22714(G22714,G22712,G22713);
  nand GNAME22715(G22715,G22470,G9184);
  nand GNAME22716(G22716,G22352,G22592);
  not GNAME22717(G22717,G22490);
  not GNAME22718(G22718,G22498);
  not GNAME22719(G22719,G22406);
  and GNAME22720(G22720,G22814,G22815);
  not GNAME22721(G22721,G22006);
  not GNAME22722(G22722,G8131);
  and GNAME22723(G22723,G8132,G22006);
  and GNAME22724(G22724,G22794,G22795);
  not GNAME22725(G22725,G8130);
  and GNAME22726(G22726,G22797,G22798);
  not GNAME22727(G22727,G8129);
  and GNAME22728(G22728,G22800,G22801);
  not GNAME22729(G22729,G8128);
  and GNAME22730(G22730,G22803,G22804);
  not GNAME22731(G22731,G8127);
  not GNAME22732(G22732,G8126);
  and GNAME22733(G22733,G22806,G22807);
  and GNAME22734(G22734,G22810,G22811);
  not GNAME22735(G22735,G21990);
  nor GNAME22736(G22736,G22782,G22735);
  not GNAME22737(G22737,G22048);
  not GNAME22738(G22738,G22051);
  nand GNAME22739(G22739,G22051,G22736,G22048);
  and GNAME22740(G22740,G22045,G22873);
  not GNAME22741(G22741,G22036);
  not GNAME22742(G22742,G22039);
  nand GNAME22743(G22743,G22039,G22740,G22036);
  and GNAME22744(G22744,G22033,G22874);
  not GNAME22745(G22745,G22027);
  not GNAME22746(G22746,G22030);
  not GNAME22747(G22747,G21988);
  nand GNAME22748(G22748,G22030,G22744,G22027);
  nand GNAME22749(G22749,G22791,G21988,G21989);
  and GNAME22750(G22750,G21987,G22875);
  not GNAME22751(G22751,G21986);
  and GNAME22752(G22752,G22750,G21986);
  not GNAME22753(G22753,G21985);
  and GNAME22754(G22754,G22812,G22734);
  nand GNAME22755(G22755,G22818,G22819);
  nand GNAME22756(G22756,G22820,G22821);
  nand GNAME22757(G22757,G22822,G22823);
  nand GNAME22758(G22758,G22824,G22825);
  nand GNAME22759(G22759,G22826,G22827);
  nand GNAME22760(G22760,G22828,G22829);
  nand GNAME22761(G22761,G22830,G22831);
  nand GNAME22762(G22762,G22832,G22833);
  nand GNAME22763(G22763,G22834,G22835);
  nand GNAME22764(G22764,G22836,G22837);
  nand GNAME22765(G22765,G22838,G22839);
  nand GNAME22766(G22766,G22840,G22841);
  nand GNAME22767(G22767,G22842,G22843);
  nand GNAME22768(G22768,G22844,G22845);
  nand GNAME22769(G22769,G22846,G22847);
  nand GNAME22770(G22770,G22848,G22849);
  and GNAME22771(G22771,G22816,G22817);
  and GNAME22772(G22772,G22852,G22853);
  and GNAME22773(G22773,G22856,G22857);
  and GNAME22774(G22774,G22860,G22861);
  and GNAME22775(G22775,G22864,G22865);
  and GNAME22776(G22776,G22868,G22869);
  nand GNAME22777(G22777,G22752,G21985);
  and GNAME22778(G22778,G21989,G22791);
  and GNAME22779(G22779,G22744,G22030);
  and GNAME22780(G22780,G22740,G22039);
  and GNAME22781(G22781,G22736,G22051);
  nor GNAME22782(G22782,G22872,G22754);
  and GNAME22783(G22783,G22850,G22851);
  not GNAME22784(G22784,G21935);
  and GNAME22785(G22785,G22854,G22855);
  and GNAME22786(G22786,G22858,G22859);
  and GNAME22787(G22787,G22862,G22863);
  and GNAME22788(G22788,G22866,G22867);
  and GNAME22789(G22789,G22870,G22871);
  not GNAME22790(G22790,G22782);
  not GNAME22791(G22791,G22748);
  nand GNAME22792(G22792,G21991,G8125);
  or GNAME22793(G22793,G21971,G8131);
  nand GNAME22794(G22794,G22793,G22723);
  nand GNAME22795(G22795,G21971,G8131);
  nand GNAME22796(G22796,G22725,G22724);
  nand GNAME22797(G22797,G22796,G21934);
  or GNAME22798(G22798,G22724,G22725);
  nand GNAME22799(G22799,G22727,G22726);
  nand GNAME22800(G22800,G22799,G21994);
  or GNAME22801(G22801,G22726,G22727);
  nand GNAME22802(G22802,G22729,G22728);
  nand GNAME22803(G22803,G22802,G21993);
  or GNAME22804(G22804,G22728,G22729);
  nand GNAME22805(G22805,G22731,G22730);
  nand GNAME22806(G22806,G22805,G21992);
  or GNAME22807(G22807,G22730,G22731);
  not GNAME22808(G22808,G22733);
  or GNAME22809(G22809,G22733,G22732);
  nand GNAME22810(G22810,G22784,G22809);
  or GNAME22811(G22811,G8126,G22808);
  or GNAME22812(G22812,G8125,G21991);
  and GNAME22813(G22813,G22792,G22812);
  or GNAME22814(G22814,G22813,G22734);
  nand GNAME22815(G22815,G22792,G22754);
  nand GNAME22816(G22816,G22722,G21971);
  or GNAME22817(G22817,G21971,G22722);
  nand GNAME22818(G22818,G22723,G22771);
  or GNAME22819(G22819,G22723,G22771);
  or GNAME22820(G22820,G8132,G22721);
  nand GNAME22821(G22821,G22721,G8132);
  nand GNAME22822(G22822,G22777,G21937);
  or GNAME22823(G22823,G21937,G22777);
  or GNAME22824(G22824,G22752,G22753);
  nand GNAME22825(G22825,G22753,G22752);
  or GNAME22826(G22826,G22750,G22751);
  nand GNAME22827(G22827,G22751,G22750);
  or GNAME22828(G22828,G21987,G22749);
  nand GNAME22829(G22829,G22749,G21987);
  or GNAME22830(G22830,G22778,G22747);
  nand GNAME22831(G22831,G22747,G22778);
  or GNAME22832(G22832,G21989,G22748);
  nand GNAME22833(G22833,G22748,G21989);
  or GNAME22834(G22834,G22779,G22745);
  nand GNAME22835(G22835,G22745,G22779);
  or GNAME22836(G22836,G22744,G22746);
  nand GNAME22837(G22837,G22746,G22744);
  or GNAME22838(G22838,G22033,G22743);
  nand GNAME22839(G22839,G22743,G22033);
  or GNAME22840(G22840,G22780,G22741);
  nand GNAME22841(G22841,G22741,G22780);
  or GNAME22842(G22842,G22740,G22742);
  nand GNAME22843(G22843,G22742,G22740);
  or GNAME22844(G22844,G22045,G22739);
  nand GNAME22845(G22845,G22739,G22045);
  or GNAME22846(G22846,G22781,G22737);
  nand GNAME22847(G22847,G22737,G22781);
  or GNAME22848(G22848,G22736,G22738);
  nand GNAME22849(G22849,G22738,G22736);
  or GNAME22850(G22850,G22782,G22735);
  or GNAME22851(G22851,G21990,G22790);
  or GNAME22852(G22852,G8126,G22784);
  or GNAME22853(G22853,G21935,G22732);
  nand GNAME22854(G22854,G22733,G22772);
  or GNAME22855(G22855,G22733,G22772);
  nand GNAME22856(G22856,G22731,G21992);
  or GNAME22857(G22857,G21992,G22731);
  nand GNAME22858(G22858,G22730,G22773);
  or GNAME22859(G22859,G22730,G22773);
  nand GNAME22860(G22860,G22729,G21993);
  or GNAME22861(G22861,G21993,G22729);
  nand GNAME22862(G22862,G22728,G22774);
  or GNAME22863(G22863,G22728,G22774);
  nand GNAME22864(G22864,G22727,G21994);
  or GNAME22865(G22865,G21994,G22727);
  nand GNAME22866(G22866,G22726,G22775);
  or GNAME22867(G22867,G22726,G22775);
  nand GNAME22868(G22868,G22725,G21934);
  or GNAME22869(G22869,G21934,G22725);
  nand GNAME22870(G22870,G22724,G22776);
  or GNAME22871(G22871,G22724,G22776);
  not GNAME22872(G22872,G22792);
  not GNAME22873(G22873,G22739);
  not GNAME22874(G22874,G22743);
  not GNAME22875(G22875,G22749);
  not GNAME22876(G22876,G9275);
  not GNAME22877(G22877,G9276);
  not GNAME22878(G22878,G8116);
  not GNAME22879(G22879,G9274);
  nor GNAME22880(G22880,G22920,G23006);
  and GNAME22881(G22881,G22973,G23004);
  nor GNAME22882(G22882,G22922,G23003);
  and GNAME22883(G22883,G23081,G23001);
  nand GNAME22884(G22884,G22974,G9866);
  not GNAME22885(G22885,G8301);
  not GNAME22886(G22886,G8302);
  not GNAME22887(G22887,G8299);
  and GNAME22888(G22888,G22975,G8299);
  not GNAME22889(G22889,G8298);
  not GNAME22890(G22890,G8297);
  and GNAME22891(G22891,G8297,G22888,G8298);
  and GNAME22892(G22892,G8296,G22891);
  not GNAME22893(G22893,G8294);
  not GNAME22894(G22894,G8295);
  and GNAME22895(G22895,G8295,G22892,G8294);
  not GNAME22896(G22896,G8293);
  nand GNAME22897(G22897,G22895,G8293);
  not GNAME22898(G22898,G8292);
  not GNAME22899(G22899,G8291);
  and GNAME22900(G22900,G8291,G22976,G8292);
  not GNAME22901(G22901,G8289);
  and GNAME22902(G22902,G8289,G8290,G22900);
  not GNAME22903(G22903,G8287);
  and GNAME22904(G22904,G8287,G8288,G22902);
  not GNAME22905(G22905,G8286);
  and GNAME22906(G22906,G22978,G22979);
  not GNAME22907(G22907,G8309);
  and GNAME22908(G22908,G22981,G22982);
  not GNAME22909(G22909,G8308);
  and GNAME22910(G22910,G22984,G22985);
  not GNAME22911(G22911,G8307);
  and GNAME22912(G22912,G22987,G22988);
  not GNAME22913(G22913,G8306);
  and GNAME22914(G22914,G22990,G22991);
  not GNAME22915(G22915,G8305);
  and GNAME22916(G22916,G22993,G22994);
  not GNAME22917(G22917,G8304);
  and GNAME22918(G22918,G22996,G22997);
  not GNAME22919(G22919,G8303);
  and GNAME22920(G22920,G9288,G22957,G9289);
  and GNAME22921(G22921,G9287,G22920);
  and GNAME22922(G22922,G22921,G9286,G9285);
  and GNAME22923(G22923,G9284,G22922);
  nand GNAME22924(G22924,G23008,G23009);
  nand GNAME22925(G22925,G23010,G23011);
  nand GNAME22926(G22926,G23012,G23013);
  nand GNAME22927(G22927,G23014,G23015);
  nand GNAME22928(G22928,G23016,G23017);
  nand GNAME22929(G22929,G23018,G23019);
  nand GNAME22930(G22930,G23020,G23021);
  nand GNAME22931(G22931,G23022,G23023);
  nand GNAME22932(G22932,G23024,G23025);
  nand GNAME22933(G22933,G23026,G23027);
  nand GNAME22934(G22934,G23028,G23029);
  nand GNAME22935(G22935,G23048,G23049);
  nand GNAME22936(G22936,G23064,G23065);
  nand GNAME22937(G22937,G23066,G23067);
  nand GNAME22938(G22938,G23068,G23069);
  nand GNAME22939(G22939,G23070,G23071);
  nand GNAME22940(G22940,G23072,G23073);
  nand GNAME22941(G22941,G23074,G23075);
  nand GNAME22942(G22942,G23076,G23077);
  nand GNAME22943(G22943,G23078,G23079);
  and GNAME22944(G22944,G23032,G23033);
  and GNAME22945(G22945,G23036,G23037);
  and GNAME22946(G22946,G23040,G23041);
  and GNAME22947(G22947,G23044,G23045);
  and GNAME22948(G22948,G23050,G23051);
  and GNAME22949(G22949,G23054,G23055);
  and GNAME22950(G22950,G23058,G23059);
  and GNAME22951(G22951,G23062,G23063);
  and GNAME22952(G22952,G22892,G8295);
  and GNAME22953(G22953,G22888,G8298);
  nand GNAME22954(G22954,G22923,G9283);
  not GNAME22955(G22955,G8300);
  nand GNAME22956(G22956,G22970,G9866);
  nand GNAME22957(G22957,G22999,G23000);
  and GNAME22958(G22958,G23030,G23031);
  and GNAME22959(G22959,G23034,G23035);
  and GNAME22960(G22960,G23038,G23039);
  and GNAME22961(G22961,G23042,G23043);
  and GNAME22962(G22962,G23046,G23047);
  and GNAME22963(G22963,G8302,G9866);
  and GNAME22964(G22964,G23052,G23053);
  and GNAME22965(G22965,G23056,G23057);
  and GNAME22966(G22966,G23060,G23061);
  and GNAME22967(G22967,G8288,G22902);
  and GNAME22968(G22968,G8290,G22900);
  and GNAME22969(G22969,G22976,G8292);
  nand GNAME22970(G22970,G8301,G8302);
  not GNAME22971(G22971,G22900);
  not GNAME22972(G22972,G22902);
  not GNAME22973(G22973,G22921);
  nand GNAME22974(G22974,G22955,G22970);
  not GNAME22975(G22975,G22884);
  not GNAME22976(G22976,G22897);
  or GNAME22977(G22977,G8286,G8310);
  nand GNAME22978(G22978,G22977,G22904);
  nand GNAME22979(G22979,G8310,G8286);
  nand GNAME22980(G22980,G22907,G22906);
  nand GNAME22981(G22981,G22980,G8285);
  or GNAME22982(G22982,G22906,G22907);
  nand GNAME22983(G22983,G22909,G22908);
  nand GNAME22984(G22984,G22983,G8284);
  or GNAME22985(G22985,G22908,G22909);
  nand GNAME22986(G22986,G22911,G22910);
  nand GNAME22987(G22987,G22986,G8283);
  or GNAME22988(G22988,G22910,G22911);
  nand GNAME22989(G22989,G22913,G22912);
  nand GNAME22990(G22990,G22989,G8282);
  or GNAME22991(G22991,G22912,G22913);
  nand GNAME22992(G22992,G22915,G22914);
  nand GNAME22993(G22993,G22992,G8281);
  or GNAME22994(G22994,G22914,G22915);
  nand GNAME22995(G22995,G22917,G22916);
  nand GNAME22996(G22996,G22995,G8280);
  or GNAME22997(G22997,G22916,G22917);
  nand GNAME22998(G22998,G22919,G22918);
  nand GNAME22999(G22999,G22998,G9290);
  or GNAME23000(G23000,G22918,G22919);
  or GNAME23001(G23001,G9284,G22922);
  and GNAME23002(G23002,G9286,G22921);
  nor GNAME23003(G23003,G23002,G9285);
  or GNAME23004(G23004,G9287,G22920);
  and GNAME23005(G23005,G22957,G9289);
  nor GNAME23006(G23006,G23005,G9288);
  not GNAME23007(G23007,G22956);
  nand GNAME23008(G23008,G22896,G22895);
  or GNAME23009(G23009,G22895,G22896);
  or GNAME23010(G23010,G22952,G22893);
  nand GNAME23011(G23011,G22893,G22952);
  or GNAME23012(G23012,G22892,G22894);
  nand GNAME23013(G23013,G22894,G22892);
  or GNAME23014(G23014,G8296,G23080);
  nand GNAME23015(G23015,G23080,G8296);
  or GNAME23016(G23016,G22953,G22890);
  nand GNAME23017(G23017,G22890,G22953);
  or GNAME23018(G23018,G22888,G22889);
  nand GNAME23019(G23019,G22889,G22888);
  nand GNAME23020(G23020,G22884,G8299);
  nand GNAME23021(G23021,G22887,G22975);
  nand GNAME23022(G23022,G22954,G8279);
  or GNAME23023(G23023,G8279,G22954);
  nand GNAME23024(G23024,G23081,G9283);
  or GNAME23025(G23025,G9283,G23081);
  nand GNAME23026(G23026,G22956,G8300);
  nand GNAME23027(G23027,G22955,G23007);
  or GNAME23028(G23028,G9286,G22973);
  nand GNAME23029(G23029,G22973,G9286);
  nand GNAME23030(G23030,G22957,G9289);
  or GNAME23031(G23031,G9289,G22957);
  nand GNAME23032(G23032,G22919,G9290);
  or GNAME23033(G23033,G9290,G22919);
  nand GNAME23034(G23034,G22918,G22944);
  or GNAME23035(G23035,G22918,G22944);
  nand GNAME23036(G23036,G22917,G8280);
  or GNAME23037(G23037,G8280,G22917);
  nand GNAME23038(G23038,G22916,G22945);
  or GNAME23039(G23039,G22916,G22945);
  nand GNAME23040(G23040,G22915,G8281);
  or GNAME23041(G23041,G8281,G22915);
  nand GNAME23042(G23042,G22914,G22946);
  or GNAME23043(G23043,G22914,G22946);
  nand GNAME23044(G23044,G22913,G8282);
  or GNAME23045(G23045,G8282,G22913);
  nand GNAME23046(G23046,G22912,G22947);
  or GNAME23047(G23047,G22912,G22947);
  or GNAME23048(G23048,G22963,G22885);
  nand GNAME23049(G23049,G22885,G22963);
  nand GNAME23050(G23050,G22911,G8283);
  or GNAME23051(G23051,G8283,G22911);
  nand GNAME23052(G23052,G22910,G22948);
  or GNAME23053(G23053,G22910,G22948);
  nand GNAME23054(G23054,G22909,G8284);
  or GNAME23055(G23055,G8284,G22909);
  nand GNAME23056(G23056,G22908,G22949);
  or GNAME23057(G23057,G22908,G22949);
  nand GNAME23058(G23058,G22907,G8285);
  or GNAME23059(G23059,G8285,G22907);
  nand GNAME23060(G23060,G22906,G22950);
  or GNAME23061(G23061,G22906,G22950);
  nand GNAME23062(G23062,G22905,G22904);
  or GNAME23063(G23063,G22904,G22905);
  nand GNAME23064(G23064,G8310,G22951);
  or GNAME23065(G23065,G8310,G22951);
  or GNAME23066(G23066,G22967,G22903);
  nand GNAME23067(G23067,G22903,G22967);
  or GNAME23068(G23068,G8288,G22972);
  nand GNAME23069(G23069,G22972,G8288);
  or GNAME23070(G23070,G22968,G22901);
  nand GNAME23071(G23071,G22901,G22968);
  or GNAME23072(G23072,G8290,G22971);
  nand GNAME23073(G23073,G22971,G8290);
  or GNAME23074(G23074,G22969,G22899);
  nand GNAME23075(G23075,G22899,G22969);
  nand GNAME23076(G23076,G22897,G8292);
  nand GNAME23077(G23077,G22898,G22976);
  or GNAME23078(G23078,G9866,G22886);
  nand GNAME23079(G23079,G22886,G9866);
  not GNAME23080(G23080,G22891);
  not GNAME23081(G23081,G22923);
  nand GNAME23082(G23082,G23084,G23085);
  not GNAME23083(G23083,G59567);
  nand GNAME23084(G23084,G23083,G59568);
  or GNAME23085(G23085,G59568,G23083);
  not GNAME23086(G23086,G9278);
  not GNAME23087(G23087,G9279);
  nand GNAME23088(G23088,G23115,G23118,G23119);
  not GNAME23089(G23089,G14132);
  not GNAME23090(G23090,G14136);
  not GNAME23091(G23091,G14143);
  not GNAME23092(G23092,G14134);
  not GNAME23093(G23093,G14141);
  not GNAME23094(G23094,G14131);
  not GNAME23095(G23095,G14137);
  nand GNAME23096(G23096,G23097,G23114);
  or GNAME23097(G23097,G14139,G23089);
  or GNAME23098(G23098,G14144,G23090);
  nand GNAME23099(G23099,G14145,G23095,G23098);
  or GNAME23100(G23100,G14135,G23091);
  nand GNAME23101(G23101,G23090,G14144);
  nand GNAME23102(G23102,G23101,G23099,G23100);
  or GNAME23103(G23103,G14142,G23092);
  nand GNAME23104(G23104,G23091,G14135);
  nand GNAME23105(G23105,G23104,G23102,G23103);
  or GNAME23106(G23106,G14133,G23093);
  nand GNAME23107(G23107,G23092,G14142);
  nand GNAME23108(G23108,G23107,G23105,G23106);
  or GNAME23109(G23109,G14140,G23089);
  nand GNAME23110(G23110,G23093,G14133);
  nand GNAME23111(G23111,G23110,G23108,G23109);
  or GNAME23112(G23112,G14140,G14139);
  nand GNAME23113(G23113,G23089,G23112);
  nand GNAME23114(G23114,G23113,G23111);
  nand GNAME23115(G23115,G23096,G23116,G23117);
  nand GNAME23116(G23116,G23094,G14138);
  or GNAME23117(G23117,G14138,G23094);
  nand GNAME23118(G23118,G23094,G14138,G14130);
  or GNAME23119(G23119,G23094,G14138,G14130);
  and GNAME23120(G23120,G23285,G23286);
  and GNAME23121(G23121,G23244,G23282);
  and GNAME23122(G23122,G23234,G23280);
  and GNAME23123(G23123,G23246,G23253);
  not GNAME23124(G23124,G14785);
  not GNAME23125(G23125,G14186);
  not GNAME23126(G23126,G14187);
  nor GNAME23127(G23127,G23243,G23155);
  nor GNAME23128(G23128,G23154,G23244);
  nor GNAME23129(G23129,G23153,G23229);
  nor GNAME23130(G23130,G23245,G23151,G23152);
  nor GNAME23131(G23131,G23150,G23246);
  not GNAME23132(G23132,G14185);
  not GNAME23133(G23133,G14184);
  not GNAME23134(G23134,G14183);
  not GNAME23135(G23135,G14182);
  not GNAME23136(G23136,G14181);
  not GNAME23137(G23137,G14180);
  not GNAME23138(G23138,G14179);
  not GNAME23139(G23139,G14178);
  nor GNAME23140(G23140,G23215,G23175);
  nor GNAME23141(G23141,G23402,G23173,G23174);
  nor GNAME23142(G23142,G23172,G23230);
  nor GNAME23143(G23143,G23277,G23170,G23171);
  nor GNAME23144(G23144,G23169,G23231);
  nor GNAME23145(G23145,G23278,G23167,G23168);
  nor GNAME23146(G23146,G23166,G23232);
  nor GNAME23147(G23147,G23279,G23164,G23165);
  or GNAME23148(G23148,G23233,G23162,G23163);
  and GNAME23149(G23149,G23264,G23236);
  and GNAME23150(G23150,G23292,G23293);
  and GNAME23151(G23151,G23306,G23307);
  and GNAME23152(G23152,G23308,G23309);
  and GNAME23153(G23153,G23294,G23295);
  and GNAME23154(G23154,G23296,G23297);
  and GNAME23155(G23155,G23304,G23305);
  nand GNAME23156(G23156,G23316,G23317);
  nand GNAME23157(G23157,G23318,G23319);
  nand GNAME23158(G23158,G23320,G23321);
  nand GNAME23159(G23159,G23322,G23323);
  nand GNAME23160(G23160,G23324,G23325);
  and GNAME23161(G23161,G23329,G23330);
  and GNAME23162(G23162,G23367,G23368);
  and GNAME23163(G23163,G23369,G23370);
  and GNAME23164(G23164,G23363,G23364);
  and GNAME23165(G23165,G23365,G23366);
  and GNAME23166(G23166,G23331,G23332);
  and GNAME23167(G23167,G23359,G23360);
  and GNAME23168(G23168,G23361,G23362);
  and GNAME23169(G23169,G23333,G23334);
  and GNAME23170(G23170,G23355,G23356);
  and GNAME23171(G23171,G23357,G23358);
  and GNAME23172(G23172,G23335,G23336);
  and GNAME23173(G23173,G23351,G23352);
  and GNAME23174(G23174,G23353,G23354);
  and GNAME23175(G23175,G23349,G23350);
  nand GNAME23176(G23176,G23373,G23374);
  nand GNAME23177(G23177,G23375,G23376);
  nand GNAME23178(G23178,G23377,G23378);
  nand GNAME23179(G23179,G23379,G23380);
  nand GNAME23180(G23180,G23381,G23382);
  nand GNAME23181(G23181,G23383,G23384);
  nand GNAME23182(G23182,G23385,G23386);
  nand GNAME23183(G23183,G23387,G23388);
  nand GNAME23184(G23184,G23389,G23390);
  nand GNAME23185(G23185,G23391,G23392);
  nand GNAME23186(G23186,G23395,G23396);
  nand GNAME23187(G23187,G23397,G23398);
  nand GNAME23188(G23188,G23399,G23400);
  nand GNAME23189(G23189,G23413,G23414);
  nand GNAME23190(G23190,G23371,G23372);
  nand GNAME23191(G23191,G23405,G23406);
  nand GNAME23192(G23192,G23411,G23412);
  not GNAME23193(G23193,G14169);
  not GNAME23194(G23194,G14176);
  not GNAME23195(G23195,G14177);
  not GNAME23196(G23196,G14168);
  nand GNAME23197(G23197,G23249,G23247);
  and GNAME23198(G23198,G23251,G23250);
  and GNAME23199(G23199,G23314,G23315);
  nand GNAME23200(G23200,G23248,G23247);
  not GNAME23201(G23201,G14146);
  not GNAME23202(G23202,G14166);
  not GNAME23203(G23203,G14165);
  not GNAME23204(G23204,G14164);
  not GNAME23205(G23205,G14162);
  nor GNAME23206(G23206,G23161,G23148);
  nor GNAME23207(G23207,G23163,G23233);
  nor GNAME23208(G23208,G23164,G23279);
  nor GNAME23209(G23209,G23167,G23278);
  nor GNAME23210(G23210,G23170,G23277);
  nand GNAME23211(G23211,G23241,G23239);
  and GNAME23212(G23212,G23242,G23238);
  and GNAME23213(G23213,G23393,G23394);
  nor GNAME23214(G23214,G23173,G23402);
  and GNAME23215(G23215,G23276,G23254);
  and GNAME23216(G23216,G23401,G23402);
  nand GNAME23217(G23217,G23274,G23237);
  and GNAME23218(G23218,G23275,G23254);
  and GNAME23219(G23219,G23403,G23404);
  and GNAME23220(G23220,G23272,G23258);
  nand GNAME23221(G23221,G23270,G23259);
  and GNAME23222(G23222,G23271,G23258);
  and GNAME23223(G23223,G23407,G23408);
  nand GNAME23224(G23224,G23268,G23260);
  and GNAME23225(G23225,G23269,G23259);
  and GNAME23226(G23226,G23409,G23410);
  nor GNAME23227(G23227,G23415,G23149);
  and GNAME23228(G23228,G23240,G23239);
  not GNAME23229(G23229,G23128);
  not GNAME23230(G23230,G23141);
  not GNAME23231(G23231,G23143);
  not GNAME23232(G23232,G23145);
  not GNAME23233(G23233,G23147);
  not GNAME23234(G23234,G23206);
  nand GNAME23235(G23235,G23256,G23138,G23255);
  nand GNAME23236(G23236,G23263,G23134,G23262);
  nand GNAME23237(G23237,G23257,G14179);
  nand GNAME23238(G23238,G23300,G14186);
  nand GNAME23239(G23239,G23303,G14187);
  nand GNAME23240(G23240,G23126,G23301,G23302);
  nand GNAME23241(G23241,G23240,G14785);
  nand GNAME23242(G23242,G23125,G23298,G23299);
  and GNAME23243(G23243,G23238,G23281);
  not GNAME23244(G23244,G23127);
  not GNAME23245(G23245,G23129);
  not GNAME23246(G23246,G23130);
  nand GNAME23247(G23247,G23310,G14185);
  nand GNAME23248(G23248,G23132,G23290,G23291);
  nand GNAME23249(G23249,G23248,G23131);
  nand GNAME23250(G23250,G23313,G14184);
  nand GNAME23251(G23251,G23133,G23311,G23312);
  or GNAME23252(G23252,G23151,G23245);
  nand GNAME23253(G23253,G23252,G23152);
  nand GNAME23254(G23254,G23348,G14178);
  or GNAME23255(G23255,G14163,G23124);
  nand GNAME23256(G23256,G23124,G14163);
  nand GNAME23257(G23257,G23256,G23255);
  nand GNAME23258(G23258,G23345,G14180);
  nand GNAME23259(G23259,G23342,G14181);
  nand GNAME23260(G23260,G23339,G14182);
  nand GNAME23261(G23261,G23135,G23337,G23338);
  or GNAME23262(G23262,G14167,G23124);
  nand GNAME23263(G23263,G23124,G14167);
  nand GNAME23264(G23264,G23250,G23284);
  nand GNAME23265(G23265,G23262,G23263);
  nand GNAME23266(G23266,G23265,G14183);
  not GNAME23267(G23267,G23227);
  nand GNAME23268(G23268,G23261,G23267);
  nand GNAME23269(G23269,G23136,G23340,G23341);
  nand GNAME23270(G23270,G23224,G23269);
  nand GNAME23271(G23271,G23137,G23343,G23344);
  nand GNAME23272(G23272,G23221,G23271);
  not GNAME23273(G23273,G23220);
  nand GNAME23274(G23274,G23235,G23273);
  nand GNAME23275(G23275,G23139,G23346,G23347);
  nand GNAME23276(G23276,G23217,G23275);
  not GNAME23277(G23277,G23142);
  not GNAME23278(G23278,G23144);
  not GNAME23279(G23279,G23146);
  nand GNAME23280(G23280,G23148,G23161);
  nand GNAME23281(G23281,G23211,G23242);
  nand GNAME23282(G23282,G23155,G23238,G23281);
  nand GNAME23283(G23283,G23236,G23266);
  nand GNAME23284(G23284,G23197,G23251);
  nand GNAME23285(G23285,G23284,G23250,G23283);
  nand GNAME23286(G23286,G23266,G23149);
  not GNAME23287(G23287,G23228);
  nand GNAME23288(G23288,G23235,G23237);
  nand GNAME23289(G23289,G23260,G23261);
  or GNAME23290(G23290,G14169,G23124);
  or GNAME23291(G23291,G14785,G23193);
  or GNAME23292(G23292,G14170,G23124);
  nand GNAME23293(G23293,G23124,G14170);
  or GNAME23294(G23294,G14173,G23124);
  nand GNAME23295(G23295,G23124,G14173);
  or GNAME23296(G23296,G14174,G23124);
  nand GNAME23297(G23297,G23124,G14174);
  or GNAME23298(G23298,G14176,G23124);
  or GNAME23299(G23299,G14785,G23194);
  nand GNAME23300(G23300,G23298,G23299);
  or GNAME23301(G23301,G14177,G23124);
  or GNAME23302(G23302,G14785,G23195);
  nand GNAME23303(G23303,G23301,G23302);
  or GNAME23304(G23304,G14175,G23124);
  nand GNAME23305(G23305,G23124,G14175);
  or GNAME23306(G23306,G14172,G23124);
  nand GNAME23307(G23307,G23124,G14172);
  or GNAME23308(G23308,G14171,G23124);
  nand GNAME23309(G23309,G23124,G14171);
  nand GNAME23310(G23310,G23290,G23291);
  or GNAME23311(G23311,G14168,G23124);
  or GNAME23312(G23312,G14785,G23196);
  nand GNAME23313(G23313,G23311,G23312);
  or GNAME23314(G23314,G23198,G23197);
  nand GNAME23315(G23315,G23197,G23198);
  nand GNAME23316(G23316,G23200,G23131);
  or GNAME23317(G23317,G23131,G23200);
  nand GNAME23318(G23318,G23130,G23150);
  or GNAME23319(G23319,G23130,G23150);
  nand GNAME23320(G23320,G23129,G23151);
  or GNAME23321(G23321,G23129,G23151);
  nand GNAME23322(G23322,G23128,G23153);
  or GNAME23323(G23323,G23128,G23153);
  nand GNAME23324(G23324,G23127,G23154);
  or GNAME23325(G23325,G23127,G23154);
  or GNAME23326(G23326,G14146,G23124);
  or GNAME23327(G23327,G14785,G23201);
  nand GNAME23328(G23328,G23326,G23327);
  or GNAME23329(G23329,G14147,G23124);
  nand GNAME23330(G23330,G23124,G14147);
  or GNAME23331(G23331,G14152,G23124);
  nand GNAME23332(G23332,G23124,G14152);
  or GNAME23333(G23333,G14155,G23124);
  nand GNAME23334(G23334,G23124,G14155);
  or GNAME23335(G23335,G14158,G23124);
  nand GNAME23336(G23336,G23124,G14158);
  or GNAME23337(G23337,G14166,G23124);
  or GNAME23338(G23338,G14785,G23202);
  nand GNAME23339(G23339,G23337,G23338);
  or GNAME23340(G23340,G14165,G23124);
  or GNAME23341(G23341,G14785,G23203);
  nand GNAME23342(G23342,G23340,G23341);
  or GNAME23343(G23343,G14164,G23124);
  or GNAME23344(G23344,G14785,G23204);
  nand GNAME23345(G23345,G23343,G23344);
  or GNAME23346(G23346,G14162,G23124);
  or GNAME23347(G23347,G14785,G23205);
  nand GNAME23348(G23348,G23346,G23347);
  or GNAME23349(G23349,G14161,G23124);
  nand GNAME23350(G23350,G23124,G14161);
  or GNAME23351(G23351,G14160,G23124);
  nand GNAME23352(G23352,G23124,G14160);
  or GNAME23353(G23353,G14159,G23124);
  nand GNAME23354(G23354,G23124,G14159);
  or GNAME23355(G23355,G14157,G23124);
  nand GNAME23356(G23356,G23124,G14157);
  or GNAME23357(G23357,G14156,G23124);
  nand GNAME23358(G23358,G23124,G14156);
  or GNAME23359(G23359,G14154,G23124);
  nand GNAME23360(G23360,G23124,G14154);
  or GNAME23361(G23361,G14153,G23124);
  nand GNAME23362(G23362,G23124,G14153);
  or GNAME23363(G23363,G14151,G23124);
  nand GNAME23364(G23364,G23124,G14151);
  or GNAME23365(G23365,G14150,G23124);
  nand GNAME23366(G23366,G23124,G14150);
  or GNAME23367(G23367,G14148,G23124);
  nand GNAME23368(G23368,G23124,G14148);
  or GNAME23369(G23369,G14149,G23124);
  nand GNAME23370(G23370,G23124,G14149);
  nand GNAME23371(G23371,G23234,G23328);
  nand GNAME23372(G23372,G23206,G23326,G23327);
  nand GNAME23373(G23373,G23162,G23207);
  or GNAME23374(G23374,G23207,G23162);
  nand GNAME23375(G23375,G23147,G23163);
  or GNAME23376(G23376,G23147,G23163);
  nand GNAME23377(G23377,G23165,G23208);
  or GNAME23378(G23378,G23208,G23165);
  nand GNAME23379(G23379,G23146,G23164);
  or GNAME23380(G23380,G23146,G23164);
  nand GNAME23381(G23381,G23145,G23166);
  or GNAME23382(G23382,G23145,G23166);
  nand GNAME23383(G23383,G23168,G23209);
  or GNAME23384(G23384,G23209,G23168);
  nand GNAME23385(G23385,G23144,G23167);
  or GNAME23386(G23386,G23144,G23167);
  nand GNAME23387(G23387,G23143,G23169);
  or GNAME23388(G23388,G23143,G23169);
  nand GNAME23389(G23389,G23171,G23210);
  or GNAME23390(G23390,G23210,G23171);
  nand GNAME23391(G23391,G23142,G23170);
  or GNAME23392(G23392,G23142,G23170);
  or GNAME23393(G23393,G23212,G23211);
  nand GNAME23394(G23394,G23211,G23212);
  nand GNAME23395(G23395,G23141,G23172);
  or GNAME23396(G23396,G23141,G23172);
  nand GNAME23397(G23397,G23174,G23214);
  or GNAME23398(G23398,G23214,G23174);
  nand GNAME23399(G23399,G23140,G23173);
  or GNAME23400(G23400,G23140,G23173);
  nand GNAME23401(G23401,G23175,G23215);
  or GNAME23402(G23402,G23215,G23175);
  or GNAME23403(G23403,G23218,G23217);
  nand GNAME23404(G23404,G23217,G23218);
  nand GNAME23405(G23405,G23273,G23288);
  nand GNAME23406(G23406,G23220,G23235,G23237);
  or GNAME23407(G23407,G23222,G23221);
  nand GNAME23408(G23408,G23221,G23222);
  or GNAME23409(G23409,G23225,G23224);
  nand GNAME23410(G23410,G23224,G23225);
  nand GNAME23411(G23411,G23267,G23289);
  nand GNAME23412(G23412,G23227,G23260,G23261);
  or GNAME23413(G23413,G23228,G23124);
  or GNAME23414(G23414,G14785,G23287);
  not GNAME23415(G23415,G23266);
  not GNAME23416(G23416,G14115);
  not GNAME23417(G23417,G14120);
  not GNAME23418(G23418,G14114);
  not GNAME23419(G23419,G14116);
  not GNAME23420(G23420,G14121);
  not GNAME23421(G23421,G14118);
  not GNAME23422(G23422,G14119);
  not GNAME23423(G23423,G14117);
  and GNAME23424(G23424,G23591,G23615);
  and GNAME23425(G23425,G23545,G23613);
  and GNAME23426(G23426,G23610,G23611);
  and GNAME23427(G23427,G23546,G23607);
  and GNAME23428(G23428,G23580,G23581);
  not GNAME23429(G23429,G14830);
  not GNAME23430(G23430,G14229);
  not GNAME23431(G23431,G14230);
  not GNAME23432(G23432,G14233);
  not GNAME23433(G23433,G14234);
  not GNAME23434(G23434,G14235);
  not GNAME23435(G23435,G14232);
  not GNAME23436(G23436,G14231);
  not GNAME23437(G23437,G14228);
  nor GNAME23438(G23438,G23495,G23460);
  and GNAME23439(G23439,G23573,G23547);
  nor GNAME23440(G23440,G23644,G23459,G23473);
  nor GNAME23441(G23441,G23472,G23591);
  nor GNAME23442(G23442,G23471,G23544);
  nor GNAME23443(G23443,G23549,G23469,G23470);
  nor GNAME23444(G23444,G23468,G23545);
  not GNAME23445(G23445,G14227);
  not GNAME23446(G23446,G14226);
  not GNAME23447(G23447,G14225);
  not GNAME23448(G23448,G14224);
  not GNAME23449(G23449,G14223);
  not GNAME23450(G23450,G14222);
  not GNAME23451(G23451,G14221);
  not GNAME23452(G23452,G14220);
  nor GNAME23453(G23453,G23516,G23474);
  nor GNAME23454(G23454,G23719,G23466,G23467);
  and GNAME23455(G23455,G23750,G23454);
  nor GNAME23456(G23456,G23464,G23751);
  nand GNAME23457(G23457,G23752,G23456);
  and GNAME23458(G23458,G23565,G23548);
  and GNAME23459(G23459,G23639,G23640);
  and GNAME23460(G23460,G23637,G23638);
  nand GNAME23461(G23461,G23641,G23642);
  and GNAME23462(G23462,G23656,G23657);
  and GNAME23463(G23463,G23658,G23659);
  and GNAME23464(G23464,G23660,G23661);
  and GNAME23465(G23465,G23662,G23663);
  and GNAME23466(G23466,G23702,G23703);
  and GNAME23467(G23467,G23704,G23705);
  and GNAME23468(G23468,G23666,G23667);
  and GNAME23469(G23469,G23674,G23675);
  and GNAME23470(G23470,G23676,G23677);
  and GNAME23471(G23471,G23668,G23669);
  and GNAME23472(G23472,G23670,G23671);
  and GNAME23473(G23473,G23672,G23673);
  and GNAME23474(G23474,G23700,G23701);
  nand GNAME23475(G23475,G23708,G23709);
  nand GNAME23476(G23476,G23710,G23711);
  nand GNAME23477(G23477,G23712,G23713);
  nand GNAME23478(G23478,G23714,G23715);
  nand GNAME23479(G23479,G23716,G23717);
  nand GNAME23480(G23480,G23736,G23737);
  nand GNAME23481(G23481,G23738,G23739);
  nand GNAME23482(G23482,G23740,G23741);
  nand GNAME23483(G23483,G23742,G23743);
  nand GNAME23484(G23484,G23744,G23745);
  nand GNAME23485(G23485,G23746,G23747);
  nand GNAME23486(G23486,G23645,G23646);
  nand GNAME23487(G23487,G23651,G23652);
  nand GNAME23488(G23488,G23706,G23707);
  not GNAME23489(G23489,G14212);
  not GNAME23490(G23490,G14214);
  not GNAME23491(G23491,G14216);
  not GNAME23492(G23492,G14218);
  not GNAME23493(G23493,G14219);
  not GNAME23494(G23494,G14215);
  and GNAME23495(G23495,G23577,G23550);
  and GNAME23496(G23496,G23643,G23644);
  nor GNAME23497(G23497,G23749,G23439);
  nand GNAME23498(G23498,G23571,G23555);
  and GNAME23499(G23499,G23572,G23552);
  and GNAME23500(G23500,G23647,G23648);
  nand GNAME23501(G23501,G23569,G23556);
  and GNAME23502(G23502,G23570,G23555);
  and GNAME23503(G23503,G23649,G23650);
  nor GNAME23504(G23504,G23748,G23458);
  not GNAME23505(G23505,G14188);
  not GNAME23506(G23506,G14203);
  not GNAME23507(G23507,G14202);
  not GNAME23508(G23508,G14201);
  not GNAME23509(G23509,G14200);
  not GNAME23510(G23510,G14199);
  not GNAME23511(G23511,G14198);
  not GNAME23512(G23512,G14197);
  not GNAME23513(G23513,G14196);
  nor GNAME23514(G23514,G23462,G23457);
  nor GNAME23515(G23515,G23467,G23719);
  and GNAME23516(G23516,G23606,G23582);
  and GNAME23517(G23517,G23718,G23719);
  nand GNAME23518(G23518,G23604,G23583);
  and GNAME23519(G23519,G23605,G23582);
  and GNAME23520(G23520,G23720,G23721);
  nand GNAME23521(G23521,G23602,G23584);
  and GNAME23522(G23522,G23603,G23583);
  and GNAME23523(G23523,G23722,G23723);
  nand GNAME23524(G23524,G23600,G23585);
  and GNAME23525(G23525,G23601,G23584);
  and GNAME23526(G23526,G23724,G23725);
  nand GNAME23527(G23527,G23598,G23586);
  and GNAME23528(G23528,G23599,G23585);
  and GNAME23529(G23529,G23726,G23727);
  nand GNAME23530(G23530,G23563,G23561);
  and GNAME23531(G23531,G23564,G23558);
  and GNAME23532(G23532,G23728,G23729);
  nand GNAME23533(G23533,G23596,G23587);
  and GNAME23534(G23534,G23597,G23586);
  and GNAME23535(G23535,G23730,G23731);
  nand GNAME23536(G23536,G23594,G23588);
  and GNAME23537(G23537,G23595,G23587);
  and GNAME23538(G23538,G23732,G23733);
  nand GNAME23539(G23539,G23592,G23589);
  and GNAME23540(G23540,G23593,G23588);
  and GNAME23541(G23541,G23734,G23735);
  nand GNAME23542(G23542,G23590,G23589);
  and GNAME23543(G23543,G23562,G23561);
  not GNAME23544(G23544,G23441);
  not GNAME23545(G23545,G23443);
  not GNAME23546(G23546,G23514);
  nand GNAME23547(G23547,G23554,G23430,G23553);
  nand GNAME23548(G23548,G23560,G23432,G23559);
  not GNAME23549(G23549,G23442);
  nand GNAME23550(G23550,G23636,G14228);
  nand GNAME23551(G23551,G23437,G23619,G23620);
  nand GNAME23552(G23552,G23623,G14230);
  or GNAME23553(G23553,G14213,G23429);
  nand GNAME23554(G23554,G23429,G14213);
  nand GNAME23555(G23555,G23635,G14231);
  nand GNAME23556(G23556,G23632,G14232);
  nand GNAME23557(G23557,G23435,G23624,G23625);
  nand GNAME23558(G23558,G23628,G14234);
  or GNAME23559(G23559,G14217,G23429);
  nand GNAME23560(G23560,G23429,G14217);
  nand GNAME23561(G23561,G23631,G14235);
  nand GNAME23562(G23562,G23434,G23629,G23630);
  nand GNAME23563(G23563,G23562,G14830);
  nand GNAME23564(G23564,G23433,G23626,G23627);
  nand GNAME23565(G23565,G23558,G23608);
  nand GNAME23566(G23566,G23559,G23560);
  nand GNAME23567(G23567,G23566,G14233);
  not GNAME23568(G23568,G23504);
  nand GNAME23569(G23569,G23557,G23568);
  nand GNAME23570(G23570,G23436,G23633,G23634);
  nand GNAME23571(G23571,G23501,G23570);
  nand GNAME23572(G23572,G23431,G23621,G23622);
  nand GNAME23573(G23573,G23552,G23578);
  nand GNAME23574(G23574,G23553,G23554);
  nand GNAME23575(G23575,G23574,G14229);
  not GNAME23576(G23576,G23497);
  nand GNAME23577(G23577,G23551,G23576);
  nand GNAME23578(G23578,G23498,G23572);
  nand GNAME23579(G23579,G23547,G23575);
  nand GNAME23580(G23580,G23579,G23552,G23578);
  nand GNAME23581(G23581,G23575,G23439);
  nand GNAME23582(G23582,G23699,G14220);
  nand GNAME23583(G23583,G23696,G14221);
  nand GNAME23584(G23584,G23693,G14222);
  nand GNAME23585(G23585,G23690,G14223);
  nand GNAME23586(G23586,G23687,G14224);
  nand GNAME23587(G23587,G23684,G14225);
  nand GNAME23588(G23588,G23681,G14226);
  nand GNAME23589(G23589,G23678,G14227);
  nand GNAME23590(G23590,G23445,G23664,G23665);
  not GNAME23591(G23591,G23440);
  nand GNAME23592(G23592,G23590,G23444);
  nand GNAME23593(G23593,G23446,G23679,G23680);
  nand GNAME23594(G23594,G23539,G23593);
  nand GNAME23595(G23595,G23447,G23682,G23683);
  nand GNAME23596(G23596,G23536,G23595);
  nand GNAME23597(G23597,G23448,G23685,G23686);
  nand GNAME23598(G23598,G23533,G23597);
  nand GNAME23599(G23599,G23449,G23688,G23689);
  nand GNAME23600(G23600,G23527,G23599);
  nand GNAME23601(G23601,G23450,G23691,G23692);
  nand GNAME23602(G23602,G23524,G23601);
  nand GNAME23603(G23603,G23451,G23694,G23695);
  nand GNAME23604(G23604,G23521,G23603);
  nand GNAME23605(G23605,G23452,G23697,G23698);
  nand GNAME23606(G23606,G23518,G23605);
  nand GNAME23607(G23607,G23457,G23462);
  nand GNAME23608(G23608,G23530,G23564);
  nand GNAME23609(G23609,G23548,G23567);
  nand GNAME23610(G23610,G23609,G23558,G23608);
  nand GNAME23611(G23611,G23567,G23458);
  or GNAME23612(G23612,G23469,G23549);
  nand GNAME23613(G23613,G23612,G23470);
  or GNAME23614(G23614,G23459,G23644);
  nand GNAME23615(G23615,G23614,G23473);
  not GNAME23616(G23616,G23543);
  nand GNAME23617(G23617,G23550,G23551);
  nand GNAME23618(G23618,G23556,G23557);
  or GNAME23619(G23619,G14212,G23429);
  or GNAME23620(G23620,G14830,G23489);
  or GNAME23621(G23621,G14214,G23429);
  or GNAME23622(G23622,G14830,G23490);
  nand GNAME23623(G23623,G23621,G23622);
  or GNAME23624(G23624,G14216,G23429);
  or GNAME23625(G23625,G14830,G23491);
  or GNAME23626(G23626,G14218,G23429);
  or GNAME23627(G23627,G14830,G23492);
  nand GNAME23628(G23628,G23626,G23627);
  or GNAME23629(G23629,G14219,G23429);
  or GNAME23630(G23630,G14830,G23493);
  nand GNAME23631(G23631,G23629,G23630);
  nand GNAME23632(G23632,G23624,G23625);
  or GNAME23633(G23633,G14215,G23429);
  or GNAME23634(G23634,G14830,G23494);
  nand GNAME23635(G23635,G23633,G23634);
  nand GNAME23636(G23636,G23619,G23620);
  or GNAME23637(G23637,G14211,G23429);
  nand GNAME23638(G23638,G23429,G14211);
  or GNAME23639(G23639,G14210,G23429);
  nand GNAME23640(G23640,G23429,G14210);
  nand GNAME23641(G23641,G23438,G23459);
  or GNAME23642(G23642,G23438,G23459);
  nand GNAME23643(G23643,G23460,G23495);
  or GNAME23644(G23644,G23495,G23460);
  nand GNAME23645(G23645,G23576,G23617);
  nand GNAME23646(G23646,G23497,G23550,G23551);
  or GNAME23647(G23647,G23499,G23498);
  nand GNAME23648(G23648,G23498,G23499);
  or GNAME23649(G23649,G23502,G23501);
  nand GNAME23650(G23650,G23501,G23502);
  nand GNAME23651(G23651,G23568,G23618);
  nand GNAME23652(G23652,G23504,G23556,G23557);
  or GNAME23653(G23653,G14188,G23429);
  or GNAME23654(G23654,G14830,G23505);
  nand GNAME23655(G23655,G23653,G23654);
  or GNAME23656(G23656,G14189,G23429);
  nand GNAME23657(G23657,G23429,G14189);
  or GNAME23658(G23658,G14190,G23429);
  nand GNAME23659(G23659,G23429,G14190);
  or GNAME23660(G23660,G14191,G23429);
  nand GNAME23661(G23661,G23429,G14191);
  or GNAME23662(G23662,G14192,G23429);
  nand GNAME23663(G23663,G23429,G14192);
  or GNAME23664(G23664,G14203,G23429);
  or GNAME23665(G23665,G14830,G23506);
  or GNAME23666(G23666,G14204,G23429);
  nand GNAME23667(G23667,G23429,G14204);
  or GNAME23668(G23668,G14207,G23429);
  nand GNAME23669(G23669,G23429,G14207);
  or GNAME23670(G23670,G14208,G23429);
  nand GNAME23671(G23671,G23429,G14208);
  or GNAME23672(G23672,G14209,G23429);
  nand GNAME23673(G23673,G23429,G14209);
  or GNAME23674(G23674,G14206,G23429);
  nand GNAME23675(G23675,G23429,G14206);
  or GNAME23676(G23676,G14205,G23429);
  nand GNAME23677(G23677,G23429,G14205);
  nand GNAME23678(G23678,G23664,G23665);
  or GNAME23679(G23679,G14202,G23429);
  or GNAME23680(G23680,G14830,G23507);
  nand GNAME23681(G23681,G23679,G23680);
  or GNAME23682(G23682,G14201,G23429);
  or GNAME23683(G23683,G14830,G23508);
  nand GNAME23684(G23684,G23682,G23683);
  or GNAME23685(G23685,G14200,G23429);
  or GNAME23686(G23686,G14830,G23509);
  nand GNAME23687(G23687,G23685,G23686);
  or GNAME23688(G23688,G14199,G23429);
  or GNAME23689(G23689,G14830,G23510);
  nand GNAME23690(G23690,G23688,G23689);
  or GNAME23691(G23691,G14198,G23429);
  or GNAME23692(G23692,G14830,G23511);
  nand GNAME23693(G23693,G23691,G23692);
  or GNAME23694(G23694,G14197,G23429);
  or GNAME23695(G23695,G14830,G23512);
  nand GNAME23696(G23696,G23694,G23695);
  or GNAME23697(G23697,G14196,G23429);
  or GNAME23698(G23698,G14830,G23513);
  nand GNAME23699(G23699,G23697,G23698);
  or GNAME23700(G23700,G14195,G23429);
  nand GNAME23701(G23701,G23429,G14195);
  or GNAME23702(G23702,G14193,G23429);
  nand GNAME23703(G23703,G23429,G14193);
  or GNAME23704(G23704,G14194,G23429);
  nand GNAME23705(G23705,G23429,G14194);
  nand GNAME23706(G23706,G23546,G23655);
  nand GNAME23707(G23707,G23514,G23653,G23654);
  nand GNAME23708(G23708,G23456,G23463);
  or GNAME23709(G23709,G23456,G23463);
  nand GNAME23710(G23710,G23455,G23464);
  or GNAME23711(G23711,G23455,G23464);
  nand GNAME23712(G23712,G23454,G23465);
  or GNAME23713(G23713,G23454,G23465);
  nand GNAME23714(G23714,G23466,G23515);
  or GNAME23715(G23715,G23515,G23466);
  nand GNAME23716(G23716,G23453,G23467);
  or GNAME23717(G23717,G23453,G23467);
  nand GNAME23718(G23718,G23474,G23516);
  or GNAME23719(G23719,G23516,G23474);
  or GNAME23720(G23720,G23519,G23518);
  nand GNAME23721(G23721,G23518,G23519);
  or GNAME23722(G23722,G23522,G23521);
  nand GNAME23723(G23723,G23521,G23522);
  or GNAME23724(G23724,G23525,G23524);
  nand GNAME23725(G23725,G23524,G23525);
  or GNAME23726(G23726,G23528,G23527);
  nand GNAME23727(G23727,G23527,G23528);
  or GNAME23728(G23728,G23531,G23530);
  nand GNAME23729(G23729,G23530,G23531);
  or GNAME23730(G23730,G23534,G23533);
  nand GNAME23731(G23731,G23533,G23534);
  or GNAME23732(G23732,G23537,G23536);
  nand GNAME23733(G23733,G23536,G23537);
  or GNAME23734(G23734,G23540,G23539);
  nand GNAME23735(G23735,G23539,G23540);
  nand GNAME23736(G23736,G23542,G23444);
  or GNAME23737(G23737,G23444,G23542);
  nand GNAME23738(G23738,G23443,G23468);
  or GNAME23739(G23739,G23443,G23468);
  nand GNAME23740(G23740,G23442,G23469);
  or GNAME23741(G23741,G23442,G23469);
  nand GNAME23742(G23742,G23441,G23471);
  or GNAME23743(G23743,G23441,G23471);
  nand GNAME23744(G23744,G23440,G23472);
  or GNAME23745(G23745,G23440,G23472);
  or GNAME23746(G23746,G23543,G23429);
  or GNAME23747(G23747,G14830,G23616);
  not GNAME23748(G23748,G23567);
  not GNAME23749(G23749,G23575);
  not GNAME23750(G23750,G23465);
  not GNAME23751(G23751,G23455);
  not GNAME23752(G23752,G23463);
  nor GNAME23753(G23753,G23756,G23784);
  and GNAME23754(G23754,G23763,G23761,G23762);
  and GNAME23755(G23755,G23758,G23800);
  nor GNAME23756(G23756,G23755,G23754,G23799,G23798);
  not GNAME23757(G23757,G23797);
  not GNAME23758(G23758,G15846);
  not GNAME23759(G23759,G23785);
  or GNAME23760(G23760,G15778,G23757);
  nand GNAME23761(G23761,G15779,G23759,G23760);
  or GNAME23762(G23762,G23800,G23758);
  nand GNAME23763(G23763,G23757,G15778);
  or GNAME23764(G23764,G15274,G23765);
  nor GNAME23765(G23765,G1551,G1550);
  and GNAME23766(G23766,G23782,G23783);
  not GNAME23767(G23767,G15277);
  not GNAME23768(G23768,G60013);
  not GNAME23769(G23769,G15275);
  not GNAME23770(G23770,G15274);
  not GNAME23771(G23771,G15278);
  or GNAME23772(G23772,G60014,G23767);
  nand GNAME23773(G23773,G60015,G23771,G23772);
  or GNAME23774(G23774,G15276,G23768);
  nand GNAME23775(G23775,G23767,G60014);
  nand GNAME23776(G23776,G23775,G23773,G23774);
  or GNAME23777(G23777,G60012,G23769);
  nand GNAME23778(G23778,G23768,G15276);
  nand GNAME23779(G23779,G23778,G23776,G23777);
  nand GNAME23780(G23780,G23770,G60011);
  nand GNAME23781(G23781,G23769,G60012);
  nand GNAME23782(G23782,G23781,G23779,G23780);
  or GNAME23783(G23783,G60011,G23770);
  nand GNAME23784(G23784,G23816,G23817);
  nand GNAME23785(G23785,G23818,G23804);
  not GNAME23786(G23786,G60010);
  not GNAME23787(G23787,G60009);
  not GNAME23788(G23788,G60014);
  and GNAME23789(G23789,G23805,G23835);
  not GNAME23790(G23790,G60008);
  not GNAME23791(G23791,G60013);
  and GNAME23792(G23792,G23808,G23809);
  not GNAME23793(G23793,G60007);
  not GNAME23794(G23794,G60012);
  and GNAME23795(G23795,G23812,G23813);
  not GNAME23796(G23796,G60006);
  nand GNAME23797(G23797,G23836,G23837);
  nand GNAME23798(G23798,G23822,G23823);
  nand GNAME23799(G23799,G23827,G23828);
  nand GNAME23800(G23800,G23832,G23833);
  and GNAME23801(G23801,G23834,G23835);
  not GNAME23802(G23802,G60011);
  nor GNAME23803(G23803,G60015,G23786);
  not GNAME23804(G23804,G23803);
  nand GNAME23805(G23805,G23804,G23834);
  not GNAME23806(G23806,G23789);
  or GNAME23807(G23807,G23806,G23790);
  nand GNAME23808(G23808,G23807,G60013);
  or GNAME23809(G23809,G60008,G23789);
  not GNAME23810(G23810,G23792);
  or GNAME23811(G23811,G23810,G23793);
  nand GNAME23812(G23812,G23811,G60012);
  or GNAME23813(G23813,G60007,G23792);
  not GNAME23814(G23814,G23795);
  or GNAME23815(G23815,G23795,G60006);
  nand GNAME23816(G23816,G23802,G23815);
  or GNAME23817(G23817,G23814,G23796);
  nand GNAME23818(G23818,G23786,G60015);
  or GNAME23819(G23819,G60006,G23802);
  or GNAME23820(G23820,G60011,G23796);
  nand GNAME23821(G23821,G23819,G23820);
  nand GNAME23822(G23822,G23814,G23821);
  nand GNAME23823(G23823,G23795,G23819,G23820);
  or GNAME23824(G23824,G60007,G23794);
  or GNAME23825(G23825,G60012,G23793);
  nand GNAME23826(G23826,G23824,G23825);
  nand GNAME23827(G23827,G23810,G23826);
  nand GNAME23828(G23828,G23792,G23824,G23825);
  or GNAME23829(G23829,G60008,G23791);
  or GNAME23830(G23830,G60013,G23790);
  nand GNAME23831(G23831,G23829,G23830);
  nand GNAME23832(G23832,G23806,G23831);
  nand GNAME23833(G23833,G23789,G23829,G23830);
  or GNAME23834(G23834,G60014,G23787);
  or GNAME23835(G23835,G60009,G23788);
  nand GNAME23836(G23836,G23801,G23803);
  or GNAME23837(G23837,G23803,G23801);
  and GNAME23838(G23838,G24080,G24081);
  and GNAME23839(G23839,G24075,G24076);
  and GNAME23840(G23840,G24069,G24070);
  and GNAME23841(G23841,G23996,G23997);
  not GNAME23842(G23842,G15181);
  not GNAME23843(G23843,G14269);
  not GNAME23844(G23844,G14270);
  not GNAME23845(G23845,G14273);
  not GNAME23846(G23846,G14274);
  not GNAME23847(G23847,G14275);
  not GNAME23848(G23848,G14272);
  not GNAME23849(G23849,G14271);
  not GNAME23850(G23850,G14268);
  and GNAME23851(G23851,G23990,G23963);
  not GNAME23852(G23852,G14267);
  and GNAME23853(G23853,G23986,G23961);
  or GNAME23854(G23854,G23998,G23929);
  not GNAME23855(G23855,G14264);
  and GNAME23856(G23856,G24001,G24002);
  not GNAME23857(G23857,G14263);
  not GNAME23858(G23858,G14262);
  nand GNAME23859(G23859,G24004,G24005);
  nand GNAME23860(G23860,G24008,G24009);
  not GNAME23861(G23861,G14261);
  and GNAME23862(G23862,G24012,G24013);
  not GNAME23863(G23863,G14260);
  and GNAME23864(G23864,G24015,G24016);
  not GNAME23865(G23865,G14259);
  and GNAME23866(G23866,G24018,G24019);
  not GNAME23867(G23867,G14258);
  and GNAME23868(G23868,G24021,G24022);
  not GNAME23869(G23869,G14257);
  and GNAME23870(G23870,G24024,G24025);
  not GNAME23871(G23871,G14256);
  and GNAME23872(G23872,G24027,G24028);
  not GNAME23873(G23873,G14255);
  and GNAME23874(G23874,G24030,G24031);
  not GNAME23875(G23875,G14254);
  and GNAME23876(G23876,G24033,G24034);
  not GNAME23877(G23877,G14253);
  and GNAME23878(G23878,G24036,G24037);
  not GNAME23879(G23879,G14252);
  and GNAME23880(G23880,G24039,G24040);
  not GNAME23881(G23881,G14251);
  and GNAME23882(G23882,G24042,G24043);
  not GNAME23883(G23883,G14250);
  and GNAME23884(G23884,G24045,G24046);
  not GNAME23885(G23885,G14249);
  and GNAME23886(G23886,G24048,G24049);
  not GNAME23887(G23887,G14248);
  and GNAME23888(G23888,G24051,G24052);
  not GNAME23889(G23889,G14247);
  not GNAME23890(G23890,G14246);
  nand GNAME23891(G23891,G24054,G24055);
  nand GNAME23892(G23892,G24058,G24059);
  not GNAME23893(G23893,G14245);
  not GNAME23894(G23894,G14244);
  and GNAME23895(G23895,G23978,G23962);
  nand GNAME23896(G23896,G15181,G14265);
  nand GNAME23897(G23897,G24072,G24073);
  nand GNAME23898(G23898,G20070,G20069);
  nand GNAME23899(G23899,G24112,G24113);
  nand GNAME23900(G23900,G24118,G24119);
  nand GNAME23901(G23901,G24120,G24121);
  nand GNAME23902(G23902,G24125,G24126);
  nand GNAME23903(G23903,G24192,G24193);
  and GNAME23904(G23904,G24104,G24105);
  and GNAME23905(G23905,G24108,G24109);
  and GNAME23906(G23906,G24127,G24128);
  and GNAME23907(G23907,G24131,G24132);
  and GNAME23908(G23908,G24135,G24136);
  and GNAME23909(G23909,G24139,G24140);
  and GNAME23910(G23910,G24143,G24144);
  and GNAME23911(G23911,G24147,G24148);
  and GNAME23912(G23912,G24151,G24152);
  and GNAME23913(G23913,G24155,G24156);
  and GNAME23914(G23914,G24159,G24160);
  and GNAME23915(G23915,G24163,G24164);
  and GNAME23916(G23916,G24169,G24170);
  and GNAME23917(G23917,G24173,G24174);
  and GNAME23918(G23918,G24177,G24178);
  and GNAME23919(G23919,G24181,G24182);
  and GNAME23920(G23920,G24185,G24186);
  and GNAME23921(G23921,G24194,G20080);
  and GNAME23922(G23922,G20077,G20076);
  not GNAME23923(G23923,G14236);
  not GNAME23924(G23924,G14238);
  not GNAME23925(G23925,G14240);
  not GNAME23926(G23926,G14242);
  not GNAME23927(G23927,G14243);
  not GNAME23928(G23928,G14239);
  and GNAME23929(G23929,G23992,G23993);
  and GNAME23930(G23930,G24106,G24107);
  and GNAME23931(G23931,G24110,G24111);
  or GNAME23932(G23932,G23988,G23853);
  nand GNAME23933(G23933,G23984,G23968);
  and GNAME23934(G23934,G23985,G23965);
  and GNAME23935(G23935,G24114,G24115);
  nand GNAME23936(G23936,G23982,G23969);
  and GNAME23937(G23937,G23983,G23968);
  and GNAME23938(G23938,G24116,G24117);
  or GNAME23939(G23939,G23980,G23895);
  and GNAME23940(G23940,G24129,G24130);
  and GNAME23941(G23941,G24133,G24134);
  and GNAME23942(G23942,G24137,G24138);
  and GNAME23943(G23943,G24141,G24142);
  and GNAME23944(G23944,G24145,G24146);
  and GNAME23945(G23945,G24149,G24150);
  and GNAME23946(G23946,G24153,G24154);
  and GNAME23947(G23947,G24157,G24158);
  and GNAME23948(G23948,G24161,G24162);
  and GNAME23949(G23949,G24165,G24166);
  nand GNAME23950(G23950,G23976,G23974);
  and GNAME23951(G23951,G23977,G23971);
  and GNAME23952(G23952,G24167,G24168);
  and GNAME23953(G23953,G24171,G24172);
  and GNAME23954(G23954,G24175,G24176);
  and GNAME23955(G23955,G24179,G24180);
  and GNAME23956(G23956,G24183,G24184);
  and GNAME23957(G23957,G24187,G24188);
  and GNAME23958(G23958,G20079,G20078);
  and GNAME23959(G23959,G20075,G20074);
  nand GNAME23960(G23960,G23975,G23974);
  nand GNAME23961(G23961,G23967,G23843,G23966);
  nand GNAME23962(G23962,G23973,G23845,G23972);
  nand GNAME23963(G23963,G24103,G14268);
  nand GNAME23964(G23964,G23850,G24086,G24087);
  nand GNAME23965(G23965,G24090,G14270);
  or GNAME23966(G23966,G14237,G23842);
  nand GNAME23967(G23967,G23842,G14237);
  nand GNAME23968(G23968,G24102,G14271);
  nand GNAME23969(G23969,G24099,G14272);
  nand GNAME23970(G23970,G23848,G24091,G24092);
  nand GNAME23971(G23971,G24095,G14274);
  or GNAME23972(G23972,G14241,G23842);
  nand GNAME23973(G23973,G23842,G14241);
  nand GNAME23974(G23974,G24098,G14275);
  nand GNAME23975(G23975,G23847,G24096,G24097);
  nand GNAME23976(G23976,G23975,G15181);
  nand GNAME23977(G23977,G23846,G24093,G24094);
  nand GNAME23978(G23978,G23971,G24067);
  nand GNAME23979(G23979,G23972,G23973);
  and GNAME23980(G23980,G23979,G14273);
  not GNAME23981(G23981,G23939);
  nand GNAME23982(G23982,G23970,G23939);
  nand GNAME23983(G23983,G23849,G24100,G24101);
  nand GNAME23984(G23984,G23936,G23983);
  nand GNAME23985(G23985,G23844,G24088,G24089);
  nand GNAME23986(G23986,G23965,G23994);
  nand GNAME23987(G23987,G23966,G23967);
  and GNAME23988(G23988,G23987,G14269);
  not GNAME23989(G23989,G23932);
  nand GNAME23990(G23990,G23964,G23932);
  nand GNAME23991(G23991,G23852,G23851);
  nand GNAME23992(G23992,G23991,G15181);
  or GNAME23993(G23993,G23851,G23852);
  nand GNAME23994(G23994,G23933,G23985);
  nand GNAME23995(G23995,G23961,G20067);
  nand GNAME23996(G23996,G23995,G23965,G23994);
  nand GNAME23997(G23997,G20067,G23853);
  nor GNAME23998(G23998,G14266,G15181);
  not GNAME23999(G23999,G23854);
  or GNAME24000(G24000,G14266,G14264,G23999,G20066);
  nand GNAME24001(G24001,G14264,G23999,G14265);
  nand GNAME24002(G24002,G24000,G15181);
  nand GNAME24003(G24003,G23857,G23856);
  nand GNAME24004(G24004,G24003,G15181);
  or GNAME24005(G24005,G23856,G23857);
  not GNAME24006(G24006,G23859);
  nand GNAME24007(G24007,G23859,G14262);
  nand GNAME24008(G24008,G23842,G24007);
  nand GNAME24009(G24009,G23858,G24006);
  not GNAME24010(G24010,G23860);
  nand GNAME24011(G24011,G23860,G23861);
  nand GNAME24012(G24012,G24011,G15181);
  nand GNAME24013(G24013,G24010,G14261);
  nand GNAME24014(G24014,G23863,G23862);
  nand GNAME24015(G24015,G24014,G15181);
  or GNAME24016(G24016,G23862,G23863);
  nand GNAME24017(G24017,G23865,G23864);
  nand GNAME24018(G24018,G24017,G15181);
  or GNAME24019(G24019,G23864,G23865);
  nand GNAME24020(G24020,G23867,G23866);
  nand GNAME24021(G24021,G24020,G15181);
  or GNAME24022(G24022,G23866,G23867);
  nand GNAME24023(G24023,G23869,G23868);
  nand GNAME24024(G24024,G24023,G15181);
  or GNAME24025(G24025,G23868,G23869);
  nand GNAME24026(G24026,G23871,G23870);
  nand GNAME24027(G24027,G24026,G15181);
  or GNAME24028(G24028,G23870,G23871);
  nand GNAME24029(G24029,G23873,G23872);
  nand GNAME24030(G24030,G24029,G15181);
  or GNAME24031(G24031,G23872,G23873);
  nand GNAME24032(G24032,G23875,G23874);
  nand GNAME24033(G24033,G24032,G15181);
  or GNAME24034(G24034,G23874,G23875);
  nand GNAME24035(G24035,G23877,G23876);
  nand GNAME24036(G24036,G24035,G15181);
  or GNAME24037(G24037,G23876,G23877);
  nand GNAME24038(G24038,G23879,G23878);
  nand GNAME24039(G24039,G24038,G15181);
  or GNAME24040(G24040,G23878,G23879);
  nand GNAME24041(G24041,G23881,G23880);
  nand GNAME24042(G24042,G24041,G15181);
  or GNAME24043(G24043,G23880,G23881);
  nand GNAME24044(G24044,G23883,G23882);
  nand GNAME24045(G24045,G24044,G15181);
  or GNAME24046(G24046,G23882,G23883);
  nand GNAME24047(G24047,G23885,G23884);
  nand GNAME24048(G24048,G24047,G15181);
  or GNAME24049(G24049,G23884,G23885);
  nand GNAME24050(G24050,G23887,G23886);
  nand GNAME24051(G24051,G24050,G15181);
  or GNAME24052(G24052,G23886,G23887);
  nand GNAME24053(G24053,G23889,G23888);
  nand GNAME24054(G24054,G24053,G15181);
  or GNAME24055(G24055,G23888,G23889);
  not GNAME24056(G24056,G23891);
  nand GNAME24057(G24057,G23891,G14246);
  nand GNAME24058(G24058,G23842,G24057);
  nand GNAME24059(G24059,G23890,G24056);
  not GNAME24060(G24060,G23892);
  nand GNAME24061(G24061,G24060,G14245);
  nand GNAME24062(G24062,G23842,G24061);
  nand GNAME24063(G24063,G23893,G23892);
  nand GNAME24064(G24064,G14244,G24062,G24063);
  nand GNAME24065(G24065,G24063,G15181);
  nand GNAME24066(G24066,G24061,G23894,G24065);
  nand GNAME24067(G24067,G23950,G23977);
  nand GNAME24068(G24068,G23962,G20068);
  nand GNAME24069(G24069,G24068,G23971,G24067);
  nand GNAME24070(G24070,G20068,G23895);
  nand GNAME24071(G24071,G23999,G14265);
  nand GNAME24072(G24072,G23842,G24071);
  or GNAME24073(G24073,G14266,G23999);
  nand GNAME24074(G24074,G23896,G23897);
  nand GNAME24075(G24075,G24074,G20071);
  nand GNAME24076(G24076,G20073,G20072,G23896,G23897);
  or GNAME24077(G24077,G14266,G23896);
  nand GNAME24078(G24078,G24077,G15181);
  nand GNAME24079(G24079,G23896,G14265);
  nand GNAME24080(G24080,G24079,G23854,G24078);
  or GNAME24081(G24081,G20066,G23897);
  not GNAME24082(G24082,G23960);
  nand GNAME24083(G24083,G23963,G23964);
  nand GNAME24084(G24084,G23969,G23970);
  nand GNAME24085(G24085,G24064,G24066);
  nand GNAME24086(G24086,G23923,G15181);
  nand GNAME24087(G24087,G23842,G14236);
  nand GNAME24088(G24088,G23924,G15181);
  nand GNAME24089(G24089,G23842,G14238);
  nand GNAME24090(G24090,G24088,G24089);
  nand GNAME24091(G24091,G23925,G15181);
  nand GNAME24092(G24092,G23842,G14240);
  nand GNAME24093(G24093,G23926,G15181);
  nand GNAME24094(G24094,G23842,G14242);
  nand GNAME24095(G24095,G24093,G24094);
  nand GNAME24096(G24096,G23927,G15181);
  nand GNAME24097(G24097,G23842,G14243);
  nand GNAME24098(G24098,G24096,G24097);
  nand GNAME24099(G24099,G24091,G24092);
  nand GNAME24100(G24100,G23928,G15181);
  nand GNAME24101(G24101,G23842,G14239);
  nand GNAME24102(G24102,G24100,G24101);
  nand GNAME24103(G24103,G24086,G24087);
  or GNAME24104(G24104,G14266,G23842);
  nand GNAME24105(G24105,G23842,G14266);
  nand GNAME24106(G24106,G23904,G23929);
  or GNAME24107(G24107,G23929,G23904);
  nand GNAME24108(G24108,G23852,G15181);
  nand GNAME24109(G24109,G23842,G14267);
  nand GNAME24110(G24110,G23851,G23905);
  or GNAME24111(G24111,G23851,G23905);
  nand GNAME24112(G24112,G23932,G24083);
  nand GNAME24113(G24113,G23989,G23963,G23964);
  or GNAME24114(G24114,G23934,G23933);
  nand GNAME24115(G24115,G23933,G23934);
  or GNAME24116(G24116,G23937,G23936);
  nand GNAME24117(G24117,G23936,G23937);
  nand GNAME24118(G24118,G23939,G24084);
  nand GNAME24119(G24119,G23981,G23969,G23970);
  nand GNAME24120(G24120,G24085,G15181);
  nand GNAME24121(G24121,G23842,G24064,G24066);
  nand GNAME24122(G24122,G23893,G15181);
  nand GNAME24123(G24123,G23842,G14245);
  nand GNAME24124(G24124,G24122,G24123);
  nand GNAME24125(G24125,G23892,G24124);
  nand GNAME24126(G24126,G24060,G24122,G24123);
  nand GNAME24127(G24127,G23890,G15181);
  nand GNAME24128(G24128,G23842,G14246);
  nand GNAME24129(G24129,G24056,G23906);
  or GNAME24130(G24130,G24056,G23906);
  nand GNAME24131(G24131,G23889,G15181);
  nand GNAME24132(G24132,G23842,G14247);
  nand GNAME24133(G24133,G23888,G23907);
  or GNAME24134(G24134,G23888,G23907);
  nand GNAME24135(G24135,G23887,G15181);
  nand GNAME24136(G24136,G23842,G14248);
  nand GNAME24137(G24137,G23886,G23908);
  or GNAME24138(G24138,G23886,G23908);
  nand GNAME24139(G24139,G23885,G15181);
  nand GNAME24140(G24140,G23842,G14249);
  nand GNAME24141(G24141,G23884,G23909);
  or GNAME24142(G24142,G23884,G23909);
  nand GNAME24143(G24143,G23883,G15181);
  nand GNAME24144(G24144,G23842,G14250);
  nand GNAME24145(G24145,G23882,G23910);
  or GNAME24146(G24146,G23882,G23910);
  nand GNAME24147(G24147,G23881,G15181);
  nand GNAME24148(G24148,G23842,G14251);
  nand GNAME24149(G24149,G23880,G23911);
  or GNAME24150(G24150,G23880,G23911);
  nand GNAME24151(G24151,G23879,G15181);
  nand GNAME24152(G24152,G23842,G14252);
  nand GNAME24153(G24153,G23878,G23912);
  or GNAME24154(G24154,G23878,G23912);
  nand GNAME24155(G24155,G23877,G15181);
  nand GNAME24156(G24156,G23842,G14253);
  nand GNAME24157(G24157,G23876,G23913);
  or GNAME24158(G24158,G23876,G23913);
  nand GNAME24159(G24159,G23875,G15181);
  nand GNAME24160(G24160,G23842,G14254);
  nand GNAME24161(G24161,G23874,G23914);
  or GNAME24162(G24162,G23874,G23914);
  nand GNAME24163(G24163,G23873,G15181);
  nand GNAME24164(G24164,G23842,G14255);
  nand GNAME24165(G24165,G23872,G23915);
  or GNAME24166(G24166,G23872,G23915);
  or GNAME24167(G24167,G23951,G23950);
  nand GNAME24168(G24168,G23950,G23951);
  nand GNAME24169(G24169,G23871,G15181);
  nand GNAME24170(G24170,G23842,G14256);
  nand GNAME24171(G24171,G23870,G23916);
  or GNAME24172(G24172,G23870,G23916);
  nand GNAME24173(G24173,G23869,G15181);
  nand GNAME24174(G24174,G23842,G14257);
  nand GNAME24175(G24175,G23868,G23917);
  or GNAME24176(G24176,G23868,G23917);
  nand GNAME24177(G24177,G23867,G15181);
  nand GNAME24178(G24178,G23842,G14258);
  nand GNAME24179(G24179,G23866,G23918);
  or GNAME24180(G24180,G23866,G23918);
  nand GNAME24181(G24181,G23865,G15181);
  nand GNAME24182(G24182,G23842,G14259);
  nand GNAME24183(G24183,G23864,G23919);
  or GNAME24184(G24184,G23864,G23919);
  nand GNAME24185(G24185,G23863,G15181);
  nand GNAME24186(G24186,G23842,G14260);
  nand GNAME24187(G24187,G23862,G23920);
  or GNAME24188(G24188,G23862,G23920);
  nand GNAME24189(G24189,G23861,G15181);
  nand GNAME24190(G24190,G23842,G14261);
  nand GNAME24191(G24191,G24189,G24190);
  nand GNAME24192(G24192,G23860,G24191);
  nand GNAME24193(G24193,G24010,G24189,G24190);
  nand GNAME24194(G24194,G23858,G15181);

endmodule