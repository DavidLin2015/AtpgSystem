module b01(CK,G1,G2,G112,G113,G114,G115,G116,G10,G11,G12,G13,G24);
input CK,G1,G2,G112,G113,G114,G115,G116;
output G10,G11,G12,G13,G24;

  wire G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,
       G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,G40,
       G41,G42,G43,G44,G45,G46,G47,G48,G49,G50,G51,G52,G53,G54,G55,G56,G57,G58,G59,G60,
       G61,G62,G63,G64,G65,G66,G67,G68,G69,G70,G71,G72,G73,G74,G75,G76,G77,G78,G79,G80,
       G81,G82,G83,G84,G85,G86,G87,G88,G89,G90,G91,G92,G93,G94,G95,G96,G97,G98,G99,G100,
       G101,G102,G103,G104,G105,G106,G107,G108,G109,G110,G111,G112,G113,G114,G115,G116;

  nand GNAME10(G10,G25,G26,G28,G29);
  nand GNAME11(G11,G25,G32,G21,G39,G40);
  nand GNAME12(G12,G26,G35,G21,G41,G42);
  nand GNAME13(G13,G23,G43,G44);
  and GNAME14(G14,G19,G113);
  not GNAME15(G15,G1);
  nor GNAME16(G16,G113,G18);
  not GNAME17(G17,G112);
  and GNAME18(G18,G2,G1);
  not GNAME19(G19,G114);
  nor GNAME20(G20,G17,G19);
  and GNAME21(G21,G30,G31);
  nand GNAME22(G22,G37,G38);
  or GNAME23(G23,G22,G113,G17);
  and GNAME24(G24,G114,G17,G113);
  nand GNAME25(G25,G17,G14);
  nand GNAME26(G26,G112,G22,G16);
  nand GNAME27(G27,G113,G112);
  nand GNAME28(G28,G27,G18);
  nand GNAME29(G29,G16,G20);
  nand GNAME30(G30,G22,G20);
  nand GNAME31(G31,G14,G18);
  nand GNAME32(G32,G16,G114);
  or GNAME33(G33,G113,G19);
  nand GNAME34(G34,G33,G17);
  nand GNAME35(G35,G16,G17,G19);
  or GNAME36(G36,G14,G17);
  or GNAME37(G37,G2,G15);
  nand GNAME38(G38,G15,G2);
  or GNAME39(G39,G18,G23);
  or GNAME40(G40,G45,G46);
  nand GNAME41(G41,G45,G24);
  nand GNAME42(G42,G34,G18);
  or GNAME43(G43,G46,G22);
  nand GNAME44(G44,G36,G22);
  not GNAME45(G45,G18);
  not GNAME46(G46,G20);

endmodule